magic
tech sky130A
magscale 1 2
timestamp 1750116991
<< viali >>
rect 1685 13957 1719 13991
rect 5549 13957 5583 13991
rect 1133 13889 1167 13923
rect 3341 13889 3375 13923
rect 4261 13889 4295 13923
rect 4537 13889 4571 13923
rect 6837 13889 6871 13923
rect 8309 13889 8343 13923
rect 8677 13889 8711 13923
rect 8861 13889 8895 13923
rect 1869 13821 1903 13855
rect 2605 13821 2639 13855
rect 6561 13821 6595 13855
rect 7849 13821 7883 13855
rect 3525 13753 3559 13787
rect 2421 13685 2455 13719
rect 3157 13685 3191 13719
rect 3617 13685 3651 13719
rect 5917 13685 5951 13719
rect 6653 13685 6687 13719
rect 8493 13685 8527 13719
rect 3985 13481 4019 13515
rect 1133 13345 1167 13379
rect 3157 13345 3191 13379
rect 4629 13345 4663 13379
rect 6377 13345 6411 13379
rect 1869 13277 1903 13311
rect 3709 13277 3743 13311
rect 5365 13277 5399 13311
rect 6837 13277 6871 13311
rect 6929 13277 6963 13311
rect 8125 13277 8159 13311
rect 2513 13209 2547 13243
rect 3525 13209 3559 13243
rect 3893 13209 3927 13243
rect 8677 13209 8711 13243
rect 8861 13209 8895 13243
rect 1685 13141 1719 13175
rect 2421 13141 2455 13175
rect 4721 13141 4755 13175
rect 8493 13141 8527 13175
rect 949 12801 983 12835
rect 5089 12801 5123 12835
rect 6192 12801 6226 12835
rect 6285 12801 6319 12835
rect 8401 12801 8435 12835
rect 1409 12733 1443 12767
rect 2513 12733 2547 12767
rect 3249 12733 3283 12767
rect 3617 12733 3651 12767
rect 6561 12733 6595 12767
rect 6929 12733 6963 12767
rect 3157 12597 3191 12631
rect 5653 12597 5687 12631
rect 6101 12597 6135 12631
rect 8961 12597 8995 12631
rect 1225 12393 1259 12427
rect 7297 12393 7331 12427
rect 1409 12325 1443 12359
rect 3893 12325 3927 12359
rect 3157 12257 3191 12291
rect 4629 12257 4663 12291
rect 7121 12257 7155 12291
rect 1133 12189 1167 12223
rect 3525 12189 3559 12223
rect 3618 12189 3652 12223
rect 4721 12189 4755 12223
rect 5089 12189 5123 12223
rect 6561 12189 6595 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 8707 12189 8741 12223
rect 8861 12189 8895 12223
rect 2881 12121 2915 12155
rect 3985 12053 4019 12087
rect 8125 12053 8159 12087
rect 8493 12053 8527 12087
rect 949 11849 983 11883
rect 8777 11849 8811 11883
rect 6101 11781 6135 11815
rect 2789 11713 2823 11747
rect 5549 11713 5583 11747
rect 6285 11713 6319 11747
rect 6377 11713 6411 11747
rect 8217 11713 8251 11747
rect 2421 11645 2455 11679
rect 2697 11645 2731 11679
rect 3065 11645 3099 11679
rect 4537 11645 4571 11679
rect 4813 11645 4847 11679
rect 6745 11645 6779 11679
rect 5733 11577 5767 11611
rect 5457 11509 5491 11543
rect 5917 11509 5951 11543
rect 2605 11305 2639 11339
rect 3065 11305 3099 11339
rect 6837 11305 6871 11339
rect 2329 11237 2363 11271
rect 2789 11169 2823 11203
rect 3433 11169 3467 11203
rect 3801 11169 3835 11203
rect 2145 11101 2179 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 5273 11101 5307 11135
rect 6193 11101 6227 11135
rect 6929 11101 6963 11135
rect 1041 11033 1075 11067
rect 1869 11033 1903 11067
rect 5837 11033 5871 11067
rect 8125 11033 8159 11067
rect 8677 11033 8711 11067
rect 8861 11033 8895 11067
rect 8493 10965 8527 10999
rect 4537 10761 4571 10795
rect 5273 10761 5307 10795
rect 6469 10761 6503 10795
rect 1041 10693 1075 10727
rect 1869 10625 1903 10659
rect 5548 10625 5582 10659
rect 5641 10625 5675 10659
rect 6101 10625 6135 10659
rect 6255 10625 6289 10659
rect 8401 10625 8435 10659
rect 1961 10557 1995 10591
rect 2237 10557 2271 10591
rect 3801 10557 3835 10591
rect 5089 10557 5123 10591
rect 6561 10557 6595 10591
rect 6929 10557 6963 10591
rect 3709 10489 3743 10523
rect 4445 10421 4479 10455
rect 8961 10421 8995 10455
rect 2053 10217 2087 10251
rect 2513 10217 2547 10251
rect 5365 10217 5399 10251
rect 6745 10217 6779 10251
rect 3341 10149 3375 10183
rect 5825 10149 5859 10183
rect 8493 10149 8527 10183
rect 1041 10081 1075 10115
rect 3065 10081 3099 10115
rect 6561 10081 6595 10115
rect 7849 10081 7883 10115
rect 2237 10013 2271 10047
rect 5089 10013 5123 10047
rect 5273 10013 5307 10047
rect 5917 10013 5951 10047
rect 6837 10013 6871 10047
rect 8309 10013 8343 10047
rect 8768 10013 8802 10047
rect 8861 10013 8895 10047
rect 1869 9945 1903 9979
rect 4813 9945 4847 9979
rect 5641 9945 5675 9979
rect 3893 9673 3927 9707
rect 5733 9673 5767 9707
rect 4261 9605 4295 9639
rect 949 9537 983 9571
rect 2881 9521 2915 9555
rect 3157 9537 3191 9571
rect 3433 9537 3467 9571
rect 3709 9537 3743 9571
rect 6101 9537 6135 9571
rect 8217 9537 8251 9571
rect 1225 9469 1259 9503
rect 2697 9469 2731 9503
rect 3985 9469 4019 9503
rect 6193 9469 6227 9503
rect 6377 9469 6411 9503
rect 6745 9469 6779 9503
rect 3065 9333 3099 9367
rect 3341 9333 3375 9367
rect 3617 9333 3651 9367
rect 8777 9333 8811 9367
rect 2973 9129 3007 9163
rect 3433 9129 3467 9163
rect 4997 9129 5031 9163
rect 7665 9129 7699 9163
rect 8309 9129 8343 9163
rect 8861 9129 8895 9163
rect 4077 9061 4111 9095
rect 1133 8993 1167 9027
rect 6745 8993 6779 9027
rect 2237 8925 2271 8959
rect 2788 8925 2822 8959
rect 2892 8925 2926 8959
rect 3157 8925 3191 8959
rect 3525 8925 3559 8959
rect 3801 8925 3835 8959
rect 4261 8925 4295 8959
rect 4353 8925 4387 8959
rect 6837 8925 6871 8959
rect 6930 8925 6964 8959
rect 7756 8925 7790 8959
rect 7849 8925 7883 8959
rect 8493 8925 8527 8959
rect 8677 8925 8711 8959
rect 6469 8857 6503 8891
rect 7941 8857 7975 8891
rect 8125 8857 8159 8891
rect 2513 8789 2547 8823
rect 3985 8789 4019 8823
rect 4537 8789 4571 8823
rect 7205 8789 7239 8823
rect 4077 8517 4111 8551
rect 4261 8517 4295 8551
rect 1041 8449 1075 8483
rect 1685 8449 1719 8483
rect 3157 8449 3191 8483
rect 3893 8449 3927 8483
rect 6377 8449 6411 8483
rect 8953 8449 8987 8483
rect 1133 8381 1167 8415
rect 1317 8381 1351 8415
rect 3717 8381 3751 8415
rect 6837 8381 6871 8415
rect 8585 8381 8619 8415
rect 7389 8313 7423 8347
rect 6193 8245 6227 8279
rect 6653 8245 6687 8279
rect 2605 7973 2639 8007
rect 1225 7905 1259 7939
rect 2053 7905 2087 7939
rect 7849 7905 7883 7939
rect 2145 7837 2179 7871
rect 4077 7837 4111 7871
rect 5641 7837 5675 7871
rect 6101 7837 6135 7871
rect 6745 7837 6779 7871
rect 8309 7837 8343 7871
rect 8493 7837 8527 7871
rect 8677 7837 8711 7871
rect 1409 7769 1443 7803
rect 5825 7769 5859 7803
rect 1317 7701 1351 7735
rect 1777 7701 1811 7735
rect 2237 7701 2271 7735
rect 4721 7701 4755 7735
rect 6009 7701 6043 7735
rect 8861 7701 8895 7735
rect 1133 7497 1167 7531
rect 1409 7497 1443 7531
rect 2237 7497 2271 7531
rect 3249 7497 3283 7531
rect 8593 7497 8627 7531
rect 8769 7497 8803 7531
rect 4721 7429 4755 7463
rect 949 7361 983 7395
rect 1225 7361 1259 7395
rect 4997 7361 5031 7395
rect 5640 7361 5674 7395
rect 5733 7361 5767 7395
rect 5917 7361 5951 7395
rect 8033 7361 8067 7395
rect 8953 7361 8987 7395
rect 2789 7293 2823 7327
rect 6009 7293 6043 7327
rect 6193 7293 6227 7327
rect 6561 7293 6595 7327
rect 5549 7157 5583 7191
rect 7297 6953 7331 6987
rect 4905 6817 4939 6851
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 6377 6749 6411 6783
rect 7849 6749 7883 6783
rect 8707 6749 8741 6783
rect 8861 6749 8895 6783
rect 6941 6681 6975 6715
rect 8493 6613 8527 6647
rect 1133 6409 1167 6443
rect 5641 6409 5675 6443
rect 4169 6341 4203 6375
rect 949 6273 983 6307
rect 3893 6273 3927 6307
rect 6009 6273 6043 6307
rect 6285 6273 6319 6307
rect 6929 6273 6963 6307
rect 8401 6273 8435 6307
rect 6377 6205 6411 6239
rect 6561 6205 6595 6239
rect 6193 6069 6227 6103
rect 8961 6069 8995 6103
rect 6561 5865 6595 5899
rect 8493 5865 8527 5899
rect 6653 5797 6687 5831
rect 1409 5729 1443 5763
rect 5089 5729 5123 5763
rect 7849 5729 7883 5763
rect 1133 5661 1167 5695
rect 4813 5661 4847 5695
rect 6837 5661 6871 5695
rect 8309 5661 8343 5695
rect 8677 5661 8711 5695
rect 8861 5593 8895 5627
rect 5733 5321 5767 5355
rect 8861 5253 8895 5287
rect 6377 5185 6411 5219
rect 7665 5185 7699 5219
rect 949 5117 983 5151
rect 1225 5117 1259 5151
rect 2697 5117 2731 5151
rect 5089 5117 5123 5151
rect 7389 5117 7423 5151
rect 1133 4777 1167 4811
rect 2145 4709 2179 4743
rect 4905 4709 4939 4743
rect 1501 4641 1535 4675
rect 4261 4641 4295 4675
rect 6653 4641 6687 4675
rect 7849 4641 7883 4675
rect 1317 4573 1351 4607
rect 1961 4573 1995 4607
rect 8309 4573 8343 4607
rect 8707 4573 8741 4607
rect 8861 4573 8895 4607
rect 6377 4505 6411 4539
rect 4813 4437 4847 4471
rect 8493 4437 8527 4471
rect 5549 4233 5583 4267
rect 6285 4233 6319 4267
rect 8961 4233 8995 4267
rect 949 4097 983 4131
rect 3801 4097 3835 4131
rect 6101 4097 6135 4131
rect 6929 4097 6963 4131
rect 8401 4097 8435 4131
rect 6561 4029 6595 4063
rect 1133 3961 1167 3995
rect 4064 3893 4098 3927
rect 3985 3689 4019 3723
rect 7849 3689 7883 3723
rect 8493 3689 8527 3723
rect 7665 3621 7699 3655
rect 5733 3553 5767 3587
rect 5917 3553 5951 3587
rect 6193 3553 6227 3587
rect 7941 3485 7975 3519
rect 8861 3485 8895 3519
rect 5457 3417 5491 3451
rect 8677 3417 8711 3451
rect 8677 3077 8711 3111
rect 4997 3009 5031 3043
rect 5168 3009 5202 3043
rect 5733 3009 5767 3043
rect 7205 3009 7239 3043
rect 7757 3009 7791 3043
rect 8493 3009 8527 3043
rect 4537 2941 4571 2975
rect 7573 2941 7607 2975
rect 8309 2941 8343 2975
rect 8861 2805 8895 2839
rect 2789 2601 2823 2635
rect 5825 2601 5859 2635
rect 8769 2601 8803 2635
rect 4905 2465 4939 2499
rect 6009 2465 6043 2499
rect 6377 2465 6411 2499
rect 2973 2397 3007 2431
rect 3157 2397 3191 2431
rect 4813 2397 4847 2431
rect 5273 2397 5307 2431
rect 7849 2397 7883 2431
rect 8585 2397 8619 2431
rect 8678 2397 8712 2431
rect 8409 2261 8443 2295
rect 7389 2057 7423 2091
rect 9045 2057 9079 2091
rect 5181 1989 5215 2023
rect 8861 1989 8895 2023
rect 4721 1921 4755 1955
rect 4905 1921 4939 1955
rect 6837 1921 6871 1955
rect 6930 1921 6964 1955
rect 7481 1921 7515 1955
rect 8677 1921 8711 1955
rect 4353 1853 4387 1887
rect 6653 1785 6687 1819
rect 7021 1717 7055 1751
rect 8861 1513 8895 1547
rect 7389 1377 7423 1411
rect 6377 1309 6411 1343
rect 9045 1309 9079 1343
<< metal1 >>
rect 3602 14424 3608 14476
rect 3660 14464 3666 14476
rect 5718 14464 5724 14476
rect 3660 14436 5724 14464
rect 3660 14424 3666 14436
rect 5718 14424 5724 14436
rect 5776 14424 5782 14476
rect 3234 14356 3240 14408
rect 3292 14396 3298 14408
rect 8202 14396 8208 14408
rect 3292 14368 8208 14396
rect 3292 14356 3298 14368
rect 8202 14356 8208 14368
rect 8260 14356 8266 14408
rect 4614 14288 4620 14340
rect 4672 14328 4678 14340
rect 7098 14328 7104 14340
rect 4672 14300 7104 14328
rect 4672 14288 4678 14300
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 1118 14220 1124 14272
rect 1176 14260 1182 14272
rect 6270 14260 6276 14272
rect 1176 14232 6276 14260
rect 1176 14220 1182 14232
rect 6270 14220 6276 14232
rect 6328 14220 6334 14272
rect 6362 14220 6368 14272
rect 6420 14260 6426 14272
rect 6822 14260 6828 14272
rect 6420 14232 6828 14260
rect 6420 14220 6426 14232
rect 6822 14220 6828 14232
rect 6880 14220 6886 14272
rect 644 14170 9384 14192
rect 644 14118 2954 14170
rect 3006 14118 3018 14170
rect 3070 14118 3082 14170
rect 3134 14118 6954 14170
rect 7006 14118 7018 14170
rect 7070 14118 7082 14170
rect 7134 14118 9384 14170
rect 644 14096 9384 14118
rect 4798 14056 4804 14068
rect 1136 14028 4804 14056
rect 1136 13929 1164 14028
rect 4798 14016 4804 14028
rect 4856 14016 4862 14068
rect 7650 14056 7656 14068
rect 5000 14028 7656 14056
rect 1673 13991 1731 13997
rect 1673 13957 1685 13991
rect 1719 13988 1731 13991
rect 4154 13988 4160 14000
rect 1719 13960 4160 13988
rect 1719 13957 1731 13960
rect 1673 13951 1731 13957
rect 4154 13948 4160 13960
rect 4212 13948 4218 14000
rect 5000 13988 5028 14028
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 4264 13960 5028 13988
rect 5537 13991 5595 13997
rect 1121 13923 1179 13929
rect 1121 13889 1133 13923
rect 1167 13889 1179 13923
rect 1121 13883 1179 13889
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13920 3387 13923
rect 3970 13920 3976 13932
rect 3375 13892 3976 13920
rect 3375 13889 3387 13892
rect 3329 13883 3387 13889
rect 3970 13880 3976 13892
rect 4028 13880 4034 13932
rect 4264 13929 4292 13960
rect 5537 13957 5549 13991
rect 5583 13988 5595 13991
rect 9582 13988 9588 14000
rect 5583 13960 9588 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 4249 13923 4307 13929
rect 4249 13889 4261 13923
rect 4295 13889 4307 13923
rect 4249 13883 4307 13889
rect 4525 13923 4583 13929
rect 4525 13889 4537 13923
rect 4571 13920 4583 13923
rect 4706 13920 4712 13932
rect 4571 13892 4712 13920
rect 4571 13889 4583 13892
rect 4525 13883 4583 13889
rect 4706 13880 4712 13892
rect 4764 13880 4770 13932
rect 6825 13923 6883 13929
rect 6825 13889 6837 13923
rect 6871 13920 6883 13923
rect 7650 13920 7656 13932
rect 6871 13892 7656 13920
rect 6871 13889 6883 13892
rect 6825 13883 6883 13889
rect 7650 13880 7656 13892
rect 7708 13880 7714 13932
rect 8297 13923 8355 13929
rect 8297 13889 8309 13923
rect 8343 13920 8355 13923
rect 8570 13920 8576 13932
rect 8343 13892 8576 13920
rect 8343 13889 8355 13892
rect 8297 13883 8355 13889
rect 8570 13880 8576 13892
rect 8628 13880 8634 13932
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 1857 13855 1915 13861
rect 1857 13821 1869 13855
rect 1903 13821 1915 13855
rect 1857 13815 1915 13821
rect 2593 13855 2651 13861
rect 2593 13821 2605 13855
rect 2639 13852 2651 13855
rect 3234 13852 3240 13864
rect 2639 13824 3240 13852
rect 2639 13821 2651 13824
rect 2593 13815 2651 13821
rect 1872 13784 1900 13815
rect 3234 13812 3240 13824
rect 3292 13812 3298 13864
rect 6549 13855 6607 13861
rect 3436 13824 5304 13852
rect 3436 13784 3464 13824
rect 1872 13756 3464 13784
rect 3513 13787 3571 13793
rect 3513 13753 3525 13787
rect 3559 13784 3571 13787
rect 5166 13784 5172 13796
rect 3559 13756 5172 13784
rect 3559 13753 3571 13756
rect 3513 13747 3571 13753
rect 5166 13744 5172 13756
rect 5224 13744 5230 13796
rect 5276 13784 5304 13824
rect 6549 13821 6561 13855
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8478 13852 8484 13864
rect 7883 13824 8484 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 6362 13784 6368 13796
rect 5276 13756 6368 13784
rect 6362 13744 6368 13756
rect 6420 13744 6426 13796
rect 6564 13784 6592 13815
rect 8478 13812 8484 13824
rect 8536 13812 8542 13864
rect 8680 13852 8708 13883
rect 8846 13880 8852 13932
rect 8904 13880 8910 13932
rect 9214 13852 9220 13864
rect 8680 13824 9220 13852
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 8018 13784 8024 13796
rect 6564 13756 8024 13784
rect 8018 13744 8024 13756
rect 8076 13744 8082 13796
rect 2314 13676 2320 13728
rect 2372 13716 2378 13728
rect 2409 13719 2467 13725
rect 2409 13716 2421 13719
rect 2372 13688 2421 13716
rect 2372 13676 2378 13688
rect 2409 13685 2421 13688
rect 2455 13685 2467 13719
rect 2409 13679 2467 13685
rect 2774 13676 2780 13728
rect 2832 13716 2838 13728
rect 3145 13719 3203 13725
rect 3145 13716 3157 13719
rect 2832 13688 3157 13716
rect 2832 13676 2838 13688
rect 3145 13685 3157 13688
rect 3191 13685 3203 13719
rect 3145 13679 3203 13685
rect 3605 13719 3663 13725
rect 3605 13685 3617 13719
rect 3651 13716 3663 13719
rect 4062 13716 4068 13728
rect 3651 13688 4068 13716
rect 3651 13685 3663 13688
rect 3605 13679 3663 13685
rect 4062 13676 4068 13688
rect 4120 13676 4126 13728
rect 4982 13676 4988 13728
rect 5040 13716 5046 13728
rect 5905 13719 5963 13725
rect 5905 13716 5917 13719
rect 5040 13688 5917 13716
rect 5040 13676 5046 13688
rect 5905 13685 5917 13688
rect 5951 13685 5963 13719
rect 5905 13679 5963 13685
rect 6178 13676 6184 13728
rect 6236 13716 6242 13728
rect 6641 13719 6699 13725
rect 6641 13716 6653 13719
rect 6236 13688 6653 13716
rect 6236 13676 6242 13688
rect 6641 13685 6653 13688
rect 6687 13685 6699 13719
rect 6641 13679 6699 13685
rect 8110 13676 8116 13728
rect 8168 13716 8174 13728
rect 8481 13719 8539 13725
rect 8481 13716 8493 13719
rect 8168 13688 8493 13716
rect 8168 13676 8174 13688
rect 8481 13685 8493 13688
rect 8527 13685 8539 13719
rect 8481 13679 8539 13685
rect 644 13626 9384 13648
rect 644 13574 2554 13626
rect 2606 13574 2618 13626
rect 2670 13574 2682 13626
rect 2734 13574 6554 13626
rect 6606 13574 6618 13626
rect 6670 13574 6682 13626
rect 6734 13574 9384 13626
rect 644 13552 9384 13574
rect 3970 13472 3976 13524
rect 4028 13472 4034 13524
rect 5994 13512 6000 13524
rect 4080 13484 6000 13512
rect 4080 13444 4108 13484
rect 5994 13472 6000 13484
rect 6052 13472 6058 13524
rect 9030 13512 9036 13524
rect 6196 13484 9036 13512
rect 2746 13416 4108 13444
rect 1118 13336 1124 13388
rect 1176 13336 1182 13388
rect 1857 13311 1915 13317
rect 1857 13277 1869 13311
rect 1903 13308 1915 13311
rect 2746 13308 2774 13416
rect 4522 13404 4528 13456
rect 4580 13444 4586 13456
rect 4580 13416 5304 13444
rect 4580 13404 4586 13416
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13376 3203 13379
rect 3602 13376 3608 13388
rect 3191 13348 3608 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 3602 13336 3608 13348
rect 3660 13336 3666 13388
rect 4614 13336 4620 13388
rect 4672 13336 4678 13388
rect 1903 13280 2774 13308
rect 3697 13311 3755 13317
rect 1903 13277 1915 13280
rect 1857 13271 1915 13277
rect 3697 13277 3709 13311
rect 3743 13308 3755 13311
rect 4430 13308 4436 13320
rect 3743 13280 4436 13308
rect 3743 13277 3755 13280
rect 3697 13271 3755 13277
rect 4430 13268 4436 13280
rect 4488 13268 4494 13320
rect 2222 13200 2228 13252
rect 2280 13240 2286 13252
rect 2501 13243 2559 13249
rect 2501 13240 2513 13243
rect 2280 13212 2513 13240
rect 2280 13200 2286 13212
rect 2501 13209 2513 13212
rect 2547 13209 2559 13243
rect 2501 13203 2559 13209
rect 3513 13243 3571 13249
rect 3513 13209 3525 13243
rect 3559 13240 3571 13243
rect 3602 13240 3608 13252
rect 3559 13212 3608 13240
rect 3559 13209 3571 13212
rect 3513 13203 3571 13209
rect 3602 13200 3608 13212
rect 3660 13200 3666 13252
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 5074 13240 5080 13252
rect 3927 13212 5080 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 5276 13240 5304 13416
rect 5350 13404 5356 13456
rect 5408 13444 5414 13456
rect 6196 13444 6224 13484
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 7190 13444 7196 13456
rect 5408 13416 6224 13444
rect 6288 13416 7196 13444
rect 5408 13404 5414 13416
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13308 5411 13311
rect 6288 13308 6316 13416
rect 7190 13404 7196 13416
rect 7248 13404 7254 13456
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 9582 13376 9588 13388
rect 6411 13348 9588 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 9582 13336 9588 13348
rect 9640 13336 9646 13388
rect 5399 13280 6316 13308
rect 5399 13277 5411 13280
rect 5353 13271 5411 13277
rect 6822 13268 6828 13320
rect 6880 13268 6886 13320
rect 6917 13311 6975 13317
rect 6917 13277 6929 13311
rect 6963 13277 6975 13311
rect 6917 13271 6975 13277
rect 8113 13311 8171 13317
rect 8113 13277 8125 13311
rect 8159 13308 8171 13311
rect 9122 13308 9128 13320
rect 8159 13280 9128 13308
rect 8159 13277 8171 13280
rect 8113 13271 8171 13277
rect 5626 13240 5632 13252
rect 5276 13212 5632 13240
rect 5626 13200 5632 13212
rect 5684 13200 5690 13252
rect 5902 13200 5908 13252
rect 5960 13240 5966 13252
rect 6932 13240 6960 13271
rect 9122 13268 9128 13280
rect 9180 13268 9186 13320
rect 5960 13212 6960 13240
rect 8665 13243 8723 13249
rect 5960 13200 5966 13212
rect 8665 13209 8677 13243
rect 8711 13209 8723 13243
rect 8665 13203 8723 13209
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 1673 13175 1731 13181
rect 1673 13172 1685 13175
rect 1636 13144 1685 13172
rect 1636 13132 1642 13144
rect 1673 13141 1685 13144
rect 1719 13141 1731 13175
rect 1673 13135 1731 13141
rect 1762 13132 1768 13184
rect 1820 13172 1826 13184
rect 2409 13175 2467 13181
rect 2409 13172 2421 13175
rect 1820 13144 2421 13172
rect 1820 13132 1826 13144
rect 2409 13141 2421 13144
rect 2455 13141 2467 13175
rect 2409 13135 2467 13141
rect 4246 13132 4252 13184
rect 4304 13172 4310 13184
rect 4709 13175 4767 13181
rect 4709 13172 4721 13175
rect 4304 13144 4721 13172
rect 4304 13132 4310 13144
rect 4709 13141 4721 13144
rect 4755 13141 4767 13175
rect 4709 13135 4767 13141
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8260 13144 8493 13172
rect 8260 13132 8266 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8680 13172 8708 13203
rect 8754 13200 8760 13252
rect 8812 13240 8818 13252
rect 8849 13243 8907 13249
rect 8849 13240 8861 13243
rect 8812 13212 8861 13240
rect 8812 13200 8818 13212
rect 8849 13209 8861 13212
rect 8895 13209 8907 13243
rect 8849 13203 8907 13209
rect 9214 13172 9220 13184
rect 8680 13144 9220 13172
rect 8481 13135 8539 13141
rect 9214 13132 9220 13144
rect 9272 13132 9278 13184
rect 644 13082 9384 13104
rect 644 13030 2954 13082
rect 3006 13030 3018 13082
rect 3070 13030 3082 13082
rect 3134 13030 6954 13082
rect 7006 13030 7018 13082
rect 7070 13030 7082 13082
rect 7134 13030 9384 13082
rect 644 13008 9384 13030
rect 6454 12928 6460 12980
rect 6512 12968 6518 12980
rect 6512 12940 7236 12968
rect 6512 12928 6518 12940
rect 4154 12860 4160 12912
rect 4212 12860 4218 12912
rect 7208 12900 7236 12940
rect 6196 12872 6408 12900
rect 7208 12872 7314 12900
rect 934 12792 940 12844
rect 992 12792 998 12844
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 6196 12841 6224 12872
rect 6180 12835 6238 12841
rect 6180 12801 6192 12835
rect 6226 12801 6238 12835
rect 6180 12795 6238 12801
rect 6270 12792 6276 12844
rect 6328 12792 6334 12844
rect 6380 12832 6408 12872
rect 6380 12804 6684 12832
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 1544 12736 2513 12764
rect 1544 12724 1550 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 3234 12724 3240 12776
rect 3292 12724 3298 12776
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3344 12736 3617 12764
rect 3344 12696 3372 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 5994 12724 6000 12776
rect 6052 12764 6058 12776
rect 6549 12767 6607 12773
rect 6549 12764 6561 12767
rect 6052 12736 6561 12764
rect 6052 12724 6058 12736
rect 6549 12733 6561 12736
rect 6595 12733 6607 12767
rect 6549 12727 6607 12733
rect 3160 12668 3372 12696
rect 2774 12588 2780 12640
rect 2832 12628 2838 12640
rect 3160 12637 3188 12668
rect 3145 12631 3203 12637
rect 3145 12628 3157 12631
rect 2832 12600 3157 12628
rect 2832 12588 2838 12600
rect 3145 12597 3157 12600
rect 3191 12597 3203 12631
rect 3145 12591 3203 12597
rect 5641 12631 5699 12637
rect 5641 12597 5653 12631
rect 5687 12628 5699 12631
rect 5810 12628 5816 12640
rect 5687 12600 5816 12628
rect 5687 12597 5699 12600
rect 5641 12591 5699 12597
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 6086 12588 6092 12640
rect 6144 12588 6150 12640
rect 6656 12628 6684 12804
rect 8386 12792 8392 12844
rect 8444 12792 8450 12844
rect 6822 12724 6828 12776
rect 6880 12764 6886 12776
rect 6917 12767 6975 12773
rect 6917 12764 6929 12767
rect 6880 12736 6929 12764
rect 6880 12724 6886 12736
rect 6917 12733 6929 12736
rect 6963 12733 6975 12767
rect 6917 12727 6975 12733
rect 8846 12628 8852 12640
rect 6656 12600 8852 12628
rect 8846 12588 8852 12600
rect 8904 12588 8910 12640
rect 8938 12588 8944 12640
rect 8996 12637 9002 12640
rect 8996 12591 9007 12637
rect 8996 12588 9002 12591
rect 644 12538 9384 12560
rect 644 12486 2554 12538
rect 2606 12486 2618 12538
rect 2670 12486 2682 12538
rect 2734 12486 6554 12538
rect 6606 12486 6618 12538
rect 6670 12486 6682 12538
rect 6734 12486 9384 12538
rect 644 12464 9384 12486
rect 1213 12427 1271 12433
rect 1213 12393 1225 12427
rect 1259 12424 1271 12427
rect 3234 12424 3240 12436
rect 1259 12396 3240 12424
rect 1259 12393 1271 12396
rect 1213 12387 1271 12393
rect 3234 12384 3240 12396
rect 3292 12384 3298 12436
rect 6362 12424 6368 12436
rect 4816 12396 6368 12424
rect 1397 12359 1455 12365
rect 1397 12325 1409 12359
rect 1443 12356 1455 12359
rect 1486 12356 1492 12368
rect 1443 12328 1492 12356
rect 1443 12325 1455 12328
rect 1397 12319 1455 12325
rect 1486 12316 1492 12328
rect 1544 12316 1550 12368
rect 3881 12359 3939 12365
rect 3881 12325 3893 12359
rect 3927 12356 3939 12359
rect 4154 12356 4160 12368
rect 3927 12328 4160 12356
rect 3927 12325 3939 12328
rect 3881 12319 3939 12325
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 2130 12248 2136 12300
rect 2188 12288 2194 12300
rect 3145 12291 3203 12297
rect 3145 12288 3157 12291
rect 2188 12260 3157 12288
rect 2188 12248 2194 12260
rect 3145 12257 3157 12260
rect 3191 12257 3203 12291
rect 4617 12291 4675 12297
rect 3145 12251 3203 12257
rect 3436 12260 4200 12288
rect 1121 12223 1179 12229
rect 1121 12189 1133 12223
rect 1167 12220 1179 12223
rect 1210 12220 1216 12232
rect 1167 12192 1216 12220
rect 1167 12189 1179 12192
rect 1121 12183 1179 12189
rect 1210 12180 1216 12192
rect 1268 12180 1274 12232
rect 1394 12112 1400 12164
rect 1452 12152 1458 12164
rect 2869 12155 2927 12161
rect 1452 12124 1702 12152
rect 1452 12112 1458 12124
rect 1596 12084 1624 12124
rect 2869 12121 2881 12155
rect 2915 12152 2927 12155
rect 3436 12152 3464 12260
rect 4172 12232 4200 12260
rect 4617 12257 4629 12291
rect 4663 12288 4675 12291
rect 4816 12288 4844 12396
rect 6362 12384 6368 12396
rect 6420 12384 6426 12436
rect 7285 12427 7343 12433
rect 7285 12393 7297 12427
rect 7331 12424 7343 12427
rect 7650 12424 7656 12436
rect 7331 12396 7656 12424
rect 7331 12393 7343 12396
rect 7285 12387 7343 12393
rect 7650 12384 7656 12396
rect 7708 12384 7714 12436
rect 7190 12356 7196 12368
rect 7116 12328 7196 12356
rect 7116 12297 7144 12328
rect 7190 12316 7196 12328
rect 7248 12316 7254 12368
rect 4663 12260 4844 12288
rect 7109 12291 7167 12297
rect 4663 12257 4675 12260
rect 4617 12251 4675 12257
rect 7109 12257 7121 12291
rect 7155 12257 7167 12291
rect 8110 12288 8116 12300
rect 7109 12251 7167 12257
rect 7484 12260 8116 12288
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 2915 12124 3464 12152
rect 2915 12121 2927 12124
rect 2869 12115 2927 12121
rect 3528 12084 3556 12183
rect 3602 12180 3608 12232
rect 3660 12220 3666 12232
rect 3660 12192 3705 12220
rect 3660 12180 3666 12192
rect 4154 12180 4160 12232
rect 4212 12180 4218 12232
rect 4706 12180 4712 12232
rect 4764 12180 4770 12232
rect 5074 12180 5080 12232
rect 5132 12180 5138 12232
rect 6549 12223 6607 12229
rect 6549 12189 6561 12223
rect 6595 12220 6607 12223
rect 7484 12220 7512 12260
rect 8110 12248 8116 12260
rect 8168 12248 8174 12300
rect 6595 12192 7512 12220
rect 6595 12189 6607 12192
rect 6549 12183 6607 12189
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 7837 12223 7895 12229
rect 7837 12220 7849 12223
rect 7708 12192 7849 12220
rect 7708 12180 7714 12192
rect 7837 12189 7849 12192
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 8662 12180 8668 12232
rect 8720 12229 8726 12232
rect 8720 12223 8753 12229
rect 8741 12189 8753 12223
rect 8720 12183 8753 12189
rect 8849 12223 8907 12229
rect 8849 12189 8861 12223
rect 8895 12220 8907 12223
rect 9214 12220 9220 12232
rect 8895 12192 9220 12220
rect 8895 12189 8907 12192
rect 8849 12183 8907 12189
rect 8720 12180 8726 12183
rect 6086 12112 6092 12164
rect 6144 12112 6150 12164
rect 8864 12152 8892 12183
rect 9214 12180 9220 12192
rect 9272 12180 9278 12232
rect 8772 12124 8892 12152
rect 8772 12096 8800 12124
rect 3602 12084 3608 12096
rect 1596 12056 3608 12084
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 3973 12087 4031 12093
rect 3973 12053 3985 12087
rect 4019 12084 4031 12087
rect 4062 12084 4068 12096
rect 4019 12056 4068 12084
rect 4019 12053 4031 12056
rect 3973 12047 4031 12053
rect 4062 12044 4068 12056
rect 4120 12044 4126 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 7650 12084 7656 12096
rect 5592 12056 7656 12084
rect 5592 12044 5598 12056
rect 7650 12044 7656 12056
rect 7708 12044 7714 12096
rect 8110 12044 8116 12096
rect 8168 12044 8174 12096
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 8754 12044 8760 12096
rect 8812 12044 8818 12096
rect 644 11994 9384 12016
rect 644 11942 2954 11994
rect 3006 11942 3018 11994
rect 3070 11942 3082 11994
rect 3134 11942 6954 11994
rect 7006 11942 7018 11994
rect 7070 11942 7082 11994
rect 7134 11942 9384 11994
rect 644 11920 9384 11942
rect 934 11840 940 11892
rect 992 11840 998 11892
rect 2406 11840 2412 11892
rect 2464 11880 2470 11892
rect 5718 11880 5724 11892
rect 2464 11852 5724 11880
rect 2464 11840 2470 11852
rect 5718 11840 5724 11852
rect 5776 11840 5782 11892
rect 6270 11880 6276 11892
rect 6104 11852 6276 11880
rect 1394 11772 1400 11824
rect 1452 11772 1458 11824
rect 2130 11772 2136 11824
rect 2188 11812 2194 11824
rect 2188 11784 2819 11812
rect 2188 11772 2194 11784
rect 2791 11753 2819 11784
rect 3602 11772 3608 11824
rect 3660 11772 3666 11824
rect 5442 11772 5448 11824
rect 5500 11812 5506 11824
rect 6104 11821 6132 11852
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 8110 11880 8116 11892
rect 6380 11852 8116 11880
rect 6089 11815 6147 11821
rect 6089 11812 6101 11815
rect 5500 11784 6101 11812
rect 5500 11772 5506 11784
rect 6089 11781 6101 11784
rect 6135 11781 6147 11815
rect 6089 11775 6147 11781
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 5350 11704 5356 11756
rect 5408 11744 5414 11756
rect 5537 11747 5595 11753
rect 5537 11744 5549 11747
rect 5408 11716 5549 11744
rect 5408 11704 5414 11716
rect 5537 11713 5549 11716
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 6178 11704 6184 11756
rect 6236 11744 6242 11756
rect 6380 11753 6408 11852
rect 8110 11840 8116 11852
rect 8168 11840 8174 11892
rect 8570 11840 8576 11892
rect 8628 11880 8634 11892
rect 8765 11883 8823 11889
rect 8765 11880 8777 11883
rect 8628 11852 8777 11880
rect 8628 11840 8634 11852
rect 8765 11849 8777 11852
rect 8811 11849 8823 11883
rect 8765 11843 8823 11849
rect 8478 11812 8484 11824
rect 7866 11784 8484 11812
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 6273 11747 6331 11753
rect 6273 11744 6285 11747
rect 6236 11716 6285 11744
rect 6236 11704 6242 11716
rect 6273 11713 6285 11716
rect 6319 11713 6331 11747
rect 6273 11707 6331 11713
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6365 11707 6423 11713
rect 8202 11704 8208 11756
rect 8260 11704 8266 11756
rect 2406 11636 2412 11688
rect 2464 11636 2470 11688
rect 2685 11679 2743 11685
rect 2685 11645 2697 11679
rect 2731 11645 2743 11679
rect 3053 11679 3111 11685
rect 3053 11676 3065 11679
rect 2685 11639 2743 11645
rect 2792 11648 3065 11676
rect 2700 11540 2728 11639
rect 2792 11620 2820 11648
rect 3053 11645 3065 11648
rect 3099 11645 3111 11679
rect 3053 11639 3111 11645
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11676 4583 11679
rect 4801 11679 4859 11685
rect 4801 11676 4813 11679
rect 4571 11648 4813 11676
rect 4571 11645 4583 11648
rect 4525 11639 4583 11645
rect 4801 11645 4813 11648
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 6086 11636 6092 11688
rect 6144 11676 6150 11688
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 6144 11648 6745 11676
rect 6144 11636 6150 11648
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 2774 11568 2780 11620
rect 2832 11568 2838 11620
rect 5721 11611 5779 11617
rect 5721 11577 5733 11611
rect 5767 11608 5779 11611
rect 6270 11608 6276 11620
rect 5767 11580 6276 11608
rect 5767 11577 5779 11580
rect 5721 11571 5779 11577
rect 6270 11568 6276 11580
rect 6328 11568 6334 11620
rect 4522 11540 4528 11552
rect 2700 11512 4528 11540
rect 4522 11500 4528 11512
rect 4580 11500 4586 11552
rect 4798 11500 4804 11552
rect 4856 11540 4862 11552
rect 5074 11540 5080 11552
rect 4856 11512 5080 11540
rect 4856 11500 4862 11512
rect 5074 11500 5080 11512
rect 5132 11540 5138 11552
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 5132 11512 5457 11540
rect 5132 11500 5138 11512
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 5445 11503 5503 11509
rect 5902 11500 5908 11552
rect 5960 11500 5966 11552
rect 644 11450 9384 11472
rect 644 11398 2554 11450
rect 2606 11398 2618 11450
rect 2670 11398 2682 11450
rect 2734 11398 6554 11450
rect 6606 11398 6618 11450
rect 6670 11398 6682 11450
rect 6734 11398 9384 11450
rect 644 11376 9384 11398
rect 2593 11339 2651 11345
rect 2593 11305 2605 11339
rect 2639 11336 2651 11339
rect 2774 11336 2780 11348
rect 2639 11308 2780 11336
rect 2639 11305 2651 11308
rect 2593 11299 2651 11305
rect 2774 11296 2780 11308
rect 2832 11296 2838 11348
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 4706 11336 4712 11348
rect 3099 11308 4712 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 6822 11296 6828 11348
rect 6880 11296 6886 11348
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 3234 11268 3240 11280
rect 2363 11240 3240 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 3234 11228 3240 11240
rect 3292 11228 3298 11280
rect 2777 11203 2835 11209
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3421 11203 3479 11209
rect 3421 11200 3433 11203
rect 2823 11172 3096 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 2130 11092 2136 11144
rect 2188 11092 2194 11144
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2280 11104 2421 11132
rect 2280 11092 2286 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2731 11104 2973 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 1026 11024 1032 11076
rect 1084 11024 1090 11076
rect 1857 11067 1915 11073
rect 1857 11033 1869 11067
rect 1903 11064 1915 11067
rect 1946 11064 1952 11076
rect 1903 11036 1952 11064
rect 1903 11033 1915 11036
rect 1857 11027 1915 11033
rect 1946 11024 1952 11036
rect 2004 11024 2010 11076
rect 2792 11008 2820 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 3068 11132 3096 11172
rect 3252 11172 3433 11200
rect 3252 11132 3280 11172
rect 3421 11169 3433 11172
rect 3467 11169 3479 11203
rect 3421 11163 3479 11169
rect 3789 11203 3847 11209
rect 3789 11169 3801 11203
rect 3835 11200 3847 11203
rect 4154 11200 4160 11212
rect 3835 11172 4160 11200
rect 3835 11169 3847 11172
rect 3789 11163 3847 11169
rect 4154 11160 4160 11172
rect 4212 11160 4218 11212
rect 5902 11200 5908 11212
rect 5276 11172 5908 11200
rect 5276 11141 5304 11172
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 3068 11104 3280 11132
rect 5261 11135 5319 11141
rect 2961 11095 3019 11101
rect 5261 11101 5273 11135
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 5718 11092 5724 11144
rect 5776 11132 5782 11144
rect 6181 11135 6239 11141
rect 6181 11132 6193 11135
rect 5776 11104 6193 11132
rect 5776 11092 5782 11104
rect 6181 11101 6193 11104
rect 6227 11101 6239 11135
rect 6181 11095 6239 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 4896 11076 4948 11082
rect 5825 11067 5883 11073
rect 5825 11033 5837 11067
rect 5871 11064 5883 11067
rect 6932 11064 6960 11095
rect 5871 11036 6960 11064
rect 5871 11033 5883 11036
rect 5825 11027 5883 11033
rect 8110 11024 8116 11076
rect 8168 11024 8174 11076
rect 8662 11064 8668 11076
rect 8220 11036 8668 11064
rect 4896 11018 4948 11024
rect 2774 10956 2780 11008
rect 2832 10956 2838 11008
rect 5626 10956 5632 11008
rect 5684 10996 5690 11008
rect 6822 10996 6828 11008
rect 5684 10968 6828 10996
rect 5684 10956 5690 10968
rect 6822 10956 6828 10968
rect 6880 10996 6886 11008
rect 8220 10996 8248 11036
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 8754 11024 8760 11076
rect 8812 11064 8818 11076
rect 8849 11067 8907 11073
rect 8849 11064 8861 11067
rect 8812 11036 8861 11064
rect 8812 11024 8818 11036
rect 8849 11033 8861 11036
rect 8895 11033 8907 11067
rect 8849 11027 8907 11033
rect 6880 10968 8248 10996
rect 6880 10956 6886 10968
rect 8478 10956 8484 11008
rect 8536 10956 8542 11008
rect 644 10906 9384 10928
rect 644 10854 2954 10906
rect 3006 10854 3018 10906
rect 3070 10854 3082 10906
rect 3134 10854 6954 10906
rect 7006 10854 7018 10906
rect 7070 10854 7082 10906
rect 7134 10854 9384 10906
rect 644 10832 9384 10854
rect 4154 10752 4160 10804
rect 4212 10792 4218 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4212 10764 4537 10792
rect 4212 10752 4218 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 4890 10752 4896 10804
rect 4948 10792 4954 10804
rect 5261 10795 5319 10801
rect 5261 10792 5273 10795
rect 4948 10764 5273 10792
rect 4948 10752 4954 10764
rect 5261 10761 5273 10764
rect 5307 10761 5319 10795
rect 6178 10792 6184 10804
rect 5261 10755 5319 10761
rect 5552 10764 6184 10792
rect 382 10684 388 10736
rect 440 10724 446 10736
rect 1029 10727 1087 10733
rect 1029 10724 1041 10727
rect 440 10696 1041 10724
rect 440 10684 446 10696
rect 1029 10693 1041 10696
rect 1075 10693 1087 10727
rect 3602 10724 3608 10736
rect 3450 10696 3608 10724
rect 1029 10687 1087 10693
rect 3602 10684 3608 10696
rect 3660 10724 3666 10736
rect 3660 10696 5488 10724
rect 3660 10684 3666 10696
rect 1857 10659 1915 10665
rect 1857 10625 1869 10659
rect 1903 10625 1915 10659
rect 1857 10619 1915 10625
rect 1210 10412 1216 10464
rect 1268 10452 1274 10464
rect 1872 10452 1900 10619
rect 1946 10548 1952 10600
rect 2004 10548 2010 10600
rect 2222 10548 2228 10600
rect 2280 10548 2286 10600
rect 3234 10548 3240 10600
rect 3292 10588 3298 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3292 10560 3801 10588
rect 3292 10548 3298 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 3789 10551 3847 10557
rect 4126 10560 5089 10588
rect 3697 10523 3755 10529
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 4126 10520 4154 10560
rect 5077 10557 5089 10560
rect 5123 10557 5135 10591
rect 5460 10588 5488 10696
rect 5552 10665 5580 10764
rect 6178 10752 6184 10764
rect 6236 10752 6242 10804
rect 6454 10752 6460 10804
rect 6512 10752 6518 10804
rect 6822 10792 6828 10804
rect 6564 10764 6828 10792
rect 6564 10724 6592 10764
rect 6822 10752 6828 10764
rect 6880 10752 6886 10804
rect 8202 10724 8208 10736
rect 6104 10696 6592 10724
rect 8050 10696 8208 10724
rect 5536 10659 5594 10665
rect 5536 10625 5548 10659
rect 5582 10625 5594 10659
rect 5536 10619 5594 10625
rect 5626 10616 5632 10668
rect 5684 10656 5690 10668
rect 5684 10628 5764 10656
rect 5684 10616 5690 10628
rect 5736 10588 5764 10628
rect 5810 10616 5816 10668
rect 5868 10656 5874 10668
rect 6104 10665 6132 10696
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 6270 10665 6276 10668
rect 6089 10659 6147 10665
rect 6089 10656 6101 10659
rect 5868 10628 6101 10656
rect 5868 10616 5874 10628
rect 6089 10625 6101 10628
rect 6135 10625 6147 10659
rect 6089 10619 6147 10625
rect 6243 10659 6276 10665
rect 6243 10625 6255 10659
rect 6243 10619 6276 10625
rect 6270 10616 6276 10619
rect 6328 10616 6334 10668
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 8478 10656 8484 10668
rect 8435 10628 8484 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 5460 10560 5764 10588
rect 5077 10551 5135 10557
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 6512 10560 6561 10588
rect 6512 10548 6518 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6917 10591 6975 10597
rect 6917 10588 6929 10591
rect 6549 10551 6607 10557
rect 6656 10560 6929 10588
rect 3743 10492 4154 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 6656 10520 6684 10560
rect 6917 10557 6929 10560
rect 6963 10557 6975 10591
rect 6917 10551 6975 10557
rect 9030 10520 9036 10532
rect 6236 10492 6684 10520
rect 8312 10492 9036 10520
rect 6236 10480 6242 10492
rect 2774 10452 2780 10464
rect 1268 10424 2780 10452
rect 1268 10412 1274 10424
rect 2774 10412 2780 10424
rect 2832 10412 2838 10464
rect 4246 10412 4252 10464
rect 4304 10452 4310 10464
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 4304 10424 4445 10452
rect 4304 10412 4310 10424
rect 4433 10421 4445 10424
rect 4479 10421 4491 10455
rect 4433 10415 4491 10421
rect 5166 10412 5172 10464
rect 5224 10452 5230 10464
rect 8312 10452 8340 10492
rect 9030 10480 9036 10492
rect 9088 10480 9094 10532
rect 5224 10424 8340 10452
rect 5224 10412 5230 10424
rect 8386 10412 8392 10464
rect 8444 10452 8450 10464
rect 8949 10455 9007 10461
rect 8949 10452 8961 10455
rect 8444 10424 8961 10452
rect 8444 10412 8450 10424
rect 8949 10421 8961 10424
rect 8995 10421 9007 10455
rect 8949 10415 9007 10421
rect 644 10362 9384 10384
rect 644 10310 2554 10362
rect 2606 10310 2618 10362
rect 2670 10310 2682 10362
rect 2734 10310 6554 10362
rect 6606 10310 6618 10362
rect 6670 10310 6682 10362
rect 6734 10310 9384 10362
rect 644 10288 9384 10310
rect 1394 10208 1400 10260
rect 1452 10248 1458 10260
rect 1670 10248 1676 10260
rect 1452 10220 1676 10248
rect 1452 10208 1458 10220
rect 1670 10208 1676 10220
rect 1728 10248 1734 10260
rect 2041 10251 2099 10257
rect 2041 10248 2053 10251
rect 1728 10220 2053 10248
rect 1728 10208 1734 10220
rect 2041 10217 2053 10220
rect 2087 10217 2099 10251
rect 2041 10211 2099 10217
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2501 10251 2559 10257
rect 2501 10248 2513 10251
rect 2280 10220 2513 10248
rect 2280 10208 2286 10220
rect 2501 10217 2513 10220
rect 2547 10217 2559 10251
rect 2501 10211 2559 10217
rect 2774 10208 2780 10260
rect 2832 10248 2838 10260
rect 5353 10251 5411 10257
rect 2832 10220 5304 10248
rect 2832 10208 2838 10220
rect 3234 10140 3240 10192
rect 3292 10180 3298 10192
rect 3329 10183 3387 10189
rect 3329 10180 3341 10183
rect 3292 10152 3341 10180
rect 3292 10140 3298 10152
rect 3329 10149 3341 10152
rect 3375 10149 3387 10183
rect 3329 10143 3387 10149
rect 474 10072 480 10124
rect 532 10112 538 10124
rect 1029 10115 1087 10121
rect 1029 10112 1041 10115
rect 532 10084 1041 10112
rect 532 10072 538 10084
rect 1029 10081 1041 10084
rect 1075 10081 1087 10115
rect 1029 10075 1087 10081
rect 2038 10072 2044 10124
rect 2096 10112 2102 10124
rect 3053 10115 3111 10121
rect 3053 10112 3065 10115
rect 2096 10084 3065 10112
rect 2096 10072 2102 10084
rect 3053 10081 3065 10084
rect 3099 10081 3111 10115
rect 3053 10075 3111 10081
rect 3602 10072 3608 10124
rect 3660 10112 3666 10124
rect 3660 10084 3740 10112
rect 3660 10072 3666 10084
rect 2130 10004 2136 10056
rect 2188 10044 2194 10056
rect 2225 10047 2283 10053
rect 2225 10044 2237 10047
rect 2188 10016 2237 10044
rect 2188 10004 2194 10016
rect 2225 10013 2237 10016
rect 2271 10013 2283 10047
rect 3712 10030 3740 10084
rect 2225 10007 2283 10013
rect 5074 10004 5080 10056
rect 5132 10004 5138 10056
rect 5276 10053 5304 10220
rect 5353 10217 5365 10251
rect 5399 10248 5411 10251
rect 5994 10248 6000 10260
rect 5399 10220 6000 10248
rect 5399 10217 5411 10220
rect 5353 10211 5411 10217
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6454 10208 6460 10260
rect 6512 10248 6518 10260
rect 6733 10251 6791 10257
rect 6733 10248 6745 10251
rect 6512 10220 6745 10248
rect 6512 10208 6518 10220
rect 6733 10217 6745 10220
rect 6779 10217 6791 10251
rect 6733 10211 6791 10217
rect 5810 10140 5816 10192
rect 5868 10140 5874 10192
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8481 10183 8539 10189
rect 8481 10180 8493 10183
rect 8260 10152 8493 10180
rect 8260 10140 8266 10152
rect 8481 10149 8493 10152
rect 8527 10149 8539 10183
rect 8481 10143 8539 10149
rect 5534 10072 5540 10124
rect 5592 10112 5598 10124
rect 6454 10112 6460 10124
rect 5592 10084 6460 10112
rect 5592 10072 5598 10084
rect 6454 10072 6460 10084
rect 6512 10112 6518 10124
rect 6549 10115 6607 10121
rect 6549 10112 6561 10115
rect 6512 10084 6561 10112
rect 6512 10072 6518 10084
rect 6549 10081 6561 10084
rect 6595 10081 6607 10115
rect 6549 10075 6607 10081
rect 7837 10115 7895 10121
rect 7837 10081 7849 10115
rect 7883 10112 7895 10115
rect 9582 10112 9588 10124
rect 7883 10084 9588 10112
rect 7883 10081 7895 10084
rect 7837 10075 7895 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 5261 10047 5319 10053
rect 5261 10013 5273 10047
rect 5307 10044 5319 10047
rect 5307 10016 5764 10044
rect 5307 10013 5319 10016
rect 5261 10007 5319 10013
rect 1854 9936 1860 9988
rect 1912 9936 1918 9988
rect 4801 9979 4859 9985
rect 4801 9945 4813 9979
rect 4847 9976 4859 9979
rect 5534 9976 5540 9988
rect 4847 9948 5540 9976
rect 4847 9945 4859 9948
rect 4801 9939 4859 9945
rect 5534 9936 5540 9948
rect 5592 9936 5598 9988
rect 5626 9936 5632 9988
rect 5684 9936 5690 9988
rect 5736 9976 5764 10016
rect 5902 10004 5908 10056
rect 5960 10004 5966 10056
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 8018 10044 8024 10056
rect 6871 10016 8024 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 5994 9976 6000 9988
rect 5736 9948 6000 9976
rect 5994 9936 6000 9948
rect 6052 9976 6058 9988
rect 6840 9976 6868 10007
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 8297 10047 8355 10053
rect 8297 10013 8309 10047
rect 8343 10044 8355 10047
rect 8386 10044 8392 10056
rect 8343 10016 8392 10044
rect 8343 10013 8355 10016
rect 8297 10007 8355 10013
rect 8386 10004 8392 10016
rect 8444 10004 8450 10056
rect 8570 10004 8576 10056
rect 8628 10044 8634 10056
rect 8754 10046 8760 10056
rect 8680 10044 8760 10046
rect 8628 10018 8760 10044
rect 8628 10016 8708 10018
rect 8628 10004 8634 10016
rect 8754 10004 8760 10018
rect 8812 10004 8818 10056
rect 8849 10047 8907 10053
rect 8849 10013 8861 10047
rect 8895 10013 8907 10047
rect 8849 10007 8907 10013
rect 8864 9976 8892 10007
rect 6052 9948 6868 9976
rect 8680 9948 8892 9976
rect 6052 9936 6058 9948
rect 8680 9920 8708 9948
rect 2314 9868 2320 9920
rect 2372 9908 2378 9920
rect 3234 9908 3240 9920
rect 2372 9880 3240 9908
rect 2372 9868 2378 9880
rect 3234 9868 3240 9880
rect 3292 9868 3298 9920
rect 6270 9868 6276 9920
rect 6328 9908 6334 9920
rect 8018 9908 8024 9920
rect 6328 9880 8024 9908
rect 6328 9868 6334 9880
rect 8018 9868 8024 9880
rect 8076 9868 8082 9920
rect 8662 9868 8668 9920
rect 8720 9868 8726 9920
rect 644 9818 9384 9840
rect 644 9766 2954 9818
rect 3006 9766 3018 9818
rect 3070 9766 3082 9818
rect 3134 9766 6954 9818
rect 7006 9766 7018 9818
rect 7070 9766 7082 9818
rect 7134 9766 9384 9818
rect 644 9744 9384 9766
rect 1946 9704 1952 9716
rect 952 9676 1952 9704
rect 952 9577 980 9676
rect 1946 9664 1952 9676
rect 2004 9704 2010 9716
rect 2004 9676 2544 9704
rect 2004 9664 2010 9676
rect 1670 9596 1676 9648
rect 1728 9596 1734 9648
rect 2516 9636 2544 9676
rect 2774 9664 2780 9716
rect 2832 9704 2838 9716
rect 3881 9707 3939 9713
rect 2832 9676 3188 9704
rect 2832 9664 2838 9676
rect 3160 9674 3188 9676
rect 3160 9646 3280 9674
rect 3881 9673 3893 9707
rect 3927 9704 3939 9707
rect 4890 9704 4896 9716
rect 3927 9676 4896 9704
rect 3927 9673 3939 9676
rect 3881 9667 3939 9673
rect 4890 9664 4896 9676
rect 4948 9664 4954 9716
rect 5718 9664 5724 9716
rect 5776 9664 5782 9716
rect 3252 9636 3280 9646
rect 3970 9636 3976 9648
rect 2516 9608 3004 9636
rect 3252 9608 3464 9636
rect 937 9571 995 9577
rect 937 9537 949 9571
rect 983 9537 995 9571
rect 2869 9555 2927 9561
rect 2869 9552 2881 9555
rect 937 9531 995 9537
rect 2791 9524 2881 9552
rect 1213 9503 1271 9509
rect 1213 9469 1225 9503
rect 1259 9500 1271 9503
rect 1670 9500 1676 9512
rect 1259 9472 1676 9500
rect 1259 9469 1271 9472
rect 1213 9463 1271 9469
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 1946 9460 1952 9512
rect 2004 9500 2010 9512
rect 2685 9503 2743 9509
rect 2685 9500 2697 9503
rect 2004 9472 2697 9500
rect 2004 9460 2010 9472
rect 2685 9469 2697 9472
rect 2731 9469 2743 9503
rect 2685 9463 2743 9469
rect 2406 9392 2412 9444
rect 2464 9432 2470 9444
rect 2791 9432 2819 9524
rect 2869 9521 2881 9524
rect 2915 9521 2927 9555
rect 2869 9515 2927 9521
rect 2464 9404 2819 9432
rect 2976 9432 3004 9608
rect 3436 9577 3464 9608
rect 3804 9608 3976 9636
rect 3145 9571 3203 9577
rect 3145 9537 3157 9571
rect 3191 9570 3203 9571
rect 3421 9571 3479 9577
rect 3191 9542 3280 9570
rect 3191 9537 3203 9542
rect 3145 9531 3203 9537
rect 3252 9512 3280 9542
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9568 3755 9571
rect 3804 9568 3832 9608
rect 3970 9596 3976 9608
rect 4028 9596 4034 9648
rect 4246 9596 4252 9648
rect 4304 9596 4310 9648
rect 5810 9636 5816 9648
rect 5474 9608 5816 9636
rect 5810 9596 5816 9608
rect 5868 9596 5874 9648
rect 7650 9596 7656 9648
rect 7708 9596 7714 9648
rect 3743 9540 3832 9568
rect 3743 9537 3755 9540
rect 3697 9531 3755 9537
rect 5994 9528 6000 9580
rect 6052 9568 6058 9580
rect 6089 9571 6147 9577
rect 6089 9568 6101 9571
rect 6052 9540 6101 9568
rect 6052 9528 6058 9540
rect 6089 9537 6101 9540
rect 6135 9537 6147 9571
rect 6089 9531 6147 9537
rect 8205 9571 8263 9577
rect 8205 9537 8217 9571
rect 8251 9568 8263 9571
rect 8846 9568 8852 9580
rect 8251 9540 8852 9568
rect 8251 9537 8263 9540
rect 8205 9531 8263 9537
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 3234 9460 3240 9512
rect 3292 9460 3298 9512
rect 3973 9503 4031 9509
rect 3973 9469 3985 9503
rect 4019 9500 4031 9503
rect 4982 9500 4988 9512
rect 4019 9472 4988 9500
rect 4019 9469 4031 9472
rect 3973 9463 4031 9469
rect 3988 9432 4016 9463
rect 4982 9460 4988 9472
rect 5040 9460 5046 9512
rect 6181 9503 6239 9509
rect 6181 9469 6193 9503
rect 6227 9500 6239 9503
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 6227 9472 6377 9500
rect 6227 9469 6239 9472
rect 6181 9463 6239 9469
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 6365 9463 6423 9469
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6733 9503 6791 9509
rect 6733 9500 6745 9503
rect 6512 9472 6745 9500
rect 6512 9460 6518 9472
rect 6733 9469 6745 9472
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 8570 9432 8576 9444
rect 2976 9404 4016 9432
rect 8128 9404 8576 9432
rect 2464 9392 2470 9404
rect 2774 9324 2780 9376
rect 2832 9364 2838 9376
rect 3053 9367 3111 9373
rect 3053 9364 3065 9367
rect 2832 9336 3065 9364
rect 2832 9324 2838 9336
rect 3053 9333 3065 9336
rect 3099 9333 3111 9367
rect 3053 9327 3111 9333
rect 3234 9324 3240 9376
rect 3292 9364 3298 9376
rect 3329 9367 3387 9373
rect 3329 9364 3341 9367
rect 3292 9336 3341 9364
rect 3292 9324 3298 9336
rect 3329 9333 3341 9336
rect 3375 9333 3387 9367
rect 3329 9327 3387 9333
rect 3605 9367 3663 9373
rect 3605 9333 3617 9367
rect 3651 9364 3663 9367
rect 8128 9364 8156 9404
rect 8570 9392 8576 9404
rect 8628 9392 8634 9444
rect 3651 9336 8156 9364
rect 3651 9333 3663 9336
rect 3605 9327 3663 9333
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 8765 9367 8823 9373
rect 8765 9364 8777 9367
rect 8260 9336 8777 9364
rect 8260 9324 8266 9336
rect 8765 9333 8777 9336
rect 8811 9333 8823 9367
rect 8765 9327 8823 9333
rect 644 9274 9384 9296
rect 644 9222 2554 9274
rect 2606 9222 2618 9274
rect 2670 9222 2682 9274
rect 2734 9222 6554 9274
rect 6606 9222 6618 9274
rect 6670 9222 6682 9274
rect 6734 9222 9384 9274
rect 644 9200 9384 9222
rect 2961 9163 3019 9169
rect 2961 9160 2973 9163
rect 2746 9132 2973 9160
rect 2746 9092 2774 9132
rect 2961 9129 2973 9132
rect 3007 9129 3019 9163
rect 2961 9123 3019 9129
rect 3421 9163 3479 9169
rect 3421 9129 3433 9163
rect 3467 9160 3479 9163
rect 4522 9160 4528 9172
rect 3467 9132 4528 9160
rect 3467 9129 3479 9132
rect 3421 9123 3479 9129
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 4985 9163 5043 9169
rect 4985 9129 4997 9163
rect 5031 9160 5043 9163
rect 5902 9160 5908 9172
rect 5031 9132 5908 9160
rect 5031 9129 5043 9132
rect 4985 9123 5043 9129
rect 5902 9120 5908 9132
rect 5960 9120 5966 9172
rect 7650 9120 7656 9172
rect 7708 9120 7714 9172
rect 8294 9120 8300 9172
rect 8352 9120 8358 9172
rect 8846 9120 8852 9172
rect 8904 9120 8910 9172
rect 4065 9095 4123 9101
rect 4065 9092 4077 9095
rect 2700 9064 2774 9092
rect 2976 9064 4077 9092
rect 382 8984 388 9036
rect 440 9024 446 9036
rect 1121 9027 1179 9033
rect 1121 9024 1133 9027
rect 440 8996 1133 9024
rect 440 8984 446 8996
rect 1121 8993 1133 8996
rect 1167 8993 1179 9027
rect 1121 8987 1179 8993
rect 2222 8916 2228 8968
rect 2280 8916 2286 8968
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 2464 8792 2513 8820
rect 2464 8780 2470 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2700 8820 2728 9064
rect 2976 9024 3004 9064
rect 4065 9061 4077 9064
rect 4111 9092 4123 9095
rect 4430 9092 4436 9104
rect 4111 9064 4436 9092
rect 4111 9061 4123 9064
rect 4065 9055 4123 9061
rect 4430 9052 4436 9064
rect 4488 9052 4494 9104
rect 5074 9024 5080 9036
rect 2791 8996 3004 9024
rect 3528 8996 5080 9024
rect 2791 8965 2819 8996
rect 2884 8965 3096 8966
rect 3528 8965 3556 8996
rect 5074 8984 5080 8996
rect 5132 9024 5138 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 5132 8996 6745 9024
rect 5132 8984 5138 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 7668 8996 8524 9024
rect 2776 8959 2834 8965
rect 2776 8925 2788 8959
rect 2822 8925 2834 8959
rect 2776 8919 2834 8925
rect 2880 8959 3096 8965
rect 2880 8925 2892 8959
rect 2926 8938 3096 8959
rect 2926 8925 2938 8938
rect 2880 8919 2938 8925
rect 2774 8820 2780 8832
rect 2700 8792 2780 8820
rect 2501 8783 2559 8789
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 3068 8820 3096 8938
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8925 3203 8959
rect 3145 8919 3203 8925
rect 3513 8959 3571 8965
rect 3513 8925 3525 8959
rect 3559 8925 3571 8959
rect 3513 8919 3571 8925
rect 3789 8959 3847 8965
rect 3789 8925 3801 8959
rect 3835 8956 3847 8959
rect 4062 8956 4068 8968
rect 3835 8928 4068 8956
rect 3835 8925 3847 8928
rect 3789 8919 3847 8925
rect 3160 8888 3188 8919
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4246 8916 4252 8968
rect 4304 8916 4310 8968
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8956 4399 8959
rect 5166 8956 5172 8968
rect 4387 8928 5172 8956
rect 4387 8925 4399 8928
rect 4341 8919 4399 8925
rect 5166 8916 5172 8928
rect 5224 8916 5230 8968
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 6918 8959 6976 8965
rect 6918 8925 6930 8959
rect 6964 8952 6976 8959
rect 7190 8956 7196 8968
rect 7116 8952 7196 8956
rect 6964 8928 7196 8952
rect 6964 8925 7144 8928
rect 6918 8924 7144 8925
rect 6918 8919 6976 8924
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 4154 8888 4160 8900
rect 3160 8860 4160 8888
rect 4154 8848 4160 8860
rect 4212 8848 4218 8900
rect 5810 8848 5816 8900
rect 5868 8848 5874 8900
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 6236 8860 6469 8888
rect 6236 8848 6242 8860
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 7668 8888 7696 8996
rect 8496 8965 8524 8996
rect 7744 8959 7802 8965
rect 7744 8925 7756 8959
rect 7790 8925 7802 8959
rect 7744 8919 7802 8925
rect 7837 8959 7895 8965
rect 7837 8925 7849 8959
rect 7883 8956 7895 8959
rect 8481 8959 8539 8965
rect 7883 8928 8156 8956
rect 7883 8925 7895 8928
rect 7837 8919 7895 8925
rect 7760 8888 7788 8919
rect 6457 8851 6515 8857
rect 7024 8860 7788 8888
rect 7929 8891 7987 8897
rect 3602 8820 3608 8832
rect 3068 8792 3608 8820
rect 3602 8780 3608 8792
rect 3660 8780 3666 8832
rect 3973 8823 4031 8829
rect 3973 8789 3985 8823
rect 4019 8820 4031 8823
rect 4338 8820 4344 8832
rect 4019 8792 4344 8820
rect 4019 8789 4031 8792
rect 3973 8783 4031 8789
rect 4338 8780 4344 8792
rect 4396 8780 4402 8832
rect 4525 8823 4583 8829
rect 4525 8789 4537 8823
rect 4571 8820 4583 8823
rect 7024 8820 7052 8860
rect 7929 8857 7941 8891
rect 7975 8888 7987 8891
rect 8018 8888 8024 8900
rect 7975 8860 8024 8888
rect 7975 8857 7987 8860
rect 7929 8851 7987 8857
rect 8018 8848 8024 8860
rect 8076 8848 8082 8900
rect 8128 8897 8156 8928
rect 8481 8925 8493 8959
rect 8527 8925 8539 8959
rect 8481 8919 8539 8925
rect 8662 8916 8668 8968
rect 8720 8916 8726 8968
rect 8113 8891 8171 8897
rect 8113 8857 8125 8891
rect 8159 8888 8171 8891
rect 8680 8888 8708 8916
rect 8159 8860 8708 8888
rect 8159 8857 8171 8860
rect 8113 8851 8171 8857
rect 4571 8792 7052 8820
rect 7193 8823 7251 8829
rect 4571 8789 4583 8792
rect 4525 8783 4583 8789
rect 7193 8789 7205 8823
rect 7239 8820 7251 8823
rect 7650 8820 7656 8832
rect 7239 8792 7656 8820
rect 7239 8789 7251 8792
rect 7193 8783 7251 8789
rect 7650 8780 7656 8792
rect 7708 8780 7714 8832
rect 644 8730 9384 8752
rect 644 8678 2954 8730
rect 3006 8678 3018 8730
rect 3070 8678 3082 8730
rect 3134 8678 6954 8730
rect 7006 8678 7018 8730
rect 7070 8678 7082 8730
rect 7134 8678 9384 8730
rect 644 8656 9384 8678
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3660 8588 4108 8616
rect 3660 8576 3666 8588
rect 2406 8508 2412 8560
rect 2464 8508 2470 8560
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 4080 8557 4108 8588
rect 4338 8576 4344 8628
rect 4396 8616 4402 8628
rect 7190 8616 7196 8628
rect 4396 8588 7196 8616
rect 4396 8576 4402 8588
rect 7190 8576 7196 8588
rect 7248 8616 7254 8628
rect 8478 8616 8484 8628
rect 7248 8588 8484 8616
rect 7248 8576 7254 8588
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 4065 8551 4123 8557
rect 3292 8520 4016 8548
rect 3292 8508 3298 8520
rect 1029 8483 1087 8489
rect 1029 8449 1041 8483
rect 1075 8480 1087 8483
rect 1210 8480 1216 8492
rect 1075 8452 1216 8480
rect 1075 8449 1087 8452
rect 1029 8443 1087 8449
rect 1210 8440 1216 8452
rect 1268 8440 1274 8492
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8480 3203 8483
rect 3881 8483 3939 8489
rect 3881 8480 3893 8483
rect 3191 8452 3893 8480
rect 3191 8449 3203 8452
rect 3145 8443 3203 8449
rect 3881 8449 3893 8452
rect 3927 8449 3939 8483
rect 3988 8480 4016 8520
rect 4065 8517 4077 8551
rect 4111 8517 4123 8551
rect 4065 8511 4123 8517
rect 4249 8551 4307 8557
rect 4249 8517 4261 8551
rect 4295 8548 4307 8551
rect 4430 8548 4436 8560
rect 4295 8520 4436 8548
rect 4295 8517 4307 8520
rect 4249 8511 4307 8517
rect 4430 8508 4436 8520
rect 4488 8508 4494 8560
rect 5718 8508 5724 8560
rect 5776 8548 5782 8560
rect 6822 8548 6828 8560
rect 5776 8520 6828 8548
rect 5776 8508 5782 8520
rect 6822 8508 6828 8520
rect 6880 8548 6886 8560
rect 8662 8548 8668 8560
rect 6880 8520 8668 8548
rect 6880 8508 6886 8520
rect 8662 8508 8668 8520
rect 8720 8508 8726 8560
rect 5810 8480 5816 8492
rect 3988 8452 5816 8480
rect 3881 8443 3939 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8449 6423 8483
rect 6365 8443 6423 8449
rect 1121 8415 1179 8421
rect 1121 8381 1133 8415
rect 1167 8412 1179 8415
rect 1305 8415 1363 8421
rect 1305 8412 1317 8415
rect 1167 8384 1317 8412
rect 1167 8381 1179 8384
rect 1121 8375 1179 8381
rect 1305 8381 1317 8384
rect 1351 8381 1363 8415
rect 1305 8375 1363 8381
rect 3602 8372 3608 8424
rect 3660 8412 3666 8424
rect 3705 8415 3763 8421
rect 3705 8412 3717 8415
rect 3660 8384 3717 8412
rect 3660 8372 3666 8384
rect 3705 8381 3717 8384
rect 3751 8381 3763 8415
rect 3705 8375 3763 8381
rect 6380 8344 6408 8443
rect 8938 8440 8944 8492
rect 8996 8440 9002 8492
rect 6822 8372 6828 8424
rect 6880 8372 6886 8424
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 9582 8412 9588 8424
rect 8619 8384 9588 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 2608 8316 6408 8344
rect 1578 8236 1584 8288
rect 1636 8276 1642 8288
rect 2608 8276 2636 8316
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 7377 8347 7435 8353
rect 7377 8344 7389 8347
rect 6512 8316 7389 8344
rect 6512 8304 6518 8316
rect 7377 8313 7389 8316
rect 7423 8313 7435 8347
rect 7377 8307 7435 8313
rect 1636 8248 2636 8276
rect 1636 8236 1642 8248
rect 5626 8236 5632 8288
rect 5684 8276 5690 8288
rect 6181 8279 6239 8285
rect 6181 8276 6193 8279
rect 5684 8248 6193 8276
rect 5684 8236 5690 8248
rect 6181 8245 6193 8248
rect 6227 8245 6239 8279
rect 6181 8239 6239 8245
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 7190 8276 7196 8288
rect 6687 8248 7196 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 644 8186 9384 8208
rect 644 8134 2554 8186
rect 2606 8134 2618 8186
rect 2670 8134 2682 8186
rect 2734 8134 6554 8186
rect 6606 8134 6618 8186
rect 6670 8134 6682 8186
rect 6734 8134 9384 8186
rect 644 8112 9384 8134
rect 1394 8032 1400 8084
rect 1452 8072 1458 8084
rect 2774 8072 2780 8084
rect 1452 8044 2780 8072
rect 1452 8032 1458 8044
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 1762 7964 1768 8016
rect 1820 8004 1826 8016
rect 2314 8004 2320 8016
rect 1820 7976 2320 8004
rect 1820 7964 1826 7976
rect 2314 7964 2320 7976
rect 2372 7964 2378 8016
rect 2593 8007 2651 8013
rect 2593 7973 2605 8007
rect 2639 8004 2651 8007
rect 6362 8004 6368 8016
rect 2639 7976 6368 8004
rect 2639 7973 2651 7976
rect 2593 7967 2651 7973
rect 6362 7964 6368 7976
rect 6420 7964 6426 8016
rect 1213 7939 1271 7945
rect 1213 7905 1225 7939
rect 1259 7936 1271 7939
rect 2041 7939 2099 7945
rect 2041 7936 2053 7939
rect 1259 7908 2053 7936
rect 1259 7905 1271 7908
rect 1213 7899 1271 7905
rect 2041 7905 2053 7908
rect 2087 7936 2099 7939
rect 2774 7936 2780 7948
rect 2087 7908 2780 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 2774 7896 2780 7908
rect 2832 7936 2838 7948
rect 3602 7936 3608 7948
rect 2832 7908 3608 7936
rect 2832 7896 2838 7908
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8386 7936 8392 7948
rect 7883 7908 8392 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 1118 7828 1124 7880
rect 1176 7868 1182 7880
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 1176 7840 2145 7868
rect 1176 7828 1182 7840
rect 2133 7837 2145 7840
rect 2179 7837 2191 7871
rect 2133 7831 2191 7837
rect 2314 7828 2320 7880
rect 2372 7868 2378 7880
rect 2372 7840 3188 7868
rect 2372 7828 2378 7840
rect 1394 7760 1400 7812
rect 1452 7760 1458 7812
rect 3160 7800 3188 7840
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3292 7840 4077 7868
rect 3292 7828 3298 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 4706 7828 4712 7880
rect 4764 7868 4770 7880
rect 5350 7868 5356 7880
rect 4764 7840 5356 7868
rect 4764 7828 4770 7840
rect 5350 7828 5356 7840
rect 5408 7868 5414 7880
rect 5534 7868 5540 7880
rect 5408 7840 5540 7868
rect 5408 7828 5414 7840
rect 5534 7828 5540 7840
rect 5592 7828 5598 7880
rect 5626 7828 5632 7880
rect 5684 7828 5690 7880
rect 5736 7840 5948 7868
rect 5736 7800 5764 7840
rect 1780 7772 2774 7800
rect 3160 7772 5764 7800
rect 5813 7803 5871 7809
rect 1302 7692 1308 7744
rect 1360 7692 1366 7744
rect 1780 7741 1808 7772
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7701 1823 7735
rect 1765 7695 1823 7701
rect 1946 7692 1952 7744
rect 2004 7732 2010 7744
rect 2225 7735 2283 7741
rect 2225 7732 2237 7735
rect 2004 7704 2237 7732
rect 2004 7692 2010 7704
rect 2225 7701 2237 7704
rect 2271 7701 2283 7735
rect 2746 7732 2774 7772
rect 5813 7769 5825 7803
rect 5859 7769 5871 7803
rect 5920 7800 5948 7840
rect 6086 7828 6092 7880
rect 6144 7828 6150 7880
rect 6270 7828 6276 7880
rect 6328 7868 6334 7880
rect 6733 7871 6791 7877
rect 6733 7868 6745 7871
rect 6328 7840 6745 7868
rect 6328 7828 6334 7840
rect 6733 7837 6745 7840
rect 6779 7837 6791 7871
rect 6733 7831 6791 7837
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 8662 7828 8668 7880
rect 8720 7828 8726 7880
rect 8110 7800 8116 7812
rect 5920 7772 8116 7800
rect 5813 7763 5871 7769
rect 4614 7732 4620 7744
rect 2746 7704 4620 7732
rect 2225 7695 2283 7701
rect 4614 7692 4620 7704
rect 4672 7692 4678 7744
rect 4709 7735 4767 7741
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 4890 7732 4896 7744
rect 4755 7704 4896 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 4890 7692 4896 7704
rect 4948 7692 4954 7744
rect 5718 7692 5724 7744
rect 5776 7732 5782 7744
rect 5828 7732 5856 7763
rect 8110 7760 8116 7772
rect 8168 7760 8174 7812
rect 5776 7704 5856 7732
rect 5997 7735 6055 7741
rect 5776 7692 5782 7704
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 6362 7732 6368 7744
rect 6043 7704 6368 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 8849 7735 8907 7741
rect 8849 7732 8861 7735
rect 8076 7704 8861 7732
rect 8076 7692 8082 7704
rect 8849 7701 8861 7704
rect 8895 7701 8907 7735
rect 8849 7695 8907 7701
rect 644 7642 9384 7664
rect 644 7590 2954 7642
rect 3006 7590 3018 7642
rect 3070 7590 3082 7642
rect 3134 7590 6954 7642
rect 7006 7590 7018 7642
rect 7070 7590 7082 7642
rect 7134 7590 9384 7642
rect 644 7568 9384 7590
rect 1121 7531 1179 7537
rect 1121 7497 1133 7531
rect 1167 7497 1179 7531
rect 1121 7491 1179 7497
rect 1136 7460 1164 7491
rect 1394 7488 1400 7540
rect 1452 7488 1458 7540
rect 1670 7488 1676 7540
rect 1728 7528 1734 7540
rect 2225 7531 2283 7537
rect 2225 7528 2237 7531
rect 1728 7500 2237 7528
rect 1728 7488 1734 7500
rect 2225 7497 2237 7500
rect 2271 7497 2283 7531
rect 2225 7491 2283 7497
rect 3234 7488 3240 7540
rect 3292 7488 3298 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8581 7531 8639 7537
rect 8581 7528 8593 7531
rect 8352 7500 8593 7528
rect 8352 7488 8358 7500
rect 8581 7497 8593 7500
rect 8627 7497 8639 7531
rect 8581 7491 8639 7497
rect 8754 7488 8760 7540
rect 8812 7488 8818 7540
rect 7656 7472 7708 7478
rect 1946 7460 1952 7472
rect 1136 7432 1952 7460
rect 1946 7420 1952 7432
rect 2004 7420 2010 7472
rect 4709 7463 4767 7469
rect 4709 7429 4721 7463
rect 4755 7460 4767 7463
rect 4798 7460 4804 7472
rect 4755 7432 4804 7460
rect 4755 7429 4767 7432
rect 4709 7423 4767 7429
rect 4798 7420 4804 7432
rect 4856 7420 4862 7472
rect 7656 7414 7708 7420
rect 934 7352 940 7404
rect 992 7352 998 7404
rect 1210 7352 1216 7404
rect 1268 7352 1274 7404
rect 2130 7352 2136 7404
rect 2188 7392 2194 7404
rect 2314 7392 2320 7404
rect 2188 7364 2320 7392
rect 2188 7352 2194 7364
rect 2314 7352 2320 7364
rect 2372 7392 2378 7404
rect 4985 7395 5043 7401
rect 2372 7378 3634 7392
rect 2372 7364 3648 7378
rect 2372 7352 2378 7364
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 2777 7327 2835 7333
rect 2777 7324 2789 7327
rect 2464 7296 2789 7324
rect 2464 7284 2470 7296
rect 2777 7293 2789 7296
rect 2823 7293 2835 7327
rect 3620 7324 3648 7364
rect 4985 7361 4997 7395
rect 5031 7392 5043 7395
rect 5074 7392 5080 7404
rect 5031 7364 5080 7392
rect 5031 7361 5043 7364
rect 4985 7355 5043 7361
rect 4706 7324 4712 7336
rect 3620 7296 4712 7324
rect 2777 7287 2835 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 3970 7148 3976 7200
rect 4028 7188 4034 7200
rect 5000 7188 5028 7355
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 5626 7392 5632 7404
rect 5587 7364 5632 7392
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 8018 7352 8024 7404
rect 8076 7352 8082 7404
rect 8110 7352 8116 7404
rect 8168 7392 8174 7404
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8168 7364 8953 7392
rect 8168 7352 8174 7364
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 5997 7327 6055 7333
rect 5997 7293 6009 7327
rect 6043 7324 6055 7327
rect 6181 7327 6239 7333
rect 6181 7324 6193 7327
rect 6043 7296 6193 7324
rect 6043 7293 6055 7296
rect 5997 7287 6055 7293
rect 6181 7293 6193 7296
rect 6227 7293 6239 7327
rect 6181 7287 6239 7293
rect 6270 7284 6276 7336
rect 6328 7324 6334 7336
rect 6549 7327 6607 7333
rect 6549 7324 6561 7327
rect 6328 7296 6561 7324
rect 6328 7284 6334 7296
rect 6549 7293 6561 7296
rect 6595 7293 6607 7327
rect 6549 7287 6607 7293
rect 4028 7160 5028 7188
rect 4028 7148 4034 7160
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 644 7098 9384 7120
rect 644 7046 2554 7098
rect 2606 7046 2618 7098
rect 2670 7046 2682 7098
rect 2734 7046 6554 7098
rect 6606 7046 6618 7098
rect 6670 7046 6682 7098
rect 6734 7046 9384 7098
rect 644 7024 9384 7046
rect 6178 6944 6184 6996
rect 6236 6984 6242 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 6236 6956 7297 6984
rect 6236 6944 6242 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 5868 6888 7972 6916
rect 5868 6876 5874 6888
rect 4890 6808 4896 6860
rect 4948 6808 4954 6860
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4387 6752 4537 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7708 6752 7849 6780
rect 7708 6740 7714 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7944 6780 7972 6888
rect 8570 6780 8576 6792
rect 7944 6752 8576 6780
rect 7837 6743 7895 6749
rect 8570 6740 8576 6752
rect 8628 6780 8634 6792
rect 8695 6783 8753 6789
rect 8695 6780 8707 6783
rect 8628 6752 8707 6780
rect 8628 6740 8634 6752
rect 8695 6749 8707 6752
rect 8741 6749 8753 6783
rect 8695 6743 8753 6749
rect 8846 6740 8852 6792
rect 8904 6740 8910 6792
rect 5534 6672 5540 6724
rect 5592 6672 5598 6724
rect 6929 6715 6987 6721
rect 6929 6681 6941 6715
rect 6975 6712 6987 6715
rect 8110 6712 8116 6724
rect 6975 6684 8116 6712
rect 6975 6681 6987 6684
rect 6929 6675 6987 6681
rect 8110 6672 8116 6684
rect 8168 6672 8174 6724
rect 8478 6604 8484 6656
rect 8536 6604 8542 6656
rect 644 6554 9384 6576
rect 644 6502 2954 6554
rect 3006 6502 3018 6554
rect 3070 6502 3082 6554
rect 3134 6502 6954 6554
rect 7006 6502 7018 6554
rect 7070 6502 7082 6554
rect 7134 6502 9384 6554
rect 644 6480 9384 6502
rect 1118 6400 1124 6452
rect 1176 6400 1182 6452
rect 3970 6400 3976 6452
rect 4028 6400 4034 6452
rect 4890 6440 4896 6452
rect 4172 6412 4896 6440
rect 3988 6372 4016 6400
rect 4172 6381 4200 6412
rect 4890 6400 4896 6412
rect 4948 6400 4954 6452
rect 5629 6443 5687 6449
rect 5629 6409 5641 6443
rect 5675 6440 5687 6443
rect 6086 6440 6092 6452
rect 5675 6412 6092 6440
rect 5675 6409 5687 6412
rect 5629 6403 5687 6409
rect 6086 6400 6092 6412
rect 6144 6400 6150 6452
rect 3896 6344 4016 6372
rect 4157 6375 4215 6381
rect 474 6264 480 6316
rect 532 6304 538 6316
rect 3896 6313 3924 6344
rect 4157 6341 4169 6375
rect 4203 6341 4215 6375
rect 8478 6372 8484 6384
rect 8050 6344 8484 6372
rect 4157 6335 4215 6341
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 937 6307 995 6313
rect 937 6304 949 6307
rect 532 6276 949 6304
rect 532 6264 538 6276
rect 937 6273 949 6276
rect 983 6273 995 6307
rect 937 6267 995 6273
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 5626 6264 5632 6316
rect 5684 6304 5690 6316
rect 5810 6304 5816 6316
rect 5684 6276 5816 6304
rect 5684 6264 5690 6276
rect 5810 6264 5816 6276
rect 5868 6304 5874 6316
rect 5997 6307 6055 6313
rect 5997 6304 6009 6307
rect 5868 6276 6009 6304
rect 5868 6264 5874 6276
rect 5997 6273 6009 6276
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6273 6331 6307
rect 6273 6267 6331 6273
rect 4246 6196 4252 6248
rect 4304 6236 4310 6248
rect 5902 6236 5908 6248
rect 4304 6208 5908 6236
rect 4304 6196 4310 6208
rect 5902 6196 5908 6208
rect 5960 6236 5966 6248
rect 6288 6236 6316 6267
rect 6454 6264 6460 6316
rect 6512 6304 6518 6316
rect 6917 6307 6975 6313
rect 6917 6304 6929 6307
rect 6512 6276 6929 6304
rect 6512 6264 6518 6276
rect 6917 6273 6929 6276
rect 6963 6273 6975 6307
rect 6917 6267 6975 6273
rect 5960 6208 6316 6236
rect 6365 6239 6423 6245
rect 5960 6196 5966 6208
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 6411 6208 6561 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6932 6236 6960 6267
rect 8386 6264 8392 6316
rect 8444 6264 8450 6316
rect 7190 6236 7196 6248
rect 6932 6208 7196 6236
rect 6549 6199 6607 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6178 6100 6184 6112
rect 5776 6072 6184 6100
rect 5776 6060 5782 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8949 6103 9007 6109
rect 8949 6100 8961 6103
rect 8352 6072 8961 6100
rect 8352 6060 8358 6072
rect 8949 6069 8961 6072
rect 8995 6069 9007 6103
rect 8949 6063 9007 6069
rect 644 6010 9384 6032
rect 644 5958 2554 6010
rect 2606 5958 2618 6010
rect 2670 5958 2682 6010
rect 2734 5958 6554 6010
rect 6606 5958 6618 6010
rect 6670 5958 6682 6010
rect 6734 5958 9384 6010
rect 644 5936 9384 5958
rect 6549 5899 6607 5905
rect 6549 5865 6561 5899
rect 6595 5896 6607 5899
rect 6822 5896 6828 5908
rect 6595 5868 6828 5896
rect 6595 5865 6607 5868
rect 6549 5859 6607 5865
rect 6822 5856 6828 5868
rect 6880 5856 6886 5908
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 8444 5868 8493 5896
rect 8444 5856 8450 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 6362 5788 6368 5840
rect 6420 5828 6426 5840
rect 6641 5831 6699 5837
rect 6641 5828 6653 5831
rect 6420 5800 6653 5828
rect 6420 5788 6426 5800
rect 6641 5797 6653 5800
rect 6687 5797 6699 5831
rect 6641 5791 6699 5797
rect 382 5720 388 5772
rect 440 5760 446 5772
rect 1397 5763 1455 5769
rect 1397 5760 1409 5763
rect 440 5732 1409 5760
rect 440 5720 446 5732
rect 1397 5729 1409 5732
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 3970 5720 3976 5772
rect 4028 5760 4034 5772
rect 5077 5763 5135 5769
rect 4028 5732 4154 5760
rect 4028 5720 4034 5732
rect 1118 5652 1124 5704
rect 1176 5652 1182 5704
rect 4126 5692 4154 5732
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 6270 5760 6276 5772
rect 5123 5732 6276 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 9582 5760 9588 5772
rect 7883 5732 9588 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 4798 5692 4804 5704
rect 4126 5664 4804 5692
rect 4798 5652 4804 5664
rect 4856 5652 4862 5704
rect 6178 5652 6184 5704
rect 6236 5652 6242 5704
rect 6825 5695 6883 5701
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 8202 5692 8208 5704
rect 6871 5664 8208 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 8202 5652 8208 5664
rect 8260 5652 8266 5704
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8662 5652 8668 5704
rect 8720 5652 8726 5704
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 8849 5627 8907 5633
rect 8849 5624 8861 5627
rect 8628 5596 8861 5624
rect 8628 5584 8634 5596
rect 8849 5593 8861 5596
rect 8895 5593 8907 5627
rect 8849 5587 8907 5593
rect 644 5466 9384 5488
rect 644 5414 2954 5466
rect 3006 5414 3018 5466
rect 3070 5414 3082 5466
rect 3134 5414 6954 5466
rect 7006 5414 7018 5466
rect 7070 5414 7082 5466
rect 7134 5414 9384 5466
rect 644 5392 9384 5414
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 5994 5352 6000 5364
rect 5767 5324 6000 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 5442 5244 5448 5296
rect 5500 5284 5506 5296
rect 5500 5256 7696 5284
rect 5500 5244 5506 5256
rect 2314 5176 2320 5228
rect 2372 5176 2378 5228
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 7668 5225 7696 5256
rect 8846 5244 8852 5296
rect 8904 5244 8910 5296
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 934 5108 940 5160
rect 992 5108 998 5160
rect 1210 5108 1216 5160
rect 1268 5108 1274 5160
rect 2406 5108 2412 5160
rect 2464 5148 2470 5160
rect 2685 5151 2743 5157
rect 2685 5148 2697 5151
rect 2464 5120 2697 5148
rect 2464 5108 2470 5120
rect 2685 5117 2697 5120
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 5074 5108 5080 5160
rect 5132 5108 5138 5160
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 9582 5148 9588 5160
rect 7423 5120 9588 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 644 4922 9384 4944
rect 644 4870 2554 4922
rect 2606 4870 2618 4922
rect 2670 4870 2682 4922
rect 2734 4870 6554 4922
rect 6606 4870 6618 4922
rect 6670 4870 6682 4922
rect 6734 4870 9384 4922
rect 644 4848 9384 4870
rect 1118 4768 1124 4820
rect 1176 4768 1182 4820
rect 4982 4768 4988 4820
rect 5040 4808 5046 4820
rect 5040 4780 8432 4808
rect 5040 4768 5046 4780
rect 2133 4743 2191 4749
rect 2133 4709 2145 4743
rect 2179 4740 2191 4743
rect 2314 4740 2320 4752
rect 2179 4712 2320 4740
rect 2179 4709 2191 4712
rect 2133 4703 2191 4709
rect 2314 4700 2320 4712
rect 2372 4700 2378 4752
rect 4893 4743 4951 4749
rect 4893 4740 4905 4743
rect 4264 4712 4905 4740
rect 1489 4675 1547 4681
rect 1489 4641 1501 4675
rect 1535 4672 1547 4675
rect 2774 4672 2780 4684
rect 1535 4644 2780 4672
rect 1535 4641 1547 4644
rect 1489 4635 1547 4641
rect 2774 4632 2780 4644
rect 2832 4632 2838 4684
rect 4264 4681 4292 4712
rect 4893 4709 4905 4712
rect 4939 4709 4951 4743
rect 4893 4703 4951 4709
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4641 4307 4675
rect 4249 4635 4307 4641
rect 4798 4632 4804 4684
rect 4856 4672 4862 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 4856 4644 6653 4672
rect 4856 4632 4862 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4672 7895 4675
rect 8202 4672 8208 4684
rect 7883 4644 8208 4672
rect 7883 4641 7895 4644
rect 7837 4635 7895 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 1302 4564 1308 4616
rect 1360 4564 1366 4616
rect 1854 4564 1860 4616
rect 1912 4604 1918 4616
rect 1949 4607 2007 4613
rect 1949 4604 1961 4607
rect 1912 4576 1961 4604
rect 1912 4564 1918 4576
rect 1949 4573 1961 4576
rect 1995 4573 2007 4607
rect 1949 4567 2007 4573
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 8404 4604 8432 4780
rect 9030 4672 9036 4684
rect 8680 4644 9036 4672
rect 8680 4613 8708 4644
rect 9030 4632 9036 4644
rect 9088 4632 9094 4684
rect 8680 4607 8753 4613
rect 8680 4604 8707 4607
rect 8404 4576 8707 4604
rect 8695 4573 8707 4576
rect 8741 4573 8753 4607
rect 8695 4567 8753 4573
rect 8849 4607 8907 4613
rect 8849 4573 8861 4607
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 6086 4496 6092 4548
rect 6144 4536 6150 4548
rect 6365 4539 6423 4545
rect 6365 4536 6377 4539
rect 6144 4508 6377 4536
rect 6144 4496 6150 4508
rect 6365 4505 6377 4508
rect 6411 4505 6423 4539
rect 6365 4499 6423 4505
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 8864 4536 8892 4567
rect 8628 4508 8892 4536
rect 8628 4496 8634 4508
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 4801 4471 4859 4477
rect 4801 4468 4813 4471
rect 4764 4440 4813 4468
rect 4764 4428 4770 4440
rect 4801 4437 4813 4440
rect 4847 4437 4859 4471
rect 4801 4431 4859 4437
rect 8478 4428 8484 4480
rect 8536 4428 8542 4480
rect 644 4378 9384 4400
rect 644 4326 2954 4378
rect 3006 4326 3018 4378
rect 3070 4326 3082 4378
rect 3134 4326 6954 4378
rect 7006 4326 7018 4378
rect 7070 4326 7082 4378
rect 7134 4326 9384 4378
rect 644 4304 9384 4326
rect 934 4224 940 4276
rect 992 4264 998 4276
rect 4154 4264 4160 4276
rect 992 4236 4160 4264
rect 992 4224 998 4236
rect 474 4088 480 4140
rect 532 4128 538 4140
rect 3804 4137 3832 4236
rect 4154 4224 4160 4236
rect 4212 4264 4218 4276
rect 4798 4264 4804 4276
rect 4212 4236 4804 4264
rect 4212 4224 4218 4236
rect 4798 4224 4804 4236
rect 4856 4224 4862 4276
rect 5534 4224 5540 4276
rect 5592 4224 5598 4276
rect 6086 4224 6092 4276
rect 6144 4264 6150 4276
rect 6273 4267 6331 4273
rect 6273 4264 6285 4267
rect 6144 4236 6285 4264
rect 6144 4224 6150 4236
rect 6273 4233 6285 4236
rect 6319 4233 6331 4267
rect 6273 4227 6331 4233
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8949 4267 9007 4273
rect 8949 4264 8961 4267
rect 8352 4236 8961 4264
rect 8352 4224 8358 4236
rect 8949 4233 8961 4236
rect 8995 4233 9007 4267
rect 8949 4227 9007 4233
rect 8478 4196 8484 4208
rect 8050 4168 8484 4196
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 937 4131 995 4137
rect 937 4128 949 4131
rect 532 4100 949 4128
rect 532 4088 538 4100
rect 937 4097 949 4100
rect 983 4097 995 4131
rect 937 4091 995 4097
rect 3789 4131 3847 4137
rect 3789 4097 3801 4131
rect 3835 4097 3847 4131
rect 3789 4091 3847 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 6052 4100 6101 4128
rect 6052 4088 6058 4100
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6089 4091 6147 4097
rect 6196 4100 6929 4128
rect 4798 4020 4804 4072
rect 4856 4060 4862 4072
rect 5258 4060 5264 4072
rect 4856 4032 5264 4060
rect 4856 4020 4862 4032
rect 5258 4020 5264 4032
rect 5316 4060 5322 4072
rect 6196 4060 6224 4100
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 5316 4032 6224 4060
rect 6549 4063 6607 4069
rect 5316 4020 5322 4032
rect 6549 4029 6561 4063
rect 6595 4060 6607 4063
rect 6822 4060 6828 4072
rect 6595 4032 6828 4060
rect 6595 4029 6607 4032
rect 6549 4023 6607 4029
rect 6822 4020 6828 4032
rect 6880 4020 6886 4072
rect 1121 3995 1179 4001
rect 1121 3961 1133 3995
rect 1167 3992 1179 3995
rect 1210 3992 1216 4004
rect 1167 3964 1216 3992
rect 1167 3961 1179 3964
rect 1121 3955 1179 3961
rect 1210 3952 1216 3964
rect 1268 3952 1274 4004
rect 5166 3952 5172 4004
rect 5224 3992 5230 4004
rect 6086 3992 6092 4004
rect 5224 3964 6092 3992
rect 5224 3952 5230 3964
rect 6086 3952 6092 3964
rect 6144 3952 6150 4004
rect 6196 3964 6408 3992
rect 4052 3927 4110 3933
rect 4052 3893 4064 3927
rect 4098 3924 4110 3927
rect 6196 3924 6224 3964
rect 4098 3896 6224 3924
rect 6380 3924 6408 3964
rect 7190 3924 7196 3936
rect 6380 3896 7196 3924
rect 4098 3893 4110 3896
rect 4052 3887 4110 3893
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 644 3834 9384 3856
rect 644 3782 6554 3834
rect 6606 3782 6618 3834
rect 6670 3782 6682 3834
rect 6734 3782 9384 3834
rect 644 3760 9384 3782
rect 3973 3723 4031 3729
rect 3973 3689 3985 3723
rect 4019 3720 4031 3723
rect 5074 3720 5080 3732
rect 4019 3692 5080 3720
rect 4019 3689 4031 3692
rect 3973 3683 4031 3689
rect 5074 3680 5080 3692
rect 5132 3680 5138 3732
rect 6822 3680 6828 3732
rect 6880 3720 6886 3732
rect 7837 3723 7895 3729
rect 7837 3720 7849 3723
rect 6880 3692 7849 3720
rect 6880 3680 6886 3692
rect 7837 3689 7849 3692
rect 7883 3689 7895 3723
rect 7837 3683 7895 3689
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8444 3692 8493 3720
rect 8444 3680 8450 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 7650 3612 7656 3664
rect 7708 3612 7714 3664
rect 4154 3544 4160 3596
rect 4212 3584 4218 3596
rect 4798 3584 4804 3596
rect 4212 3556 4804 3584
rect 4212 3544 4218 3556
rect 4798 3544 4804 3556
rect 4856 3584 4862 3596
rect 5721 3587 5779 3593
rect 5721 3584 5733 3587
rect 4856 3556 5733 3584
rect 4856 3544 4862 3556
rect 5721 3553 5733 3556
rect 5767 3584 5779 3587
rect 5905 3587 5963 3593
rect 5905 3584 5917 3587
rect 5767 3556 5917 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 5905 3553 5917 3556
rect 5951 3553 5963 3587
rect 5905 3547 5963 3553
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 7190 3584 7196 3596
rect 6227 3556 7196 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3516 7987 3519
rect 8018 3516 8024 3528
rect 7975 3488 8024 3516
rect 7975 3485 7987 3488
rect 7929 3479 7987 3485
rect 8018 3476 8024 3488
rect 8076 3476 8082 3528
rect 8849 3519 8907 3525
rect 8849 3485 8861 3519
rect 8895 3516 8907 3519
rect 9030 3516 9036 3528
rect 8895 3488 9036 3516
rect 8895 3485 8907 3488
rect 8849 3479 8907 3485
rect 9030 3476 9036 3488
rect 9088 3476 9094 3528
rect 5166 3448 5172 3460
rect 5014 3420 5172 3448
rect 5166 3408 5172 3420
rect 5224 3408 5230 3460
rect 5442 3408 5448 3460
rect 5500 3408 5506 3460
rect 6086 3408 6092 3460
rect 6144 3448 6150 3460
rect 6270 3448 6276 3460
rect 6144 3420 6276 3448
rect 6144 3408 6150 3420
rect 6270 3408 6276 3420
rect 6328 3448 6334 3460
rect 8665 3451 8723 3457
rect 6328 3420 6670 3448
rect 6328 3408 6334 3420
rect 6564 3380 6592 3420
rect 8665 3417 8677 3451
rect 8711 3417 8723 3451
rect 8665 3411 8723 3417
rect 8570 3380 8576 3392
rect 6564 3352 8576 3380
rect 8570 3340 8576 3352
rect 8628 3380 8634 3392
rect 8680 3380 8708 3411
rect 8628 3352 8708 3380
rect 8628 3340 8634 3352
rect 644 3290 9384 3312
rect 644 3238 6954 3290
rect 7006 3238 7018 3290
rect 7070 3238 7082 3290
rect 7134 3238 9384 3290
rect 644 3216 9384 3238
rect 9030 3176 9036 3188
rect 5736 3148 9036 3176
rect 5736 3049 5764 3148
rect 9030 3136 9036 3148
rect 9088 3136 9094 3188
rect 6822 3068 6828 3120
rect 6880 3068 6886 3120
rect 8570 3068 8576 3120
rect 8628 3108 8634 3120
rect 8665 3111 8723 3117
rect 8665 3108 8677 3111
rect 8628 3080 8677 3108
rect 8628 3068 8634 3080
rect 8665 3077 8677 3080
rect 8711 3077 8723 3111
rect 8665 3071 8723 3077
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5156 3043 5214 3049
rect 5156 3040 5168 3043
rect 5031 3012 5168 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5156 3009 5168 3012
rect 5202 3009 5214 3043
rect 5156 3003 5214 3009
rect 5721 3043 5779 3049
rect 5721 3009 5733 3043
rect 5767 3009 5779 3043
rect 5721 3003 5779 3009
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7745 3043 7803 3049
rect 7745 3040 7757 3043
rect 7248 3012 7757 3040
rect 7248 3000 7254 3012
rect 7745 3009 7757 3012
rect 7791 3009 7803 3043
rect 8481 3043 8539 3049
rect 8481 3040 8493 3043
rect 7745 3003 7803 3009
rect 7852 3012 8493 3040
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2972 4583 2975
rect 5626 2972 5632 2984
rect 4571 2944 5632 2972
rect 4571 2941 4583 2944
rect 4525 2935 4583 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2972 7619 2975
rect 7650 2972 7656 2984
rect 7607 2944 7656 2972
rect 7607 2941 7619 2944
rect 7561 2935 7619 2941
rect 7650 2932 7656 2944
rect 7708 2932 7714 2984
rect 6454 2796 6460 2848
rect 6512 2836 6518 2848
rect 7852 2836 7880 3012
rect 8481 3009 8493 3012
rect 8527 3009 8539 3043
rect 8481 3003 8539 3009
rect 8294 2932 8300 2984
rect 8352 2932 8358 2984
rect 6512 2808 7880 2836
rect 6512 2796 6518 2808
rect 8110 2796 8116 2848
rect 8168 2836 8174 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 8168 2808 8861 2836
rect 8168 2796 8174 2808
rect 8849 2805 8861 2808
rect 8895 2805 8907 2839
rect 8849 2799 8907 2805
rect 2484 2746 9384 2768
rect 2484 2694 6554 2746
rect 6606 2694 6618 2746
rect 6670 2694 6682 2746
rect 6734 2694 9384 2746
rect 2484 2672 9384 2694
rect 2222 2592 2228 2644
rect 2280 2632 2286 2644
rect 2777 2635 2835 2641
rect 2777 2632 2789 2635
rect 2280 2604 2789 2632
rect 2280 2592 2286 2604
rect 2777 2601 2789 2604
rect 2823 2601 2835 2635
rect 2777 2595 2835 2601
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 5500 2604 5825 2632
rect 5500 2592 5506 2604
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 5813 2595 5871 2601
rect 5828 2564 5856 2595
rect 6822 2592 6828 2644
rect 6880 2632 6886 2644
rect 8757 2635 8815 2641
rect 8757 2632 8769 2635
rect 6880 2604 8769 2632
rect 6880 2592 6886 2604
rect 8757 2601 8769 2604
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 5828 2536 6132 2564
rect 1302 2456 1308 2508
rect 1360 2496 1366 2508
rect 4893 2499 4951 2505
rect 1360 2468 3188 2496
rect 1360 2456 1366 2468
rect 3160 2440 3188 2468
rect 4893 2465 4905 2499
rect 4939 2496 4951 2499
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 4939 2468 6009 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 6104 2496 6132 2536
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 6104 2468 6377 2496
rect 5997 2459 6055 2465
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 2961 2431 3019 2437
rect 2961 2428 2973 2431
rect 1872 2400 2973 2428
rect 1872 1544 1900 2400
rect 2961 2397 2973 2400
rect 3007 2397 3019 2431
rect 2961 2391 3019 2397
rect 3142 2388 3148 2440
rect 3200 2388 3206 2440
rect 4706 2388 4712 2440
rect 4764 2428 4770 2440
rect 4801 2431 4859 2437
rect 4801 2428 4813 2431
rect 4764 2400 4813 2428
rect 4764 2388 4770 2400
rect 4801 2397 4813 2400
rect 4847 2397 4859 2431
rect 4801 2391 4859 2397
rect 5261 2431 5319 2437
rect 5261 2397 5273 2431
rect 5307 2428 5319 2431
rect 5534 2428 5540 2440
rect 5307 2400 5540 2428
rect 5307 2397 5319 2400
rect 5261 2391 5319 2397
rect 4816 2360 4844 2391
rect 5534 2388 5540 2400
rect 5592 2388 5598 2440
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8110 2428 8116 2440
rect 7883 2400 8116 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8110 2388 8116 2400
rect 8168 2388 8174 2440
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 8662 2388 8668 2440
rect 8720 2428 8726 2440
rect 8720 2400 8765 2428
rect 8720 2388 8726 2400
rect 4816 2332 6040 2360
rect 6012 2292 6040 2332
rect 6822 2320 6828 2372
rect 6880 2320 6886 2372
rect 8018 2292 8024 2304
rect 6012 2264 8024 2292
rect 8018 2252 8024 2264
rect 8076 2252 8082 2304
rect 8110 2252 8116 2304
rect 8168 2292 8174 2304
rect 8397 2295 8455 2301
rect 8397 2292 8409 2295
rect 8168 2264 8409 2292
rect 8168 2252 8174 2264
rect 8397 2261 8409 2264
rect 8443 2261 8455 2295
rect 8397 2255 8455 2261
rect 2484 2202 9384 2224
rect 2484 2150 6954 2202
rect 7006 2150 7018 2202
rect 7070 2150 7082 2202
rect 7134 2150 9384 2202
rect 2484 2128 9384 2150
rect 7377 2091 7435 2097
rect 4724 2060 7052 2088
rect 4724 1961 4752 2060
rect 5169 2023 5227 2029
rect 5169 1989 5181 2023
rect 5215 2020 5227 2023
rect 5258 2020 5264 2032
rect 5215 1992 5264 2020
rect 5215 1989 5227 1992
rect 5169 1983 5227 1989
rect 5258 1980 5264 1992
rect 5316 1980 5322 2032
rect 6454 1980 6460 2032
rect 6512 2020 6518 2032
rect 7024 2020 7052 2060
rect 7377 2057 7389 2091
rect 7423 2088 7435 2091
rect 7650 2088 7656 2100
rect 7423 2060 7656 2088
rect 7423 2057 7435 2060
rect 7377 2051 7435 2057
rect 7650 2048 7656 2060
rect 7708 2048 7714 2100
rect 9030 2048 9036 2100
rect 9088 2048 9094 2100
rect 8110 2020 8116 2032
rect 6512 1992 6960 2020
rect 7024 1992 8116 2020
rect 6512 1980 6518 1992
rect 4709 1955 4767 1961
rect 4709 1921 4721 1955
rect 4755 1921 4767 1955
rect 4709 1915 4767 1921
rect 4798 1912 4804 1964
rect 4856 1952 4862 1964
rect 4893 1955 4951 1961
rect 4893 1952 4905 1955
rect 4856 1924 4905 1952
rect 4856 1912 4862 1924
rect 4893 1921 4905 1924
rect 4939 1921 4951 1955
rect 4893 1915 4951 1921
rect 6270 1912 6276 1964
rect 6328 1952 6334 1964
rect 6932 1961 6960 1992
rect 8110 1980 8116 1992
rect 8168 1980 8174 2032
rect 8570 1980 8576 2032
rect 8628 2020 8634 2032
rect 8849 2023 8907 2029
rect 8849 2020 8861 2023
rect 8628 1992 8861 2020
rect 8628 1980 8634 1992
rect 8849 1989 8861 1992
rect 8895 1989 8907 2023
rect 8849 1983 8907 1989
rect 6825 1955 6883 1961
rect 6825 1952 6837 1955
rect 6328 1924 6837 1952
rect 6328 1912 6334 1924
rect 6825 1921 6837 1924
rect 6871 1921 6883 1955
rect 6825 1915 6883 1921
rect 6918 1955 6976 1961
rect 6918 1921 6930 1955
rect 6964 1921 6976 1955
rect 6918 1915 6976 1921
rect 7469 1955 7527 1961
rect 7469 1921 7481 1955
rect 7515 1952 7527 1955
rect 8018 1952 8024 1964
rect 7515 1924 8024 1952
rect 7515 1921 7527 1924
rect 7469 1915 7527 1921
rect 8018 1912 8024 1924
rect 8076 1912 8082 1964
rect 8662 1912 8668 1964
rect 8720 1912 8726 1964
rect 4341 1887 4399 1893
rect 4341 1853 4353 1887
rect 4387 1884 4399 1887
rect 9582 1884 9588 1896
rect 4387 1856 9588 1884
rect 4387 1853 4399 1856
rect 4341 1847 4399 1853
rect 9582 1844 9588 1856
rect 9640 1844 9646 1896
rect 6641 1819 6699 1825
rect 6641 1785 6653 1819
rect 6687 1816 6699 1819
rect 8294 1816 8300 1828
rect 6687 1788 8300 1816
rect 6687 1785 6699 1788
rect 6641 1779 6699 1785
rect 8294 1776 8300 1788
rect 8352 1776 8358 1828
rect 2866 1708 2872 1760
rect 2924 1748 2930 1760
rect 6454 1748 6460 1760
rect 2924 1720 6460 1748
rect 2924 1708 2930 1720
rect 6454 1708 6460 1720
rect 6512 1708 6518 1760
rect 6822 1708 6828 1760
rect 6880 1748 6886 1760
rect 7009 1751 7067 1757
rect 7009 1748 7021 1751
rect 6880 1720 7021 1748
rect 6880 1708 6886 1720
rect 7009 1717 7021 1720
rect 7055 1717 7067 1751
rect 7009 1711 7067 1717
rect 2484 1658 9384 1680
rect 2484 1606 6554 1658
rect 6606 1606 6618 1658
rect 6670 1606 6682 1658
rect 6734 1606 9384 1658
rect 2484 1584 9384 1606
rect 1702 1516 1900 1544
rect 3142 1504 3148 1556
rect 3200 1544 3206 1556
rect 8849 1547 8907 1553
rect 8849 1544 8861 1547
rect 3200 1516 8861 1544
rect 3200 1504 3206 1516
rect 8849 1513 8861 1516
rect 8895 1513 8907 1547
rect 8849 1507 8907 1513
rect 6454 1436 6460 1488
rect 6512 1476 6518 1488
rect 8662 1476 8668 1488
rect 6512 1448 8668 1476
rect 6512 1436 6518 1448
rect 8662 1436 8668 1448
rect 8720 1436 8726 1488
rect 7377 1411 7435 1417
rect 7377 1377 7389 1411
rect 7423 1408 7435 1411
rect 8386 1408 8392 1420
rect 7423 1380 8392 1408
rect 7423 1377 7435 1380
rect 7377 1371 7435 1377
rect 8386 1368 8392 1380
rect 8444 1368 8450 1420
rect 6365 1343 6423 1349
rect 6365 1309 6377 1343
rect 6411 1340 6423 1343
rect 8202 1340 8208 1352
rect 6411 1312 8208 1340
rect 6411 1309 6423 1312
rect 6365 1303 6423 1309
rect 8202 1300 8208 1312
rect 8260 1300 8266 1352
rect 9030 1300 9036 1352
rect 9088 1300 9094 1352
rect 2484 1114 9384 1136
rect 2484 1062 6954 1114
rect 7006 1062 7018 1114
rect 7070 1062 7082 1114
rect 7134 1062 9384 1114
rect 2484 1040 9384 1062
<< via1 >>
rect 3608 14424 3660 14476
rect 5724 14424 5776 14476
rect 3240 14356 3292 14408
rect 8208 14356 8260 14408
rect 4620 14288 4672 14340
rect 7104 14288 7156 14340
rect 1124 14220 1176 14272
rect 6276 14220 6328 14272
rect 6368 14220 6420 14272
rect 6828 14220 6880 14272
rect 2954 14118 3006 14170
rect 3018 14118 3070 14170
rect 3082 14118 3134 14170
rect 6954 14118 7006 14170
rect 7018 14118 7070 14170
rect 7082 14118 7134 14170
rect 4804 14016 4856 14068
rect 4160 13948 4212 14000
rect 7656 14016 7708 14068
rect 3976 13880 4028 13932
rect 9588 13948 9640 14000
rect 4712 13880 4764 13932
rect 7656 13880 7708 13932
rect 8576 13880 8628 13932
rect 3240 13812 3292 13864
rect 5172 13744 5224 13796
rect 6368 13744 6420 13796
rect 8484 13812 8536 13864
rect 8852 13923 8904 13932
rect 8852 13889 8861 13923
rect 8861 13889 8895 13923
rect 8895 13889 8904 13923
rect 8852 13880 8904 13889
rect 9220 13812 9272 13864
rect 8024 13744 8076 13796
rect 2320 13676 2372 13728
rect 2780 13676 2832 13728
rect 4068 13676 4120 13728
rect 4988 13676 5040 13728
rect 6184 13676 6236 13728
rect 8116 13676 8168 13728
rect 2554 13574 2606 13626
rect 2618 13574 2670 13626
rect 2682 13574 2734 13626
rect 6554 13574 6606 13626
rect 6618 13574 6670 13626
rect 6682 13574 6734 13626
rect 3976 13515 4028 13524
rect 3976 13481 3985 13515
rect 3985 13481 4019 13515
rect 4019 13481 4028 13515
rect 3976 13472 4028 13481
rect 6000 13472 6052 13524
rect 1124 13379 1176 13388
rect 1124 13345 1133 13379
rect 1133 13345 1167 13379
rect 1167 13345 1176 13379
rect 1124 13336 1176 13345
rect 4528 13404 4580 13456
rect 3608 13336 3660 13388
rect 4620 13379 4672 13388
rect 4620 13345 4629 13379
rect 4629 13345 4663 13379
rect 4663 13345 4672 13379
rect 4620 13336 4672 13345
rect 4436 13268 4488 13320
rect 2228 13200 2280 13252
rect 3608 13200 3660 13252
rect 5080 13200 5132 13252
rect 5356 13404 5408 13456
rect 9036 13472 9088 13524
rect 7196 13404 7248 13456
rect 9588 13336 9640 13388
rect 6828 13311 6880 13320
rect 6828 13277 6837 13311
rect 6837 13277 6871 13311
rect 6871 13277 6880 13311
rect 6828 13268 6880 13277
rect 5632 13200 5684 13252
rect 5908 13200 5960 13252
rect 9128 13268 9180 13320
rect 1584 13132 1636 13184
rect 1768 13132 1820 13184
rect 4252 13132 4304 13184
rect 8208 13132 8260 13184
rect 8760 13200 8812 13252
rect 9220 13132 9272 13184
rect 2954 13030 3006 13082
rect 3018 13030 3070 13082
rect 3082 13030 3134 13082
rect 6954 13030 7006 13082
rect 7018 13030 7070 13082
rect 7082 13030 7134 13082
rect 6460 12928 6512 12980
rect 4160 12860 4212 12912
rect 940 12835 992 12844
rect 940 12801 949 12835
rect 949 12801 983 12835
rect 983 12801 992 12835
rect 940 12792 992 12801
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 6276 12835 6328 12844
rect 6276 12801 6285 12835
rect 6285 12801 6319 12835
rect 6319 12801 6328 12835
rect 6276 12792 6328 12801
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 1492 12724 1544 12776
rect 3240 12767 3292 12776
rect 3240 12733 3249 12767
rect 3249 12733 3283 12767
rect 3283 12733 3292 12767
rect 3240 12724 3292 12733
rect 6000 12724 6052 12776
rect 2780 12588 2832 12640
rect 5816 12588 5868 12640
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 6828 12724 6880 12776
rect 8852 12588 8904 12640
rect 8944 12631 8996 12640
rect 8944 12597 8961 12631
rect 8961 12597 8995 12631
rect 8995 12597 8996 12631
rect 8944 12588 8996 12597
rect 2554 12486 2606 12538
rect 2618 12486 2670 12538
rect 2682 12486 2734 12538
rect 6554 12486 6606 12538
rect 6618 12486 6670 12538
rect 6682 12486 6734 12538
rect 3240 12384 3292 12436
rect 1492 12316 1544 12368
rect 4160 12316 4212 12368
rect 2136 12248 2188 12300
rect 1216 12180 1268 12232
rect 1400 12112 1452 12164
rect 6368 12384 6420 12436
rect 7656 12384 7708 12436
rect 7196 12316 7248 12368
rect 3608 12223 3660 12232
rect 3608 12189 3618 12223
rect 3618 12189 3652 12223
rect 3652 12189 3660 12223
rect 3608 12180 3660 12189
rect 4160 12180 4212 12232
rect 4712 12223 4764 12232
rect 4712 12189 4721 12223
rect 4721 12189 4755 12223
rect 4755 12189 4764 12223
rect 4712 12180 4764 12189
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 8116 12248 8168 12300
rect 7656 12180 7708 12232
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8668 12223 8720 12232
rect 8668 12189 8707 12223
rect 8707 12189 8720 12223
rect 8668 12180 8720 12189
rect 6092 12112 6144 12164
rect 9220 12180 9272 12232
rect 3608 12044 3660 12096
rect 4068 12044 4120 12096
rect 5540 12044 5592 12096
rect 7656 12044 7708 12096
rect 8116 12087 8168 12096
rect 8116 12053 8125 12087
rect 8125 12053 8159 12087
rect 8159 12053 8168 12087
rect 8116 12044 8168 12053
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 8760 12044 8812 12096
rect 2954 11942 3006 11994
rect 3018 11942 3070 11994
rect 3082 11942 3134 11994
rect 6954 11942 7006 11994
rect 7018 11942 7070 11994
rect 7082 11942 7134 11994
rect 940 11883 992 11892
rect 940 11849 949 11883
rect 949 11849 983 11883
rect 983 11849 992 11883
rect 940 11840 992 11849
rect 2412 11840 2464 11892
rect 5724 11840 5776 11892
rect 1400 11772 1452 11824
rect 2136 11772 2188 11824
rect 3608 11772 3660 11824
rect 5448 11772 5500 11824
rect 6276 11840 6328 11892
rect 5356 11704 5408 11756
rect 6184 11704 6236 11756
rect 8116 11840 8168 11892
rect 8576 11840 8628 11892
rect 8484 11772 8536 11824
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 2412 11679 2464 11688
rect 2412 11645 2421 11679
rect 2421 11645 2455 11679
rect 2455 11645 2464 11679
rect 2412 11636 2464 11645
rect 6092 11636 6144 11688
rect 2780 11568 2832 11620
rect 6276 11568 6328 11620
rect 4528 11500 4580 11552
rect 4804 11500 4856 11552
rect 5080 11500 5132 11552
rect 5908 11543 5960 11552
rect 5908 11509 5917 11543
rect 5917 11509 5951 11543
rect 5951 11509 5960 11543
rect 5908 11500 5960 11509
rect 2554 11398 2606 11450
rect 2618 11398 2670 11450
rect 2682 11398 2734 11450
rect 6554 11398 6606 11450
rect 6618 11398 6670 11450
rect 6682 11398 6734 11450
rect 2780 11296 2832 11348
rect 4712 11296 4764 11348
rect 6828 11339 6880 11348
rect 6828 11305 6837 11339
rect 6837 11305 6871 11339
rect 6871 11305 6880 11339
rect 6828 11296 6880 11305
rect 3240 11228 3292 11280
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2228 11092 2280 11144
rect 1032 11067 1084 11076
rect 1032 11033 1041 11067
rect 1041 11033 1075 11067
rect 1075 11033 1084 11067
rect 1032 11024 1084 11033
rect 1952 11024 2004 11076
rect 4160 11160 4212 11212
rect 5908 11160 5960 11212
rect 5724 11092 5776 11144
rect 4896 11024 4948 11076
rect 8116 11067 8168 11076
rect 8116 11033 8125 11067
rect 8125 11033 8159 11067
rect 8159 11033 8168 11067
rect 8116 11024 8168 11033
rect 8668 11067 8720 11076
rect 2780 10956 2832 11008
rect 5632 10956 5684 11008
rect 6828 10956 6880 11008
rect 8668 11033 8677 11067
rect 8677 11033 8711 11067
rect 8711 11033 8720 11067
rect 8668 11024 8720 11033
rect 8760 11024 8812 11076
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 2954 10854 3006 10906
rect 3018 10854 3070 10906
rect 3082 10854 3134 10906
rect 6954 10854 7006 10906
rect 7018 10854 7070 10906
rect 7082 10854 7134 10906
rect 4160 10752 4212 10804
rect 4896 10752 4948 10804
rect 388 10684 440 10736
rect 3608 10684 3660 10736
rect 1216 10412 1268 10464
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 2228 10591 2280 10600
rect 2228 10557 2237 10591
rect 2237 10557 2271 10591
rect 2271 10557 2280 10591
rect 2228 10548 2280 10557
rect 3240 10548 3292 10600
rect 6184 10752 6236 10804
rect 6460 10795 6512 10804
rect 6460 10761 6469 10795
rect 6469 10761 6503 10795
rect 6503 10761 6512 10795
rect 6460 10752 6512 10761
rect 6828 10752 6880 10804
rect 5632 10659 5684 10668
rect 5632 10625 5641 10659
rect 5641 10625 5675 10659
rect 5675 10625 5684 10659
rect 5632 10616 5684 10625
rect 5816 10616 5868 10668
rect 8208 10684 8260 10736
rect 6276 10659 6328 10668
rect 6276 10625 6289 10659
rect 6289 10625 6328 10659
rect 6276 10616 6328 10625
rect 8484 10616 8536 10668
rect 6460 10548 6512 10600
rect 6184 10480 6236 10532
rect 2780 10412 2832 10464
rect 4252 10412 4304 10464
rect 5172 10412 5224 10464
rect 9036 10480 9088 10532
rect 8392 10412 8444 10464
rect 2554 10310 2606 10362
rect 2618 10310 2670 10362
rect 2682 10310 2734 10362
rect 6554 10310 6606 10362
rect 6618 10310 6670 10362
rect 6682 10310 6734 10362
rect 1400 10208 1452 10260
rect 1676 10208 1728 10260
rect 2228 10208 2280 10260
rect 2780 10208 2832 10260
rect 3240 10140 3292 10192
rect 480 10072 532 10124
rect 2044 10072 2096 10124
rect 3608 10072 3660 10124
rect 2136 10004 2188 10056
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 6000 10208 6052 10260
rect 6460 10208 6512 10260
rect 5816 10183 5868 10192
rect 5816 10149 5825 10183
rect 5825 10149 5859 10183
rect 5859 10149 5868 10183
rect 5816 10140 5868 10149
rect 8208 10140 8260 10192
rect 5540 10072 5592 10124
rect 6460 10072 6512 10124
rect 9588 10072 9640 10124
rect 1860 9979 1912 9988
rect 1860 9945 1869 9979
rect 1869 9945 1903 9979
rect 1903 9945 1912 9979
rect 1860 9936 1912 9945
rect 5540 9936 5592 9988
rect 5632 9979 5684 9988
rect 5632 9945 5641 9979
rect 5641 9945 5675 9979
rect 5675 9945 5684 9979
rect 5632 9936 5684 9945
rect 5908 10047 5960 10056
rect 5908 10013 5917 10047
rect 5917 10013 5951 10047
rect 5951 10013 5960 10047
rect 5908 10004 5960 10013
rect 6000 9936 6052 9988
rect 8024 10004 8076 10056
rect 8392 10004 8444 10056
rect 8576 10004 8628 10056
rect 8760 10047 8812 10056
rect 8760 10013 8768 10047
rect 8768 10013 8802 10047
rect 8802 10013 8812 10047
rect 8760 10004 8812 10013
rect 2320 9868 2372 9920
rect 3240 9868 3292 9920
rect 6276 9868 6328 9920
rect 8024 9868 8076 9920
rect 8668 9868 8720 9920
rect 2954 9766 3006 9818
rect 3018 9766 3070 9818
rect 3082 9766 3134 9818
rect 6954 9766 7006 9818
rect 7018 9766 7070 9818
rect 7082 9766 7134 9818
rect 1952 9664 2004 9716
rect 1676 9596 1728 9648
rect 2780 9664 2832 9716
rect 4896 9664 4948 9716
rect 5724 9707 5776 9716
rect 5724 9673 5733 9707
rect 5733 9673 5767 9707
rect 5767 9673 5776 9707
rect 5724 9664 5776 9673
rect 1676 9460 1728 9512
rect 1952 9460 2004 9512
rect 2412 9392 2464 9444
rect 3976 9596 4028 9648
rect 4252 9639 4304 9648
rect 4252 9605 4261 9639
rect 4261 9605 4295 9639
rect 4295 9605 4304 9639
rect 4252 9596 4304 9605
rect 5816 9596 5868 9648
rect 7656 9596 7708 9648
rect 6000 9528 6052 9580
rect 8852 9528 8904 9580
rect 3240 9460 3292 9512
rect 4988 9460 5040 9512
rect 6460 9460 6512 9512
rect 2780 9324 2832 9376
rect 3240 9324 3292 9376
rect 8576 9392 8628 9444
rect 8208 9324 8260 9376
rect 2554 9222 2606 9274
rect 2618 9222 2670 9274
rect 2682 9222 2734 9274
rect 6554 9222 6606 9274
rect 6618 9222 6670 9274
rect 6682 9222 6734 9274
rect 4528 9120 4580 9172
rect 5908 9120 5960 9172
rect 7656 9163 7708 9172
rect 7656 9129 7665 9163
rect 7665 9129 7699 9163
rect 7699 9129 7708 9163
rect 7656 9120 7708 9129
rect 8300 9163 8352 9172
rect 8300 9129 8309 9163
rect 8309 9129 8343 9163
rect 8343 9129 8352 9163
rect 8300 9120 8352 9129
rect 8852 9163 8904 9172
rect 8852 9129 8861 9163
rect 8861 9129 8895 9163
rect 8895 9129 8904 9163
rect 8852 9120 8904 9129
rect 388 8984 440 9036
rect 2228 8959 2280 8968
rect 2228 8925 2237 8959
rect 2237 8925 2271 8959
rect 2271 8925 2280 8959
rect 2228 8916 2280 8925
rect 2412 8780 2464 8832
rect 4436 9052 4488 9104
rect 5080 8984 5132 9036
rect 2780 8780 2832 8832
rect 4068 8916 4120 8968
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 5172 8916 5224 8968
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 7196 8916 7248 8968
rect 4160 8848 4212 8900
rect 5816 8848 5868 8900
rect 6184 8848 6236 8900
rect 3608 8780 3660 8832
rect 4344 8780 4396 8832
rect 8024 8848 8076 8900
rect 8668 8959 8720 8968
rect 8668 8925 8677 8959
rect 8677 8925 8711 8959
rect 8711 8925 8720 8959
rect 8668 8916 8720 8925
rect 7656 8780 7708 8832
rect 2954 8678 3006 8730
rect 3018 8678 3070 8730
rect 3082 8678 3134 8730
rect 6954 8678 7006 8730
rect 7018 8678 7070 8730
rect 7082 8678 7134 8730
rect 3608 8576 3660 8628
rect 2412 8508 2464 8560
rect 3240 8508 3292 8560
rect 4344 8576 4396 8628
rect 7196 8576 7248 8628
rect 8484 8576 8536 8628
rect 1216 8440 1268 8492
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 4436 8508 4488 8560
rect 5724 8508 5776 8560
rect 6828 8508 6880 8560
rect 8668 8508 8720 8560
rect 5816 8440 5868 8492
rect 3608 8372 3660 8424
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 6828 8415 6880 8424
rect 6828 8381 6837 8415
rect 6837 8381 6871 8415
rect 6871 8381 6880 8415
rect 6828 8372 6880 8381
rect 9588 8372 9640 8424
rect 1584 8236 1636 8288
rect 6460 8304 6512 8356
rect 5632 8236 5684 8288
rect 7196 8236 7248 8288
rect 2554 8134 2606 8186
rect 2618 8134 2670 8186
rect 2682 8134 2734 8186
rect 6554 8134 6606 8186
rect 6618 8134 6670 8186
rect 6682 8134 6734 8186
rect 1400 8032 1452 8084
rect 2780 8032 2832 8084
rect 1768 7964 1820 8016
rect 2320 7964 2372 8016
rect 6368 7964 6420 8016
rect 2780 7896 2832 7948
rect 3608 7896 3660 7948
rect 8392 7896 8444 7948
rect 1124 7828 1176 7880
rect 2320 7828 2372 7880
rect 1400 7803 1452 7812
rect 1400 7769 1409 7803
rect 1409 7769 1443 7803
rect 1443 7769 1452 7803
rect 1400 7760 1452 7769
rect 3240 7828 3292 7880
rect 4712 7828 4764 7880
rect 5356 7828 5408 7880
rect 5540 7828 5592 7880
rect 5632 7871 5684 7880
rect 5632 7837 5641 7871
rect 5641 7837 5675 7871
rect 5675 7837 5684 7871
rect 5632 7828 5684 7837
rect 1308 7735 1360 7744
rect 1308 7701 1317 7735
rect 1317 7701 1351 7735
rect 1351 7701 1360 7735
rect 1308 7692 1360 7701
rect 1952 7692 2004 7744
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 6276 7828 6328 7880
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8668 7871 8720 7880
rect 8668 7837 8677 7871
rect 8677 7837 8711 7871
rect 8711 7837 8720 7871
rect 8668 7828 8720 7837
rect 4620 7692 4672 7744
rect 4896 7692 4948 7744
rect 5724 7692 5776 7744
rect 8116 7760 8168 7812
rect 6368 7692 6420 7744
rect 8024 7692 8076 7744
rect 2954 7590 3006 7642
rect 3018 7590 3070 7642
rect 3082 7590 3134 7642
rect 6954 7590 7006 7642
rect 7018 7590 7070 7642
rect 7082 7590 7134 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 1676 7488 1728 7540
rect 3240 7531 3292 7540
rect 3240 7497 3249 7531
rect 3249 7497 3283 7531
rect 3283 7497 3292 7531
rect 3240 7488 3292 7497
rect 8300 7488 8352 7540
rect 8760 7531 8812 7540
rect 8760 7497 8769 7531
rect 8769 7497 8803 7531
rect 8803 7497 8812 7531
rect 8760 7488 8812 7497
rect 1952 7420 2004 7472
rect 4804 7420 4856 7472
rect 7656 7420 7708 7472
rect 940 7395 992 7404
rect 940 7361 949 7395
rect 949 7361 983 7395
rect 983 7361 992 7395
rect 940 7352 992 7361
rect 1216 7395 1268 7404
rect 1216 7361 1225 7395
rect 1225 7361 1259 7395
rect 1259 7361 1268 7395
rect 1216 7352 1268 7361
rect 2136 7352 2188 7404
rect 2320 7352 2372 7404
rect 2412 7284 2464 7336
rect 4712 7284 4764 7336
rect 3976 7148 4028 7200
rect 5080 7352 5132 7404
rect 5632 7395 5684 7404
rect 5632 7361 5640 7395
rect 5640 7361 5674 7395
rect 5674 7361 5684 7395
rect 5632 7352 5684 7361
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 8024 7395 8076 7404
rect 8024 7361 8033 7395
rect 8033 7361 8067 7395
rect 8067 7361 8076 7395
rect 8024 7352 8076 7361
rect 8116 7352 8168 7404
rect 6276 7284 6328 7336
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 2554 7046 2606 7098
rect 2618 7046 2670 7098
rect 2682 7046 2734 7098
rect 6554 7046 6606 7098
rect 6618 7046 6670 7098
rect 6682 7046 6734 7098
rect 6184 6944 6236 6996
rect 5816 6876 5868 6928
rect 4896 6851 4948 6860
rect 4896 6817 4905 6851
rect 4905 6817 4939 6851
rect 4939 6817 4948 6851
rect 4896 6808 4948 6817
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 7656 6740 7708 6792
rect 8576 6740 8628 6792
rect 8852 6783 8904 6792
rect 8852 6749 8861 6783
rect 8861 6749 8895 6783
rect 8895 6749 8904 6783
rect 8852 6740 8904 6749
rect 5540 6672 5592 6724
rect 8116 6672 8168 6724
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 2954 6502 3006 6554
rect 3018 6502 3070 6554
rect 3082 6502 3134 6554
rect 6954 6502 7006 6554
rect 7018 6502 7070 6554
rect 7082 6502 7134 6554
rect 1124 6443 1176 6452
rect 1124 6409 1133 6443
rect 1133 6409 1167 6443
rect 1167 6409 1176 6443
rect 1124 6400 1176 6409
rect 3976 6400 4028 6452
rect 4896 6400 4948 6452
rect 6092 6400 6144 6452
rect 480 6264 532 6316
rect 8484 6332 8536 6384
rect 5264 6264 5316 6316
rect 5632 6264 5684 6316
rect 5816 6264 5868 6316
rect 4252 6196 4304 6248
rect 5908 6196 5960 6248
rect 6460 6264 6512 6316
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 7196 6196 7248 6248
rect 5724 6060 5776 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 8300 6060 8352 6112
rect 2554 5958 2606 6010
rect 2618 5958 2670 6010
rect 2682 5958 2734 6010
rect 6554 5958 6606 6010
rect 6618 5958 6670 6010
rect 6682 5958 6734 6010
rect 6828 5856 6880 5908
rect 8392 5856 8444 5908
rect 6368 5788 6420 5840
rect 388 5720 440 5772
rect 3976 5720 4028 5772
rect 1124 5695 1176 5704
rect 1124 5661 1133 5695
rect 1133 5661 1167 5695
rect 1167 5661 1176 5695
rect 1124 5652 1176 5661
rect 6276 5720 6328 5772
rect 9588 5720 9640 5772
rect 4804 5695 4856 5704
rect 4804 5661 4813 5695
rect 4813 5661 4847 5695
rect 4847 5661 4856 5695
rect 4804 5652 4856 5661
rect 6184 5652 6236 5704
rect 8208 5652 8260 5704
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 8668 5695 8720 5704
rect 8668 5661 8677 5695
rect 8677 5661 8711 5695
rect 8711 5661 8720 5695
rect 8668 5652 8720 5661
rect 8576 5584 8628 5636
rect 2954 5414 3006 5466
rect 3018 5414 3070 5466
rect 3082 5414 3134 5466
rect 6954 5414 7006 5466
rect 7018 5414 7070 5466
rect 7082 5414 7134 5466
rect 6000 5312 6052 5364
rect 5448 5244 5500 5296
rect 2320 5176 2372 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 8852 5287 8904 5296
rect 8852 5253 8861 5287
rect 8861 5253 8895 5287
rect 8895 5253 8904 5287
rect 8852 5244 8904 5253
rect 940 5151 992 5160
rect 940 5117 949 5151
rect 949 5117 983 5151
rect 983 5117 992 5151
rect 940 5108 992 5117
rect 1216 5151 1268 5160
rect 1216 5117 1225 5151
rect 1225 5117 1259 5151
rect 1259 5117 1268 5151
rect 1216 5108 1268 5117
rect 2412 5108 2464 5160
rect 5080 5151 5132 5160
rect 5080 5117 5089 5151
rect 5089 5117 5123 5151
rect 5123 5117 5132 5151
rect 5080 5108 5132 5117
rect 9588 5108 9640 5160
rect 2554 4870 2606 4922
rect 2618 4870 2670 4922
rect 2682 4870 2734 4922
rect 6554 4870 6606 4922
rect 6618 4870 6670 4922
rect 6682 4870 6734 4922
rect 1124 4811 1176 4820
rect 1124 4777 1133 4811
rect 1133 4777 1167 4811
rect 1167 4777 1176 4811
rect 1124 4768 1176 4777
rect 4988 4768 5040 4820
rect 2320 4700 2372 4752
rect 2780 4632 2832 4684
rect 4804 4632 4856 4684
rect 8208 4632 8260 4684
rect 1308 4607 1360 4616
rect 1308 4573 1317 4607
rect 1317 4573 1351 4607
rect 1351 4573 1360 4607
rect 1308 4564 1360 4573
rect 1860 4564 1912 4616
rect 5264 4564 5316 4616
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 9036 4632 9088 4684
rect 6092 4496 6144 4548
rect 8576 4496 8628 4548
rect 4712 4428 4764 4480
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 2954 4326 3006 4378
rect 3018 4326 3070 4378
rect 3082 4326 3134 4378
rect 6954 4326 7006 4378
rect 7018 4326 7070 4378
rect 7082 4326 7134 4378
rect 940 4224 992 4276
rect 480 4088 532 4140
rect 4160 4224 4212 4276
rect 4804 4224 4856 4276
rect 5540 4267 5592 4276
rect 5540 4233 5549 4267
rect 5549 4233 5583 4267
rect 5583 4233 5592 4267
rect 5540 4224 5592 4233
rect 6092 4224 6144 4276
rect 8300 4224 8352 4276
rect 8484 4156 8536 4208
rect 5172 4088 5224 4140
rect 6000 4088 6052 4140
rect 4804 4020 4856 4072
rect 5264 4020 5316 4072
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 6828 4020 6880 4072
rect 1216 3952 1268 4004
rect 5172 3952 5224 4004
rect 6092 3952 6144 4004
rect 7196 3884 7248 3936
rect 6554 3782 6606 3834
rect 6618 3782 6670 3834
rect 6682 3782 6734 3834
rect 5080 3680 5132 3732
rect 6828 3680 6880 3732
rect 8392 3680 8444 3732
rect 7656 3655 7708 3664
rect 7656 3621 7665 3655
rect 7665 3621 7699 3655
rect 7699 3621 7708 3655
rect 7656 3612 7708 3621
rect 4160 3544 4212 3596
rect 4804 3544 4856 3596
rect 7196 3544 7248 3596
rect 8024 3476 8076 3528
rect 9036 3476 9088 3528
rect 5172 3408 5224 3460
rect 5448 3451 5500 3460
rect 5448 3417 5457 3451
rect 5457 3417 5491 3451
rect 5491 3417 5500 3451
rect 5448 3408 5500 3417
rect 6092 3408 6144 3460
rect 6276 3408 6328 3460
rect 8576 3340 8628 3392
rect 6954 3238 7006 3290
rect 7018 3238 7070 3290
rect 7082 3238 7134 3290
rect 9036 3136 9088 3188
rect 6828 3068 6880 3120
rect 8576 3068 8628 3120
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 5632 2932 5684 2984
rect 7656 2932 7708 2984
rect 6460 2796 6512 2848
rect 8300 2975 8352 2984
rect 8300 2941 8309 2975
rect 8309 2941 8343 2975
rect 8343 2941 8352 2975
rect 8300 2932 8352 2941
rect 8116 2796 8168 2848
rect 6554 2694 6606 2746
rect 6618 2694 6670 2746
rect 6682 2694 6734 2746
rect 2228 2592 2280 2644
rect 5448 2592 5500 2644
rect 6828 2592 6880 2644
rect 1308 2456 1360 2508
rect 3148 2431 3200 2440
rect 3148 2397 3157 2431
rect 3157 2397 3191 2431
rect 3191 2397 3200 2431
rect 3148 2388 3200 2397
rect 4712 2388 4764 2440
rect 5540 2388 5592 2440
rect 8116 2388 8168 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 8668 2431 8720 2440
rect 8668 2397 8678 2431
rect 8678 2397 8712 2431
rect 8712 2397 8720 2431
rect 8668 2388 8720 2397
rect 6828 2320 6880 2372
rect 8024 2252 8076 2304
rect 8116 2252 8168 2304
rect 6954 2150 7006 2202
rect 7018 2150 7070 2202
rect 7082 2150 7134 2202
rect 5264 1980 5316 2032
rect 6460 1980 6512 2032
rect 7656 2048 7708 2100
rect 9036 2091 9088 2100
rect 9036 2057 9045 2091
rect 9045 2057 9079 2091
rect 9079 2057 9088 2091
rect 9036 2048 9088 2057
rect 4804 1912 4856 1964
rect 6276 1912 6328 1964
rect 8116 1980 8168 2032
rect 8576 1980 8628 2032
rect 8024 1912 8076 1964
rect 8668 1955 8720 1964
rect 8668 1921 8677 1955
rect 8677 1921 8711 1955
rect 8711 1921 8720 1955
rect 8668 1912 8720 1921
rect 9588 1844 9640 1896
rect 8300 1776 8352 1828
rect 2872 1708 2924 1760
rect 6460 1708 6512 1760
rect 6828 1708 6880 1760
rect 6554 1606 6606 1658
rect 6618 1606 6670 1658
rect 6682 1606 6734 1658
rect 3148 1504 3200 1556
rect 6460 1436 6512 1488
rect 8668 1436 8720 1488
rect 8392 1368 8444 1420
rect 8208 1300 8260 1352
rect 9036 1343 9088 1352
rect 9036 1309 9045 1343
rect 9045 1309 9079 1343
rect 9079 1309 9088 1343
rect 9036 1300 9088 1309
rect 6954 1062 7006 1114
rect 7018 1062 7070 1114
rect 7082 1062 7134 1114
<< metal2 >>
rect 5078 14498 5134 15000
rect 3608 14476 3660 14482
rect 3608 14418 3660 14424
rect 4816 14470 5134 14498
rect 3240 14408 3292 14414
rect 3240 14350 3292 14356
rect 1124 14272 1176 14278
rect 1124 14214 1176 14220
rect 1136 13394 1164 14214
rect 2320 13728 2372 13734
rect 2320 13670 2372 13676
rect 1124 13388 1176 13394
rect 1124 13330 1176 13336
rect 2228 13252 2280 13258
rect 2228 13194 2280 13200
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 1768 13184 1820 13190
rect 1768 13126 1820 13132
rect 940 12844 992 12850
rect 940 12786 992 12792
rect 952 11898 980 12786
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1412 12617 1440 12718
rect 1398 12608 1454 12617
rect 1398 12543 1454 12552
rect 1504 12374 1532 12718
rect 1492 12368 1544 12374
rect 1492 12310 1544 12316
rect 1216 12232 1268 12238
rect 1216 12174 1268 12180
rect 940 11892 992 11898
rect 940 11834 992 11840
rect 386 11792 442 11801
rect 386 11727 442 11736
rect 400 10742 428 11727
rect 1032 11076 1084 11082
rect 1032 11018 1084 11024
rect 1044 10985 1072 11018
rect 1030 10976 1086 10985
rect 1030 10911 1086 10920
rect 388 10736 440 10742
rect 388 10678 440 10684
rect 1228 10470 1256 12174
rect 1400 12164 1452 12170
rect 1400 12106 1452 12112
rect 1412 11830 1440 12106
rect 1400 11824 1452 11830
rect 1400 11766 1452 11772
rect 1216 10464 1268 10470
rect 1216 10406 1268 10412
rect 478 10160 534 10169
rect 478 10095 480 10104
rect 532 10095 534 10104
rect 480 10066 532 10072
rect 386 9344 442 9353
rect 386 9279 442 9288
rect 400 9042 428 9279
rect 388 9036 440 9042
rect 388 8978 440 8984
rect 1228 8498 1256 10406
rect 1412 10266 1440 11766
rect 1400 10260 1452 10266
rect 1400 10202 1452 10208
rect 1216 8492 1268 8498
rect 1216 8434 1268 8440
rect 1596 8294 1624 13126
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1688 9654 1716 10202
rect 1676 9648 1728 9654
rect 1676 9590 1728 9596
rect 1676 9512 1728 9518
rect 1676 9454 1728 9460
rect 1688 8498 1716 9454
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1584 8288 1636 8294
rect 1584 8230 1636 8236
rect 1400 8084 1452 8090
rect 1400 8026 1452 8032
rect 1124 7880 1176 7886
rect 1124 7822 1176 7828
rect 938 7712 994 7721
rect 938 7647 994 7656
rect 952 7410 980 7647
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 1136 6458 1164 7822
rect 1412 7818 1440 8026
rect 1400 7812 1452 7818
rect 1400 7754 1452 7760
rect 1308 7744 1360 7750
rect 1360 7692 1440 7698
rect 1308 7686 1440 7692
rect 1320 7670 1440 7686
rect 1412 7546 1440 7670
rect 1688 7546 1716 8434
rect 1780 8022 1808 13126
rect 2136 12300 2188 12306
rect 2136 12242 2188 12248
rect 2148 11830 2176 12242
rect 2136 11824 2188 11830
rect 1964 11784 2136 11812
rect 1964 11082 1992 11784
rect 2136 11766 2188 11772
rect 2134 11248 2190 11257
rect 2134 11183 2190 11192
rect 2148 11150 2176 11183
rect 2240 11150 2268 13194
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 1952 11076 2004 11082
rect 1952 11018 2004 11024
rect 1964 10606 1992 11018
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 1860 9988 1912 9994
rect 1860 9930 1912 9936
rect 1768 8016 1820 8022
rect 1768 7958 1820 7964
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 1676 7540 1728 7546
rect 1676 7482 1728 7488
rect 1216 7404 1268 7410
rect 1216 7346 1268 7352
rect 1228 6905 1256 7346
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1124 6452 1176 6458
rect 1124 6394 1176 6400
rect 480 6316 532 6322
rect 480 6258 532 6264
rect 492 6089 520 6258
rect 478 6080 534 6089
rect 478 6015 534 6024
rect 388 5772 440 5778
rect 388 5714 440 5720
rect 400 5273 428 5714
rect 1124 5704 1176 5710
rect 1124 5646 1176 5652
rect 386 5264 442 5273
rect 386 5199 442 5208
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 478 4448 534 4457
rect 478 4383 534 4392
rect 492 4146 520 4383
rect 952 4282 980 5102
rect 1136 4826 1164 5646
rect 1216 5160 1268 5166
rect 1216 5102 1268 5108
rect 1124 4820 1176 4826
rect 1124 4762 1176 4768
rect 940 4276 992 4282
rect 940 4218 992 4224
rect 480 4140 532 4146
rect 480 4082 532 4088
rect 952 2825 980 4218
rect 1228 4010 1256 5102
rect 1872 4622 1900 9930
rect 1964 9722 1992 10542
rect 2240 10266 2268 10542
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2044 10124 2096 10130
rect 2044 10066 2096 10072
rect 1952 9716 2004 9722
rect 1952 9658 2004 9664
rect 1952 9512 2004 9518
rect 2056 9500 2084 10066
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2004 9472 2084 9500
rect 1952 9454 2004 9460
rect 1952 7744 2004 7750
rect 1952 7686 2004 7692
rect 1964 7478 1992 7686
rect 1952 7472 2004 7478
rect 1952 7414 2004 7420
rect 2148 7410 2176 9998
rect 2332 9926 2360 13670
rect 2544 13626 2744 14192
rect 2944 14170 3144 14192
rect 2944 14118 2954 14170
rect 3006 14118 3018 14170
rect 3070 14118 3082 14170
rect 3134 14118 3144 14170
rect 2780 13728 2832 13734
rect 2832 13688 2912 13716
rect 2780 13670 2832 13676
rect 2544 13574 2554 13626
rect 2606 13574 2618 13626
rect 2670 13574 2682 13626
rect 2734 13574 2744 13626
rect 2544 13156 2744 13574
rect 2544 13100 2576 13156
rect 2632 13100 2656 13156
rect 2712 13100 2744 13156
rect 2544 13076 2744 13100
rect 2544 13020 2576 13076
rect 2632 13020 2656 13076
rect 2712 13020 2744 13076
rect 2544 12538 2744 13020
rect 2780 12640 2832 12646
rect 2780 12582 2832 12588
rect 2544 12486 2554 12538
rect 2606 12486 2618 12538
rect 2670 12486 2682 12538
rect 2734 12486 2744 12538
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2424 11694 2452 11834
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2544 11450 2744 12486
rect 2792 11626 2820 12582
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2778 11520 2834 11529
rect 2778 11455 2834 11464
rect 2544 11398 2554 11450
rect 2606 11398 2618 11450
rect 2670 11398 2682 11450
rect 2734 11398 2744 11450
rect 2410 10568 2466 10577
rect 2410 10503 2466 10512
rect 2320 9920 2372 9926
rect 2320 9862 2372 9868
rect 2424 9450 2452 10503
rect 2544 10362 2744 11398
rect 2792 11354 2820 11455
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2780 11008 2832 11014
rect 2780 10950 2832 10956
rect 2792 10470 2820 10950
rect 2780 10464 2832 10470
rect 2780 10406 2832 10412
rect 2544 10310 2554 10362
rect 2606 10310 2618 10362
rect 2670 10310 2682 10362
rect 2734 10310 2744 10362
rect 2412 9444 2464 9450
rect 2412 9386 2464 9392
rect 2544 9274 2744 10310
rect 2792 10266 2820 10406
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2780 9716 2832 9722
rect 2884 9704 2912 13688
rect 2832 9676 2912 9704
rect 2944 13556 3144 14118
rect 3252 13870 3280 14350
rect 3344 13956 3544 14192
rect 3344 13900 3376 13956
rect 3432 13900 3456 13956
rect 3512 13900 3544 13956
rect 3344 13876 3544 13900
rect 3240 13864 3292 13870
rect 3240 13806 3292 13812
rect 3344 13820 3376 13876
rect 3432 13820 3456 13876
rect 3512 13820 3544 13876
rect 2944 13500 2976 13556
rect 3032 13500 3056 13556
rect 3112 13500 3144 13556
rect 2944 13476 3144 13500
rect 2944 13420 2976 13476
rect 3032 13420 3056 13476
rect 3112 13420 3144 13476
rect 2944 13082 3144 13420
rect 2944 13030 2954 13082
rect 3006 13030 3018 13082
rect 3070 13030 3082 13082
rect 3134 13030 3144 13082
rect 2944 11994 3144 13030
rect 3240 12776 3292 12782
rect 3240 12718 3292 12724
rect 3252 12442 3280 12718
rect 3240 12436 3292 12442
rect 3240 12378 3292 12384
rect 3238 12064 3294 12073
rect 3238 11999 3294 12008
rect 2944 11942 2954 11994
rect 3006 11942 3018 11994
rect 3070 11942 3082 11994
rect 3134 11942 3144 11994
rect 2944 10906 3144 11942
rect 3252 11286 3280 11999
rect 3240 11280 3292 11286
rect 3240 11222 3292 11228
rect 2944 10854 2954 10906
rect 3006 10854 3018 10906
rect 3070 10854 3082 10906
rect 3134 10854 3144 10906
rect 2944 9818 3144 10854
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3252 10198 3280 10542
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3344 9956 3544 13820
rect 3620 13394 3648 14418
rect 4620 14340 4672 14346
rect 4620 14282 4672 14288
rect 3608 13388 3660 13394
rect 3608 13330 3660 13336
rect 3608 13252 3660 13258
rect 3608 13194 3660 13200
rect 3620 12238 3648 13194
rect 3608 12232 3660 12238
rect 3606 12200 3608 12209
rect 3660 12200 3662 12209
rect 3606 12135 3662 12144
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11830 3648 12038
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3620 10742 3648 11766
rect 3608 10736 3660 10742
rect 3608 10678 3660 10684
rect 3620 10130 3648 10678
rect 3744 10356 3944 14192
rect 4160 14000 4212 14006
rect 4212 13948 4384 13954
rect 4160 13942 4384 13948
rect 3976 13932 4028 13938
rect 4172 13926 4384 13942
rect 3976 13874 4028 13880
rect 3988 13530 4016 13874
rect 4068 13728 4120 13734
rect 4068 13670 4120 13676
rect 3976 13524 4028 13530
rect 3976 13466 4028 13472
rect 4080 12186 4108 13670
rect 4252 13184 4304 13190
rect 4252 13126 4304 13132
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4172 12374 4200 12854
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 3744 10300 3776 10356
rect 3832 10300 3856 10356
rect 3912 10300 3944 10356
rect 3744 10276 3944 10300
rect 3744 10220 3776 10276
rect 3832 10220 3856 10276
rect 3912 10220 3944 10276
rect 3608 10124 3660 10130
rect 3608 10066 3660 10072
rect 3240 9920 3292 9926
rect 3240 9862 3292 9868
rect 3344 9900 3376 9956
rect 3432 9900 3456 9956
rect 3512 9900 3544 9956
rect 3344 9876 3544 9900
rect 2944 9766 2954 9818
rect 3006 9766 3018 9818
rect 3070 9766 3082 9818
rect 3134 9766 3144 9818
rect 2780 9658 2832 9664
rect 2944 9556 3144 9766
rect 2944 9500 2976 9556
rect 3032 9500 3056 9556
rect 3112 9500 3144 9556
rect 3252 9518 3280 9862
rect 3344 9820 3376 9876
rect 3432 9820 3456 9876
rect 3512 9820 3544 9876
rect 2944 9476 3144 9500
rect 2944 9420 2976 9476
rect 3032 9420 3056 9476
rect 3112 9420 3144 9476
rect 3240 9512 3292 9518
rect 3240 9454 3292 9460
rect 2780 9376 2832 9382
rect 2780 9318 2832 9324
rect 2544 9222 2554 9274
rect 2606 9222 2618 9274
rect 2670 9222 2682 9274
rect 2734 9222 2744 9274
rect 2544 9156 2744 9222
rect 2544 9100 2576 9156
rect 2632 9100 2656 9156
rect 2712 9100 2744 9156
rect 2544 9076 2744 9100
rect 2544 9020 2576 9076
rect 2632 9020 2656 9076
rect 2712 9020 2744 9076
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2136 7404 2188 7410
rect 2136 7346 2188 7352
rect 1308 4616 1360 4622
rect 1308 4558 1360 4564
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1216 4004 1268 4010
rect 1216 3946 1268 3952
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 386 2544 442 2553
rect 1320 2514 1348 4558
rect 1872 2774 1900 4558
rect 1872 2746 1992 2774
rect 1964 2553 1992 2746
rect 2240 2650 2268 8910
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2424 8566 2452 8774
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2544 8186 2744 9020
rect 2792 8922 2820 9318
rect 2792 8894 2912 8922
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2544 8134 2554 8186
rect 2606 8134 2618 8186
rect 2670 8134 2682 8186
rect 2734 8134 2744 8186
rect 2320 8016 2372 8022
rect 2320 7958 2372 7964
rect 2332 7886 2360 7958
rect 2320 7880 2372 7886
rect 2320 7822 2372 7828
rect 2320 7404 2372 7410
rect 2320 7346 2372 7352
rect 2332 5234 2360 7346
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2332 4758 2360 5170
rect 2424 5166 2452 7278
rect 2544 7098 2744 8134
rect 2792 8090 2820 8774
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2780 7948 2832 7954
rect 2780 7890 2832 7896
rect 2544 7046 2554 7098
rect 2606 7046 2618 7098
rect 2670 7046 2682 7098
rect 2734 7046 2744 7098
rect 2544 6010 2744 7046
rect 2544 5958 2554 6010
rect 2606 5958 2618 6010
rect 2670 5958 2682 6010
rect 2734 5958 2744 6010
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2544 5156 2744 5958
rect 2544 5100 2576 5156
rect 2632 5100 2656 5156
rect 2712 5100 2744 5156
rect 2544 5076 2744 5100
rect 2544 5020 2576 5076
rect 2632 5020 2656 5076
rect 2712 5020 2744 5076
rect 2544 4922 2744 5020
rect 2544 4870 2554 4922
rect 2606 4870 2618 4922
rect 2670 4870 2682 4922
rect 2734 4870 2744 4922
rect 2320 4752 2372 4758
rect 2320 4694 2372 4700
rect 2544 4094 2744 4870
rect 2792 4690 2820 7890
rect 2780 4684 2832 4690
rect 2780 4626 2832 4632
rect 2228 2644 2280 2650
rect 2228 2586 2280 2592
rect 1950 2544 2006 2553
rect 386 2479 442 2488
rect 1308 2508 1360 2514
rect 400 2009 428 2479
rect 1950 2479 2006 2488
rect 1308 2450 1360 2456
rect 900 2356 1100 2365
rect 900 2300 932 2356
rect 988 2300 1012 2356
rect 1068 2300 1100 2356
rect 900 2276 1100 2300
rect 900 2220 932 2276
rect 988 2220 1012 2276
rect 1068 2220 1100 2276
rect 900 2211 1100 2220
rect 386 2000 442 2009
rect 386 1935 442 1944
rect 1500 1956 1700 1965
rect 1500 1900 1532 1956
rect 1588 1900 1612 1956
rect 1668 1900 1700 1956
rect 1500 1876 1700 1900
rect 1500 1820 1532 1876
rect 1588 1820 1612 1876
rect 1668 1820 1700 1876
rect 1500 1811 1700 1820
rect 2884 1766 2912 8894
rect 2944 8730 3144 9420
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 2944 8678 2954 8730
rect 3006 8678 3018 8730
rect 3070 8678 3082 8730
rect 3134 8678 3144 8730
rect 2944 7642 3144 8678
rect 3252 8566 3280 9318
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 2944 7590 2954 7642
rect 3006 7590 3018 7642
rect 3070 7590 3082 7642
rect 3134 7590 3144 7642
rect 2944 6554 3144 7590
rect 3252 7546 3280 7822
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 2944 6502 2954 6554
rect 3006 6502 3018 6554
rect 3070 6502 3082 6554
rect 3134 6502 3144 6554
rect 2944 5556 3144 6502
rect 2944 5500 2976 5556
rect 3032 5500 3056 5556
rect 3112 5500 3144 5556
rect 2944 5476 3144 5500
rect 2944 5466 2976 5476
rect 3032 5466 3056 5476
rect 3112 5466 3144 5476
rect 2944 5414 2954 5466
rect 3006 5414 3018 5420
rect 3070 5414 3082 5420
rect 3134 5414 3144 5466
rect 2944 4378 3144 5414
rect 2944 4326 2954 4378
rect 3006 4326 3018 4378
rect 3070 4326 3082 4378
rect 3134 4326 3144 4378
rect 2944 4094 3144 4326
rect 3344 5956 3544 9820
rect 3620 8838 3648 10066
rect 3608 8832 3660 8838
rect 3608 8774 3660 8780
rect 3620 8634 3648 8774
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 3608 8424 3660 8430
rect 3608 8366 3660 8372
rect 3620 7954 3648 8366
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3344 5900 3376 5956
rect 3432 5900 3456 5956
rect 3512 5900 3544 5956
rect 3344 5876 3544 5900
rect 3344 5820 3376 5876
rect 3432 5820 3456 5876
rect 3512 5820 3544 5876
rect 3344 4094 3544 5820
rect 3744 6356 3944 10220
rect 3988 12158 4108 12186
rect 4160 12232 4212 12238
rect 4160 12174 4212 12180
rect 3988 9654 4016 12158
rect 4068 12096 4120 12102
rect 4068 12038 4120 12044
rect 3976 9648 4028 9654
rect 3976 9590 4028 9596
rect 4080 8974 4108 12038
rect 4172 11218 4200 12174
rect 4264 11257 4292 13126
rect 4250 11248 4306 11257
rect 4160 11212 4212 11218
rect 4250 11183 4306 11192
rect 4160 11154 4212 11160
rect 4172 10810 4200 11154
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 4252 10464 4304 10470
rect 4252 10406 4304 10412
rect 4264 9654 4292 10406
rect 4252 9648 4304 9654
rect 4252 9590 4304 9596
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4252 8968 4304 8974
rect 4356 8956 4384 13926
rect 4528 13456 4580 13462
rect 4448 13416 4528 13444
rect 4448 13326 4476 13416
rect 4528 13398 4580 13404
rect 4632 13394 4660 14282
rect 4816 14074 4844 14470
rect 5078 14400 5134 14470
rect 5354 14400 5410 15000
rect 5630 14498 5686 15000
rect 5906 14498 5962 15000
rect 6182 14498 6238 15000
rect 6458 14498 6514 15000
rect 6734 14498 6790 15000
rect 7010 14498 7066 15000
rect 7286 14498 7342 15000
rect 7562 14498 7618 15000
rect 7838 14498 7894 15000
rect 8114 14498 8170 15000
rect 8390 14498 8446 15000
rect 5552 14470 5686 14498
rect 5736 14482 5962 14498
rect 4804 14068 4856 14074
rect 4804 14010 4856 14016
rect 4712 13932 4764 13938
rect 4712 13874 4764 13880
rect 4620 13388 4672 13394
rect 4620 13330 4672 13336
rect 4436 13320 4488 13326
rect 4436 13262 4488 13268
rect 4724 12434 4752 13874
rect 5172 13796 5224 13802
rect 5172 13738 5224 13744
rect 4988 13728 5040 13734
rect 4988 13670 5040 13676
rect 4632 12406 4752 12434
rect 4528 11552 4580 11558
rect 4528 11494 4580 11500
rect 4540 9178 4568 11494
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4436 9104 4488 9110
rect 4436 9046 4488 9052
rect 4304 8928 4384 8956
rect 4252 8910 4304 8916
rect 4160 8900 4212 8906
rect 4160 8842 4212 8848
rect 4172 8537 4200 8842
rect 4344 8832 4396 8838
rect 4344 8774 4396 8780
rect 4356 8634 4384 8774
rect 4344 8628 4396 8634
rect 4344 8570 4396 8576
rect 4448 8566 4476 9046
rect 4436 8560 4488 8566
rect 4158 8528 4214 8537
rect 4436 8502 4488 8508
rect 4158 8463 4214 8472
rect 4632 7750 4660 12406
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4724 11354 4752 12174
rect 4804 11552 4856 11558
rect 4804 11494 4856 11500
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4712 7880 4764 7886
rect 4712 7822 4764 7828
rect 4620 7744 4672 7750
rect 4620 7686 4672 7692
rect 4724 7342 4752 7822
rect 4816 7478 4844 11494
rect 4896 11076 4948 11082
rect 4896 11018 4948 11024
rect 4908 10810 4936 11018
rect 4896 10804 4948 10810
rect 4896 10746 4948 10752
rect 5000 10577 5028 13670
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 5092 12850 5120 13194
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5184 12434 5212 13738
rect 5356 13456 5408 13462
rect 5356 13398 5408 13404
rect 5184 12406 5304 12434
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5092 11558 5120 12174
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 4986 10568 5042 10577
rect 4986 10503 5042 10512
rect 5172 10464 5224 10470
rect 5172 10406 5224 10412
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 4896 9716 4948 9722
rect 4896 9658 4948 9664
rect 4908 7834 4936 9658
rect 4988 9512 5040 9518
rect 5092 9466 5120 9998
rect 5040 9460 5120 9466
rect 4988 9454 5120 9460
rect 5000 9438 5120 9454
rect 5092 9042 5120 9438
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 4908 7806 5028 7834
rect 4896 7744 4948 7750
rect 4896 7686 4948 7692
rect 4804 7472 4856 7478
rect 4804 7414 4856 7420
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 3976 7200 4028 7206
rect 3976 7142 4028 7148
rect 3988 6458 4016 7142
rect 4908 6866 4936 7686
rect 4896 6860 4948 6866
rect 4896 6802 4948 6808
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3744 6300 3776 6356
rect 3832 6300 3856 6356
rect 3912 6300 3944 6356
rect 3744 6276 3944 6300
rect 3744 6220 3776 6276
rect 3832 6220 3856 6276
rect 3912 6220 3944 6276
rect 3148 2440 3200 2446
rect 3148 2382 3200 2388
rect 2872 1760 2924 1766
rect 2872 1702 2924 1708
rect 3160 1562 3188 2382
rect 3744 2356 3944 6220
rect 3988 5778 4016 6394
rect 4264 6254 4292 6734
rect 4908 6458 4936 6802
rect 4896 6452 4948 6458
rect 4896 6394 4948 6400
rect 4252 6248 4304 6254
rect 4252 6190 4304 6196
rect 3976 5772 4028 5778
rect 3976 5714 4028 5720
rect 4160 4276 4212 4282
rect 4160 4218 4212 4224
rect 4172 3602 4200 4218
rect 4264 3641 4292 6190
rect 4804 5704 4856 5710
rect 4804 5646 4856 5652
rect 4816 4690 4844 5646
rect 5000 4826 5028 7806
rect 5092 7410 5120 8978
rect 5184 8974 5212 10406
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 5276 7562 5304 12406
rect 5368 11762 5396 13398
rect 5552 12102 5580 14470
rect 5630 14400 5686 14470
rect 5724 14476 5962 14482
rect 5776 14470 5962 14476
rect 5724 14418 5776 14424
rect 5906 14400 5962 14470
rect 6012 14470 6238 14498
rect 6012 13530 6040 14470
rect 6182 14400 6238 14470
rect 6288 14470 6514 14498
rect 6288 14278 6316 14470
rect 6458 14400 6514 14470
rect 6564 14470 6790 14498
rect 6564 14362 6592 14470
rect 6734 14400 6790 14470
rect 6840 14470 7066 14498
rect 6472 14334 6592 14362
rect 6276 14272 6328 14278
rect 6276 14214 6328 14220
rect 6368 14272 6420 14278
rect 6368 14214 6420 14220
rect 6380 13802 6408 14214
rect 6368 13796 6420 13802
rect 6368 13738 6420 13744
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6000 13524 6052 13530
rect 6000 13466 6052 13472
rect 5632 13252 5684 13258
rect 5632 13194 5684 13200
rect 5908 13252 5960 13258
rect 5908 13194 5960 13200
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5644 11937 5672 13194
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5630 11928 5686 11937
rect 5630 11863 5686 11872
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5356 11756 5408 11762
rect 5356 11698 5408 11704
rect 5460 11054 5488 11766
rect 5630 11656 5686 11665
rect 5630 11591 5686 11600
rect 5368 11026 5488 11054
rect 5368 7886 5396 11026
rect 5644 11014 5672 11591
rect 5736 11150 5764 11834
rect 5724 11144 5776 11150
rect 5724 11086 5776 11092
rect 5632 11008 5684 11014
rect 5632 10950 5684 10956
rect 5446 10840 5502 10849
rect 5446 10775 5502 10784
rect 5356 7880 5408 7886
rect 5356 7822 5408 7828
rect 5276 7534 5396 7562
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5080 5160 5132 5166
rect 5080 5102 5132 5108
rect 4988 4820 5040 4826
rect 4988 4762 5040 4768
rect 4804 4684 4856 4690
rect 4804 4626 4856 4632
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4724 4154 4752 4422
rect 4816 4282 4844 4626
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4724 4126 4844 4154
rect 4816 4078 4844 4126
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 5092 3738 5120 5102
rect 5276 4622 5304 6258
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 4154 5304 4558
rect 5184 4146 5304 4154
rect 5172 4140 5304 4146
rect 5224 4126 5304 4140
rect 5172 4082 5224 4088
rect 5184 4010 5212 4082
rect 5264 4072 5316 4078
rect 5264 4014 5316 4020
rect 5172 4004 5224 4010
rect 5172 3946 5224 3952
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4250 3632 4306 3641
rect 4160 3596 4212 3602
rect 4250 3567 4306 3576
rect 4710 3632 4766 3641
rect 4710 3567 4766 3576
rect 4804 3596 4856 3602
rect 4160 3538 4212 3544
rect 4724 2446 4752 3567
rect 4804 3538 4856 3544
rect 4712 2440 4764 2446
rect 4712 2382 4764 2388
rect 3744 2300 3776 2356
rect 3832 2300 3856 2356
rect 3912 2300 3944 2356
rect 3744 2276 3944 2300
rect 3744 2220 3776 2276
rect 3832 2220 3856 2276
rect 3912 2220 3944 2276
rect 3148 1556 3200 1562
rect 3148 1498 3200 1504
rect 3744 1040 3944 2220
rect 4816 1970 4844 3538
rect 5184 3466 5212 3946
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5276 2038 5304 4014
rect 5368 3505 5396 7534
rect 5460 5302 5488 10775
rect 5632 10668 5684 10674
rect 5632 10610 5684 10616
rect 5540 10124 5592 10130
rect 5540 10066 5592 10072
rect 5552 9994 5580 10066
rect 5644 9994 5672 10610
rect 5540 9988 5592 9994
rect 5540 9930 5592 9936
rect 5632 9988 5684 9994
rect 5632 9930 5684 9936
rect 5736 9722 5764 11086
rect 5828 10849 5856 12582
rect 5920 11665 5948 13194
rect 6000 12776 6052 12782
rect 6000 12718 6052 12724
rect 5906 11656 5962 11665
rect 5906 11591 5962 11600
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11218 5948 11494
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5814 10840 5870 10849
rect 5814 10775 5870 10784
rect 5816 10668 5868 10674
rect 5816 10610 5868 10616
rect 5828 10198 5856 10610
rect 6012 10266 6040 12718
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6104 12170 6132 12582
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6196 11762 6224 13670
rect 6472 13138 6500 14334
rect 6840 14278 6868 14470
rect 7010 14400 7066 14470
rect 7116 14470 7342 14498
rect 7116 14346 7144 14470
rect 7286 14400 7342 14470
rect 7392 14470 7618 14498
rect 7392 14362 7420 14470
rect 7562 14400 7618 14470
rect 7668 14470 7894 14498
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7208 14334 7420 14362
rect 6828 14272 6880 14278
rect 6828 14214 6880 14220
rect 6380 13110 6500 13138
rect 6544 13626 6744 14192
rect 6544 13574 6554 13626
rect 6606 13574 6618 13626
rect 6670 13574 6682 13626
rect 6734 13574 6744 13626
rect 6544 13156 6744 13574
rect 6944 14170 7144 14192
rect 6944 14118 6954 14170
rect 7006 14118 7018 14170
rect 7070 14118 7082 14170
rect 7134 14118 7144 14170
rect 6944 13556 7144 14118
rect 6944 13500 6976 13556
rect 7032 13500 7056 13556
rect 7112 13500 7144 13556
rect 6944 13476 7144 13500
rect 6944 13420 6976 13476
rect 7032 13420 7056 13476
rect 7112 13420 7144 13476
rect 7208 13462 7236 14334
rect 7344 13956 7544 14192
rect 7668 14074 7696 14470
rect 7838 14400 7894 14470
rect 8036 14470 8170 14498
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7344 13900 7376 13956
rect 7432 13900 7456 13956
rect 7512 13900 7544 13956
rect 7344 13876 7544 13900
rect 7344 13820 7376 13876
rect 7432 13820 7456 13876
rect 7512 13820 7544 13876
rect 7656 13932 7708 13938
rect 7656 13874 7708 13880
rect 6828 13320 6880 13326
rect 6828 13262 6880 13268
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 6288 11898 6316 12786
rect 6380 12442 6408 13110
rect 6544 13100 6576 13156
rect 6632 13100 6656 13156
rect 6712 13100 6744 13156
rect 6544 13076 6744 13100
rect 6544 13020 6576 13076
rect 6632 13020 6656 13076
rect 6712 13020 6744 13076
rect 6460 12980 6512 12986
rect 6460 12922 6512 12928
rect 6368 12436 6420 12442
rect 6368 12378 6420 12384
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5816 10192 5868 10198
rect 5816 10134 5868 10140
rect 5724 9716 5776 9722
rect 5724 9658 5776 9664
rect 5828 9654 5856 10134
rect 5908 10056 5960 10062
rect 5908 9998 5960 10004
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5828 8906 5856 9590
rect 5920 9178 5948 9998
rect 6000 9988 6052 9994
rect 6000 9930 6052 9936
rect 6012 9586 6040 9930
rect 6000 9580 6052 9586
rect 6000 9522 6052 9528
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 5816 8900 5868 8906
rect 5816 8842 5868 8848
rect 6012 8786 6040 9522
rect 5920 8758 6040 8786
rect 5724 8560 5776 8566
rect 5724 8502 5776 8508
rect 5632 8288 5684 8294
rect 5632 8230 5684 8236
rect 5644 7886 5672 8230
rect 5540 7880 5592 7886
rect 5540 7822 5592 7828
rect 5632 7880 5684 7886
rect 5632 7822 5684 7828
rect 5552 7290 5580 7822
rect 5644 7410 5672 7822
rect 5736 7750 5764 8502
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5724 7744 5776 7750
rect 5724 7686 5776 7692
rect 5736 7410 5764 7686
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5552 7262 5672 7290
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6730 5580 7142
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5644 6322 5672 7262
rect 5632 6316 5684 6322
rect 5632 6258 5684 6264
rect 5736 6118 5764 7346
rect 5828 6934 5856 8434
rect 5920 7410 5948 8758
rect 6104 7970 6132 11630
rect 6196 10810 6224 11698
rect 6366 11656 6422 11665
rect 6276 11620 6328 11626
rect 6366 11591 6422 11600
rect 6276 11562 6328 11568
rect 6184 10804 6236 10810
rect 6184 10746 6236 10752
rect 6288 10674 6316 11562
rect 6276 10668 6328 10674
rect 6276 10610 6328 10616
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 6196 8906 6224 10474
rect 6288 9926 6316 10610
rect 6276 9920 6328 9926
rect 6276 9862 6328 9868
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6012 7942 6132 7970
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5448 5296 5500 5302
rect 5448 5238 5500 5244
rect 5540 4276 5592 4282
rect 5540 4218 5592 4224
rect 5354 3496 5410 3505
rect 5354 3431 5410 3440
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 5460 2650 5488 3402
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5552 2446 5580 4218
rect 5828 4154 5856 6258
rect 5920 6254 5948 7346
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 6012 5370 6040 7942
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6104 6458 6132 7822
rect 6196 7002 6224 8842
rect 6380 8022 6408 11591
rect 6472 10810 6500 12922
rect 6544 12538 6744 13020
rect 6840 12889 6868 13262
rect 6944 13082 7144 13420
rect 7196 13456 7248 13462
rect 7196 13398 7248 13404
rect 6944 13030 6954 13082
rect 7006 13030 7018 13082
rect 7070 13030 7082 13082
rect 7134 13030 7144 13082
rect 6826 12880 6882 12889
rect 6826 12815 6882 12824
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6544 12486 6554 12538
rect 6606 12486 6618 12538
rect 6670 12486 6682 12538
rect 6734 12486 6744 12538
rect 6544 11450 6744 12486
rect 6544 11398 6554 11450
rect 6606 11398 6618 11450
rect 6670 11398 6682 11450
rect 6734 11398 6744 11450
rect 6460 10804 6512 10810
rect 6460 10746 6512 10752
rect 6460 10600 6512 10606
rect 6460 10542 6512 10548
rect 6472 10266 6500 10542
rect 6544 10362 6744 11398
rect 6840 11354 6868 12718
rect 6944 11994 7144 13030
rect 7194 12880 7250 12889
rect 7194 12815 7250 12824
rect 7208 12374 7236 12815
rect 7196 12368 7248 12374
rect 7196 12310 7248 12316
rect 6944 11942 6954 11994
rect 7006 11942 7018 11994
rect 7070 11942 7082 11994
rect 7134 11942 7144 11994
rect 6828 11348 6880 11354
rect 6828 11290 6880 11296
rect 6828 11008 6880 11014
rect 6828 10950 6880 10956
rect 6840 10810 6868 10950
rect 6944 10906 7144 11942
rect 6944 10854 6954 10906
rect 7006 10854 7018 10906
rect 7070 10854 7082 10906
rect 7134 10854 7144 10906
rect 6828 10804 6880 10810
rect 6828 10746 6880 10752
rect 6544 10310 6554 10362
rect 6606 10310 6618 10362
rect 6670 10310 6682 10362
rect 6734 10310 6744 10362
rect 6460 10260 6512 10266
rect 6460 10202 6512 10208
rect 6460 10124 6512 10130
rect 6460 10066 6512 10072
rect 6472 9518 6500 10066
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6544 9274 6744 10310
rect 6544 9222 6554 9274
rect 6606 9222 6618 9274
rect 6670 9222 6682 9274
rect 6734 9222 6744 9274
rect 6544 9156 6744 9222
rect 6544 9100 6576 9156
rect 6632 9100 6656 9156
rect 6712 9100 6744 9156
rect 6544 9076 6744 9100
rect 6544 9020 6576 9076
rect 6632 9020 6656 9076
rect 6712 9020 6744 9076
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6368 8016 6420 8022
rect 6368 7958 6420 7964
rect 6276 7880 6328 7886
rect 6276 7822 6328 7828
rect 6288 7342 6316 7822
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6092 6452 6144 6458
rect 6092 6394 6144 6400
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5710 6224 6054
rect 6288 5778 6316 7278
rect 6380 6798 6408 7686
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6472 6322 6500 8298
rect 6544 8186 6744 9020
rect 6944 9818 7144 10854
rect 6944 9766 6954 9818
rect 7006 9766 7018 9818
rect 7070 9766 7082 9818
rect 7134 9766 7144 9818
rect 6944 9556 7144 9766
rect 6944 9500 6976 9556
rect 7032 9500 7056 9556
rect 7112 9500 7144 9556
rect 6944 9476 7144 9500
rect 6944 9420 6976 9476
rect 7032 9420 7056 9476
rect 7112 9420 7144 9476
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6840 8566 6868 8910
rect 6944 8730 7144 9420
rect 7344 9956 7544 13820
rect 7668 12442 7696 13874
rect 7656 12436 7708 12442
rect 7656 12378 7708 12384
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7668 12102 7696 12174
rect 7656 12096 7708 12102
rect 7656 12038 7708 12044
rect 7344 9900 7376 9956
rect 7432 9900 7456 9956
rect 7512 9900 7544 9956
rect 7344 9876 7544 9900
rect 7344 9820 7376 9876
rect 7432 9820 7456 9876
rect 7512 9820 7544 9876
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 6944 8678 6954 8730
rect 7006 8678 7018 8730
rect 7070 8678 7082 8730
rect 7134 8678 7144 8730
rect 6828 8560 6880 8566
rect 6828 8502 6880 8508
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6544 8134 6554 8186
rect 6606 8134 6618 8186
rect 6670 8134 6682 8186
rect 6734 8134 6744 8186
rect 6544 7098 6744 8134
rect 6544 7046 6554 7098
rect 6606 7046 6618 7098
rect 6670 7046 6682 7098
rect 6734 7046 6744 7098
rect 6460 6316 6512 6322
rect 6460 6258 6512 6264
rect 6544 6010 6744 7046
rect 6544 5958 6554 6010
rect 6606 5958 6618 6010
rect 6670 5958 6682 6010
rect 6734 5958 6744 6010
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 6012 4570 6040 5306
rect 6380 5234 6408 5782
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6544 5156 6744 5958
rect 6840 5914 6868 8366
rect 6944 7642 7144 8678
rect 7208 8634 7236 8910
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7196 8288 7248 8294
rect 7194 8256 7196 8265
rect 7248 8256 7250 8265
rect 7194 8191 7250 8200
rect 6944 7590 6954 7642
rect 7006 7590 7018 7642
rect 7070 7590 7082 7642
rect 7134 7590 7144 7642
rect 6944 6554 7144 7590
rect 6944 6502 6954 6554
rect 7006 6502 7018 6554
rect 7070 6502 7082 6554
rect 7134 6502 7144 6554
rect 6828 5908 6880 5914
rect 6828 5850 6880 5856
rect 6544 5100 6576 5156
rect 6632 5100 6656 5156
rect 6712 5100 6744 5156
rect 6544 5076 6744 5100
rect 6544 5020 6576 5076
rect 6632 5020 6656 5076
rect 6712 5020 6744 5076
rect 6544 4922 6744 5020
rect 6544 4870 6554 4922
rect 6606 4870 6618 4922
rect 6670 4870 6682 4922
rect 6734 4870 6744 4922
rect 6012 4554 6132 4570
rect 6012 4548 6144 4554
rect 6012 4542 6092 4548
rect 6092 4490 6144 4496
rect 6092 4276 6144 4282
rect 6092 4218 6144 4224
rect 5828 4146 6040 4154
rect 5828 4140 6052 4146
rect 5828 4126 6000 4140
rect 6000 4082 6052 4088
rect 6104 4010 6132 4218
rect 6092 4004 6144 4010
rect 6092 3946 6144 3952
rect 6104 3466 6132 3946
rect 6544 3834 6744 4870
rect 6944 5556 7144 6502
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 6944 5500 6976 5556
rect 7032 5500 7056 5556
rect 7112 5500 7144 5556
rect 6944 5476 7144 5500
rect 6944 5466 6976 5476
rect 7032 5466 7056 5476
rect 7112 5466 7144 5476
rect 6944 5414 6954 5466
rect 7006 5414 7018 5420
rect 7070 5414 7082 5420
rect 7134 5414 7144 5466
rect 6944 4378 7144 5414
rect 6944 4326 6954 4378
rect 7006 4326 7018 4378
rect 7070 4326 7082 4378
rect 7134 4326 7144 4378
rect 6828 4072 6880 4078
rect 6828 4014 6880 4020
rect 6544 3782 6554 3834
rect 6606 3782 6618 3834
rect 6670 3782 6682 3834
rect 6734 3782 6744 3834
rect 6458 3496 6514 3505
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 6276 3460 6328 3466
rect 6458 3431 6514 3440
rect 6276 3402 6328 3408
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5644 2553 5672 2926
rect 5630 2544 5686 2553
rect 5630 2479 5686 2488
rect 5540 2440 5592 2446
rect 5540 2382 5592 2388
rect 5264 2032 5316 2038
rect 5264 1974 5316 1980
rect 6288 1970 6316 3402
rect 6472 2854 6500 3431
rect 6460 2848 6512 2854
rect 6460 2790 6512 2796
rect 6472 2038 6500 2790
rect 6544 2746 6744 3782
rect 6840 3738 6868 4014
rect 6828 3732 6880 3738
rect 6828 3674 6880 3680
rect 6944 3290 7144 4326
rect 7208 3942 7236 6190
rect 7344 5956 7544 9820
rect 7744 10356 7944 14192
rect 8036 13802 8064 14470
rect 8114 14400 8170 14470
rect 8220 14470 8446 14498
rect 8220 14414 8248 14470
rect 8208 14408 8260 14414
rect 8390 14400 8446 14470
rect 8666 14498 8722 15000
rect 8666 14470 8892 14498
rect 8666 14400 8722 14470
rect 8208 14350 8260 14356
rect 8864 14090 8892 14470
rect 8942 14400 8998 15000
rect 9218 14498 9274 15000
rect 9048 14470 9274 14498
rect 8864 14062 8984 14090
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8852 13932 8904 13938
rect 8852 13874 8904 13880
rect 8484 13864 8536 13870
rect 8484 13806 8536 13812
rect 8024 13796 8076 13802
rect 8024 13738 8076 13744
rect 8116 13728 8168 13734
rect 8116 13670 8168 13676
rect 8128 12306 8156 13670
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8116 12300 8168 12306
rect 8116 12242 8168 12248
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7744 10300 7776 10356
rect 7832 10300 7856 10356
rect 7912 10300 7944 10356
rect 7744 10276 7944 10300
rect 7744 10220 7776 10276
rect 7832 10220 7856 10276
rect 7912 10220 7944 10276
rect 7656 9648 7708 9654
rect 7656 9590 7708 9596
rect 7668 9178 7696 9590
rect 7656 9172 7708 9178
rect 7656 9114 7708 9120
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7668 7478 7696 8774
rect 7656 7472 7708 7478
rect 7656 7414 7708 7420
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7344 5900 7376 5956
rect 7432 5900 7456 5956
rect 7512 5900 7544 5956
rect 7344 5876 7544 5900
rect 7344 5820 7376 5876
rect 7432 5820 7456 5876
rect 7512 5820 7544 5876
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 6944 3238 6954 3290
rect 7006 3238 7018 3290
rect 7070 3238 7082 3290
rect 7134 3238 7144 3290
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6544 2694 6554 2746
rect 6606 2694 6618 2746
rect 6670 2694 6682 2746
rect 6734 2694 6744 2746
rect 6460 2032 6512 2038
rect 6460 1974 6512 1980
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 6276 1964 6328 1970
rect 6276 1906 6328 1912
rect 6460 1760 6512 1766
rect 6460 1702 6512 1708
rect 6472 1494 6500 1702
rect 6544 1658 6744 2694
rect 6840 2650 6868 3062
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6840 1766 6868 2314
rect 6944 2202 7144 3238
rect 7208 3058 7236 3538
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6944 2150 6954 2202
rect 7006 2150 7018 2202
rect 7070 2150 7082 2202
rect 7134 2150 7144 2202
rect 6828 1760 6880 1766
rect 6828 1702 6880 1708
rect 6544 1606 6554 1658
rect 6606 1606 6618 1658
rect 6670 1606 6682 1658
rect 6734 1606 6744 1658
rect 6460 1488 6512 1494
rect 6460 1430 6512 1436
rect 6544 1156 6744 1606
rect 6544 1100 6576 1156
rect 6632 1100 6656 1156
rect 6712 1100 6744 1156
rect 6544 1076 6744 1100
rect 6544 1020 6576 1076
rect 6632 1020 6656 1076
rect 6712 1020 6744 1076
rect 6944 1556 7144 2150
rect 6944 1500 6976 1556
rect 7032 1500 7056 1556
rect 7112 1500 7144 1556
rect 6944 1476 7144 1500
rect 6944 1420 6976 1476
rect 7032 1420 7056 1476
rect 7112 1420 7144 1476
rect 6944 1114 7144 1420
rect 6944 1062 6954 1114
rect 7006 1062 7018 1114
rect 7070 1062 7082 1114
rect 7134 1062 7144 1114
rect 6944 1040 7144 1062
rect 7344 1956 7544 5820
rect 7668 3670 7696 6734
rect 7744 6356 7944 10220
rect 8036 10062 8064 12174
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8128 11898 8156 12038
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8220 11762 8248 13126
rect 8392 12844 8444 12850
rect 8312 12804 8392 12832
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8128 10713 8156 11018
rect 8208 10736 8260 10742
rect 8114 10704 8170 10713
rect 8208 10678 8260 10684
rect 8114 10639 8170 10648
rect 8220 10198 8248 10678
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8024 9920 8076 9926
rect 8024 9862 8076 9868
rect 8036 8906 8064 9862
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7410 8064 7686
rect 8128 7410 8156 7754
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8116 7404 8168 7410
rect 8116 7346 8168 7352
rect 8116 6724 8168 6730
rect 8116 6666 8168 6672
rect 7744 6300 7776 6356
rect 7832 6300 7856 6356
rect 7912 6300 7944 6356
rect 7744 6276 7944 6300
rect 7744 6220 7776 6276
rect 7832 6220 7856 6276
rect 7912 6220 7944 6276
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7656 2984 7708 2990
rect 7656 2926 7708 2932
rect 7668 2106 7696 2926
rect 7744 2356 7944 6220
rect 8024 3528 8076 3534
rect 8024 3470 8076 3476
rect 7744 2300 7776 2356
rect 7832 2300 7856 2356
rect 7912 2300 7944 2356
rect 8036 2310 8064 3470
rect 8128 2938 8156 6666
rect 8220 5710 8248 9318
rect 8312 9178 8340 12804
rect 8392 12786 8444 12792
rect 8496 12345 8524 13806
rect 8482 12336 8538 12345
rect 8482 12271 8538 12280
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11830 8524 12038
rect 8588 11898 8616 13874
rect 8760 13252 8812 13258
rect 8680 13212 8760 13240
rect 8680 12238 8708 13212
rect 8760 13194 8812 13200
rect 8864 12646 8892 13874
rect 8956 12730 8984 14062
rect 9048 13530 9076 14470
rect 9218 14400 9274 14470
rect 9588 14000 9640 14006
rect 9586 13968 9588 13977
rect 9640 13968 9642 13977
rect 9586 13903 9642 13912
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9128 13320 9180 13326
rect 9128 13262 9180 13268
rect 8956 12702 9076 12730
rect 8852 12640 8904 12646
rect 8852 12582 8904 12588
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8680 12073 8708 12174
rect 8760 12096 8812 12102
rect 8666 12064 8722 12073
rect 8760 12038 8812 12044
rect 8666 11999 8722 12008
rect 8772 11914 8800 12038
rect 8576 11892 8628 11898
rect 8576 11834 8628 11840
rect 8680 11886 8800 11914
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8680 11082 8708 11886
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8760 11076 8812 11082
rect 8760 11018 8812 11024
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8496 10674 8524 10950
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8392 10464 8444 10470
rect 8392 10406 8444 10412
rect 8404 10062 8432 10406
rect 8392 10056 8444 10062
rect 8392 9998 8444 10004
rect 8576 10056 8628 10062
rect 8576 9998 8628 10004
rect 8588 9450 8616 9998
rect 8680 9926 8708 11018
rect 8772 10062 8800 11018
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8668 9920 8720 9926
rect 8668 9862 8720 9868
rect 8576 9444 8628 9450
rect 8576 9386 8628 9392
rect 8300 9172 8352 9178
rect 8300 9114 8352 9120
rect 8680 8974 8708 9862
rect 8864 9738 8892 12582
rect 8772 9710 8892 9738
rect 8668 8968 8720 8974
rect 8668 8910 8720 8916
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8312 7546 8340 7822
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8404 7449 8432 7890
rect 8496 7886 8524 8570
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8680 7886 8708 8502
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8390 7440 8446 7449
rect 8390 7375 8446 7384
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8680 6746 8708 7822
rect 8772 7546 8800 9710
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8864 9178 8892 9522
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8956 8498 8984 12582
rect 9048 10538 9076 12702
rect 9140 11529 9168 13262
rect 9232 13190 9260 13806
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9220 13184 9272 13190
rect 9600 13161 9628 13330
rect 9220 13126 9272 13132
rect 9586 13152 9642 13161
rect 9232 12238 9260 13126
rect 9586 13087 9642 13096
rect 9220 12232 9272 12238
rect 9220 12174 9272 12180
rect 9126 11520 9182 11529
rect 9126 11455 9182 11464
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9600 9897 9628 10066
rect 9586 9888 9642 9897
rect 9586 9823 9642 9832
rect 9586 9072 9642 9081
rect 9586 9007 9642 9016
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 9600 8430 9628 9007
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 8760 7540 8812 7546
rect 8760 7482 8812 7488
rect 8852 6792 8904 6798
rect 8680 6740 8852 6746
rect 8680 6734 8904 6740
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6390 8524 6598
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5710 8340 6054
rect 8404 5914 8432 6258
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8588 5642 8616 6734
rect 8680 6718 8892 6734
rect 8680 5710 8708 6718
rect 8850 6624 8906 6633
rect 8850 6559 8906 6568
rect 8668 5704 8720 5710
rect 8668 5646 8720 5652
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8864 5302 8892 6559
rect 9586 5808 9642 5817
rect 9586 5743 9588 5752
rect 9640 5743 9642 5752
rect 9588 5714 9640 5720
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 5001 9628 5102
rect 9586 4992 9642 5001
rect 9586 4927 9642 4936
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 9036 4684 9088 4690
rect 9036 4626 9088 4632
rect 8220 4185 8248 4626
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4282 8340 4558
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8496 4214 8524 4422
rect 8484 4208 8536 4214
rect 8206 4176 8262 4185
rect 8484 4150 8536 4156
rect 8206 4111 8262 4120
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8404 3738 8432 4082
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8588 3398 8616 4490
rect 9048 3534 9076 4626
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8576 3392 8628 3398
rect 8390 3360 8446 3369
rect 8576 3334 8628 3340
rect 8390 3295 8446 3304
rect 8300 2984 8352 2990
rect 8128 2910 8248 2938
rect 8300 2926 8352 2932
rect 8116 2848 8168 2854
rect 8116 2790 8168 2796
rect 8128 2446 8156 2790
rect 8116 2440 8168 2446
rect 8116 2382 8168 2388
rect 7744 2276 7944 2300
rect 7744 2220 7776 2276
rect 7832 2220 7856 2276
rect 7912 2220 7944 2276
rect 8024 2304 8076 2310
rect 8024 2246 8076 2252
rect 8116 2304 8168 2310
rect 8116 2246 8168 2252
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7344 1900 7376 1956
rect 7432 1900 7456 1956
rect 7512 1900 7544 1956
rect 7344 1876 7544 1900
rect 7344 1820 7376 1876
rect 7432 1820 7456 1876
rect 7512 1820 7544 1876
rect 7344 1040 7544 1820
rect 7744 1040 7944 2220
rect 8036 1970 8064 2246
rect 8128 2038 8156 2246
rect 8116 2032 8168 2038
rect 8116 1974 8168 1980
rect 8024 1964 8076 1970
rect 8024 1906 8076 1912
rect 8220 1358 8248 2910
rect 8312 1834 8340 2926
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 8404 1426 8432 3295
rect 8588 3126 8616 3334
rect 9036 3188 9088 3194
rect 9036 3130 9088 3136
rect 8576 3120 8628 3126
rect 8576 3062 8628 3068
rect 8588 2446 8616 3062
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8668 2440 8720 2446
rect 8668 2382 8720 2388
rect 8588 2038 8616 2382
rect 8576 2032 8628 2038
rect 8576 1974 8628 1980
rect 8680 1970 8708 2382
rect 9048 2106 9076 3130
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8680 1494 8708 1906
rect 9588 1896 9640 1902
rect 9588 1838 9640 1844
rect 9600 1737 9628 1838
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 8668 1488 8720 1494
rect 8668 1430 8720 1436
rect 8392 1420 8444 1426
rect 8392 1362 8444 1368
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 6544 988 6744 1020
rect 9048 921 9076 1294
rect 9034 912 9090 921
rect 9034 847 9090 856
<< via2 >>
rect 1398 12552 1454 12608
rect 386 11736 442 11792
rect 1030 10920 1086 10976
rect 478 10124 534 10160
rect 478 10104 480 10124
rect 480 10104 532 10124
rect 532 10104 534 10124
rect 386 9288 442 9344
rect 938 7656 994 7712
rect 2134 11192 2190 11248
rect 1214 6840 1270 6896
rect 478 6024 534 6080
rect 386 5208 442 5264
rect 478 4392 534 4448
rect 2576 13100 2632 13156
rect 2656 13100 2712 13156
rect 2576 13020 2632 13076
rect 2656 13020 2712 13076
rect 2778 11464 2834 11520
rect 2410 10512 2466 10568
rect 3376 13900 3432 13956
rect 3456 13900 3512 13956
rect 3376 13820 3432 13876
rect 3456 13820 3512 13876
rect 2976 13500 3032 13556
rect 3056 13500 3112 13556
rect 2976 13420 3032 13476
rect 3056 13420 3112 13476
rect 3238 12008 3294 12064
rect 3606 12180 3608 12200
rect 3608 12180 3660 12200
rect 3660 12180 3662 12200
rect 3606 12144 3662 12180
rect 3776 10300 3832 10356
rect 3856 10300 3912 10356
rect 3776 10220 3832 10276
rect 3856 10220 3912 10276
rect 3376 9900 3432 9956
rect 3456 9900 3512 9956
rect 2976 9500 3032 9556
rect 3056 9500 3112 9556
rect 3376 9820 3432 9876
rect 3456 9820 3512 9876
rect 2976 9420 3032 9476
rect 3056 9420 3112 9476
rect 2576 9100 2632 9156
rect 2656 9100 2712 9156
rect 2576 9020 2632 9076
rect 2656 9020 2712 9076
rect 938 2760 994 2816
rect 386 2488 442 2544
rect 2576 5100 2632 5156
rect 2656 5100 2712 5156
rect 2576 5020 2632 5076
rect 2656 5020 2712 5076
rect 1950 2488 2006 2544
rect 932 2300 988 2356
rect 1012 2300 1068 2356
rect 932 2220 988 2276
rect 1012 2220 1068 2276
rect 386 1944 442 2000
rect 1532 1900 1588 1956
rect 1612 1900 1668 1956
rect 1532 1820 1588 1876
rect 1612 1820 1668 1876
rect 2976 5500 3032 5556
rect 3056 5500 3112 5556
rect 2976 5466 3032 5476
rect 3056 5466 3112 5476
rect 2976 5420 3006 5466
rect 3006 5420 3018 5466
rect 3018 5420 3032 5466
rect 3056 5420 3070 5466
rect 3070 5420 3082 5466
rect 3082 5420 3112 5466
rect 3376 5900 3432 5956
rect 3456 5900 3512 5956
rect 3376 5820 3432 5876
rect 3456 5820 3512 5876
rect 4250 11192 4306 11248
rect 4158 8472 4214 8528
rect 4986 10512 5042 10568
rect 3776 6300 3832 6356
rect 3856 6300 3912 6356
rect 3776 6220 3832 6276
rect 3856 6220 3912 6276
rect 5630 11872 5686 11928
rect 5630 11600 5686 11656
rect 5446 10784 5502 10840
rect 4250 3576 4306 3632
rect 4710 3576 4766 3632
rect 3776 2300 3832 2356
rect 3856 2300 3912 2356
rect 3776 2220 3832 2276
rect 3856 2220 3912 2276
rect 5906 11600 5962 11656
rect 5814 10784 5870 10840
rect 6976 13500 7032 13556
rect 7056 13500 7112 13556
rect 6976 13420 7032 13476
rect 7056 13420 7112 13476
rect 7376 13900 7432 13956
rect 7456 13900 7512 13956
rect 7376 13820 7432 13876
rect 7456 13820 7512 13876
rect 6576 13100 6632 13156
rect 6656 13100 6712 13156
rect 6576 13020 6632 13076
rect 6656 13020 6712 13076
rect 6366 11600 6422 11656
rect 5354 3440 5410 3496
rect 6826 12824 6882 12880
rect 7194 12824 7250 12880
rect 6576 9100 6632 9156
rect 6656 9100 6712 9156
rect 6576 9020 6632 9076
rect 6656 9020 6712 9076
rect 6976 9500 7032 9556
rect 7056 9500 7112 9556
rect 6976 9420 7032 9476
rect 7056 9420 7112 9476
rect 7376 9900 7432 9956
rect 7456 9900 7512 9956
rect 7376 9820 7432 9876
rect 7456 9820 7512 9876
rect 7194 8236 7196 8256
rect 7196 8236 7248 8256
rect 7248 8236 7250 8256
rect 7194 8200 7250 8236
rect 6576 5100 6632 5156
rect 6656 5100 6712 5156
rect 6576 5020 6632 5076
rect 6656 5020 6712 5076
rect 6976 5500 7032 5556
rect 7056 5500 7112 5556
rect 6976 5466 7032 5476
rect 7056 5466 7112 5476
rect 6976 5420 7006 5466
rect 7006 5420 7018 5466
rect 7018 5420 7032 5466
rect 7056 5420 7070 5466
rect 7070 5420 7082 5466
rect 7082 5420 7112 5466
rect 6458 3440 6514 3496
rect 5630 2488 5686 2544
rect 7776 10300 7832 10356
rect 7856 10300 7912 10356
rect 7776 10220 7832 10276
rect 7856 10220 7912 10276
rect 7376 5900 7432 5956
rect 7456 5900 7512 5956
rect 7376 5820 7432 5876
rect 7456 5820 7512 5876
rect 6576 1100 6632 1156
rect 6656 1100 6712 1156
rect 6576 1020 6632 1076
rect 6656 1020 6712 1076
rect 6976 1500 7032 1556
rect 7056 1500 7112 1556
rect 6976 1420 7032 1476
rect 7056 1420 7112 1476
rect 8114 10648 8170 10704
rect 7776 6300 7832 6356
rect 7856 6300 7912 6356
rect 7776 6220 7832 6276
rect 7856 6220 7912 6276
rect 7776 2300 7832 2356
rect 7856 2300 7912 2356
rect 8482 12280 8538 12336
rect 9586 13948 9588 13968
rect 9588 13948 9640 13968
rect 9640 13948 9642 13968
rect 9586 13912 9642 13948
rect 8666 12008 8722 12064
rect 8390 7384 8446 7440
rect 9586 13096 9642 13152
rect 9126 11464 9182 11520
rect 9586 9832 9642 9888
rect 9586 9016 9642 9072
rect 8850 6568 8906 6624
rect 9586 5772 9642 5808
rect 9586 5752 9588 5772
rect 9588 5752 9640 5772
rect 9640 5752 9642 5772
rect 9586 4936 9642 4992
rect 8206 4120 8262 4176
rect 8390 3304 8446 3360
rect 7776 2220 7832 2276
rect 7856 2220 7912 2276
rect 7376 1900 7432 1956
rect 7456 1900 7512 1956
rect 7376 1820 7432 1876
rect 7456 1820 7512 1876
rect 9586 1672 9642 1728
rect 9034 856 9090 912
<< metal3 >>
rect 596 13956 9432 13988
rect 9600 13973 10200 14000
rect 596 13900 3376 13956
rect 3432 13900 3456 13956
rect 3512 13900 7376 13956
rect 7432 13900 7456 13956
rect 7512 13900 9432 13956
rect 9581 13968 10200 13973
rect 9581 13912 9586 13968
rect 9642 13912 10200 13968
rect 9581 13907 10200 13912
rect 596 13876 9432 13900
rect 9600 13880 10200 13907
rect 596 13820 3376 13876
rect 3432 13820 3456 13876
rect 3512 13820 7376 13876
rect 7432 13820 7456 13876
rect 7512 13820 9432 13876
rect 596 13788 9432 13820
rect 596 13556 9432 13588
rect 596 13500 2976 13556
rect 3032 13500 3056 13556
rect 3112 13500 6976 13556
rect 7032 13500 7056 13556
rect 7112 13500 9432 13556
rect 596 13476 9432 13500
rect 596 13420 2976 13476
rect 3032 13420 3056 13476
rect 3112 13420 6976 13476
rect 7032 13420 7056 13476
rect 7112 13420 9432 13476
rect 596 13388 9432 13420
rect 596 13156 9432 13188
rect 9600 13157 10200 13184
rect 596 13100 2576 13156
rect 2632 13100 2656 13156
rect 2712 13100 6576 13156
rect 6632 13100 6656 13156
rect 6712 13100 9432 13156
rect 596 13076 9432 13100
rect 9581 13152 10200 13157
rect 9581 13096 9586 13152
rect 9642 13096 10200 13152
rect 9581 13091 10200 13096
rect 596 13020 2576 13076
rect 2632 13020 2656 13076
rect 2712 13020 6576 13076
rect 6632 13020 6656 13076
rect 6712 13020 9432 13076
rect 9600 13064 10200 13091
rect 596 12988 9432 13020
rect 6821 12882 6887 12885
rect 7189 12882 7255 12885
rect 6821 12880 7255 12882
rect 6821 12824 6826 12880
rect 6882 12824 7194 12880
rect 7250 12824 7255 12880
rect 6821 12822 7255 12824
rect 6821 12819 6887 12822
rect 7189 12819 7255 12822
rect -200 12610 400 12640
rect 1393 12610 1459 12613
rect -200 12608 1459 12610
rect -200 12552 1398 12608
rect 1454 12552 1459 12608
rect -200 12550 1459 12552
rect -200 12520 400 12550
rect 1393 12547 1459 12550
rect 8477 12338 8543 12341
rect 9600 12338 10200 12368
rect 8477 12336 10200 12338
rect 8477 12280 8482 12336
rect 8538 12280 10200 12336
rect 8477 12278 10200 12280
rect 8477 12275 8543 12278
rect 9600 12248 10200 12278
rect 3601 12202 3667 12205
rect 2822 12200 3667 12202
rect 2822 12144 3606 12200
rect 3662 12144 3667 12200
rect 2822 12142 3667 12144
rect -200 11797 400 11824
rect -200 11792 447 11797
rect -200 11736 386 11792
rect 442 11736 447 11792
rect -200 11731 447 11736
rect -200 11704 400 11731
rect 2822 11525 2882 12142
rect 3601 12139 3667 12142
rect 3233 12066 3299 12069
rect 8661 12066 8727 12069
rect 3233 12064 8727 12066
rect 3233 12008 3238 12064
rect 3294 12008 8666 12064
rect 8722 12008 8727 12064
rect 3233 12006 8727 12008
rect 3233 12003 3299 12006
rect 8661 12003 8727 12006
rect 5625 11930 5691 11933
rect 5582 11928 5691 11930
rect 5582 11872 5630 11928
rect 5686 11872 5691 11928
rect 5582 11867 5691 11872
rect 5582 11661 5642 11867
rect 5582 11656 5691 11661
rect 5582 11600 5630 11656
rect 5686 11600 5691 11656
rect 5582 11598 5691 11600
rect 5625 11595 5691 11598
rect 5901 11658 5967 11661
rect 6361 11658 6427 11661
rect 5901 11656 6427 11658
rect 5901 11600 5906 11656
rect 5962 11600 6366 11656
rect 6422 11600 6427 11656
rect 5901 11598 6427 11600
rect 5901 11595 5967 11598
rect 6361 11595 6427 11598
rect 2773 11520 2882 11525
rect 2773 11464 2778 11520
rect 2834 11464 2882 11520
rect 2773 11462 2882 11464
rect 9121 11522 9187 11525
rect 9600 11522 10200 11552
rect 9121 11520 10200 11522
rect 9121 11464 9126 11520
rect 9182 11464 10200 11520
rect 9121 11462 10200 11464
rect 2773 11459 2839 11462
rect 9121 11459 9187 11462
rect 9600 11432 10200 11462
rect 2129 11250 2195 11253
rect 4245 11250 4311 11253
rect 2129 11248 4311 11250
rect 2129 11192 2134 11248
rect 2190 11192 4250 11248
rect 4306 11192 4311 11248
rect 2129 11190 4311 11192
rect 2129 11187 2195 11190
rect 4245 11187 4311 11190
rect -200 10978 400 11008
rect 1025 10978 1091 10981
rect -200 10976 1091 10978
rect -200 10920 1030 10976
rect 1086 10920 1091 10976
rect -200 10918 1091 10920
rect -200 10888 400 10918
rect 1025 10915 1091 10918
rect 5441 10842 5507 10845
rect 5809 10842 5875 10845
rect 5441 10840 5875 10842
rect 5441 10784 5446 10840
rect 5502 10784 5814 10840
rect 5870 10784 5875 10840
rect 5441 10782 5875 10784
rect 5441 10779 5507 10782
rect 5809 10779 5875 10782
rect 8109 10706 8175 10709
rect 9600 10706 10200 10736
rect 8109 10704 10200 10706
rect 8109 10648 8114 10704
rect 8170 10648 10200 10704
rect 8109 10646 10200 10648
rect 8109 10643 8175 10646
rect 9600 10616 10200 10646
rect 2405 10570 2471 10573
rect 4981 10570 5047 10573
rect 2405 10568 5047 10570
rect 2405 10512 2410 10568
rect 2466 10512 4986 10568
rect 5042 10512 5047 10568
rect 2405 10510 5047 10512
rect 2405 10507 2471 10510
rect 4981 10507 5047 10510
rect 596 10356 9432 10388
rect 596 10300 3776 10356
rect 3832 10300 3856 10356
rect 3912 10300 7776 10356
rect 7832 10300 7856 10356
rect 7912 10300 9432 10356
rect 596 10276 9432 10300
rect 596 10220 3776 10276
rect 3832 10220 3856 10276
rect 3912 10220 7776 10276
rect 7832 10220 7856 10276
rect 7912 10220 9432 10276
rect -200 10162 400 10192
rect 596 10188 9432 10220
rect 473 10162 539 10165
rect -200 10160 539 10162
rect -200 10104 478 10160
rect 534 10104 539 10160
rect -200 10102 539 10104
rect -200 10072 400 10102
rect 473 10099 539 10102
rect 596 9956 9432 9988
rect 596 9900 3376 9956
rect 3432 9900 3456 9956
rect 3512 9900 7376 9956
rect 7432 9900 7456 9956
rect 7512 9900 9432 9956
rect 596 9876 9432 9900
rect 9600 9893 10200 9920
rect 596 9820 3376 9876
rect 3432 9820 3456 9876
rect 3512 9820 7376 9876
rect 7432 9820 7456 9876
rect 7512 9820 9432 9876
rect 9581 9888 10200 9893
rect 9581 9832 9586 9888
rect 9642 9832 10200 9888
rect 9581 9827 10200 9832
rect 596 9788 9432 9820
rect 9600 9800 10200 9827
rect 596 9556 9432 9588
rect 596 9500 2976 9556
rect 3032 9500 3056 9556
rect 3112 9500 6976 9556
rect 7032 9500 7056 9556
rect 7112 9500 9432 9556
rect 596 9476 9432 9500
rect 596 9420 2976 9476
rect 3032 9420 3056 9476
rect 3112 9420 6976 9476
rect 7032 9420 7056 9476
rect 7112 9420 9432 9476
rect 596 9388 9432 9420
rect -200 9349 400 9376
rect -200 9344 447 9349
rect -200 9288 386 9344
rect 442 9288 447 9344
rect -200 9283 447 9288
rect -200 9256 400 9283
rect 596 9156 9432 9188
rect 596 9100 2576 9156
rect 2632 9100 2656 9156
rect 2712 9100 6576 9156
rect 6632 9100 6656 9156
rect 6712 9100 9432 9156
rect 596 9076 9432 9100
rect 9600 9077 10200 9104
rect 596 9020 2576 9076
rect 2632 9020 2656 9076
rect 2712 9020 6576 9076
rect 6632 9020 6656 9076
rect 6712 9020 9432 9076
rect 596 8988 9432 9020
rect 9581 9072 10200 9077
rect 9581 9016 9586 9072
rect 9642 9016 10200 9072
rect 9581 9011 10200 9016
rect 9600 8984 10200 9011
rect -200 8530 400 8560
rect 4153 8530 4219 8533
rect -200 8528 4219 8530
rect -200 8472 4158 8528
rect 4214 8472 4219 8528
rect -200 8470 4219 8472
rect -200 8440 400 8470
rect 4153 8467 4219 8470
rect 7189 8258 7255 8261
rect 9600 8258 10200 8288
rect 7189 8256 10200 8258
rect 7189 8200 7194 8256
rect 7250 8200 10200 8256
rect 7189 8198 10200 8200
rect 7189 8195 7255 8198
rect 9600 8168 10200 8198
rect -200 7714 400 7744
rect 933 7714 999 7717
rect -200 7712 999 7714
rect -200 7656 938 7712
rect 994 7656 999 7712
rect -200 7654 999 7656
rect -200 7624 400 7654
rect 933 7651 999 7654
rect 8385 7442 8451 7445
rect 9600 7442 10200 7472
rect 8385 7440 10200 7442
rect 8385 7384 8390 7440
rect 8446 7384 10200 7440
rect 8385 7382 10200 7384
rect 8385 7379 8451 7382
rect 9600 7352 10200 7382
rect -200 6898 400 6928
rect 1209 6898 1275 6901
rect -200 6896 1275 6898
rect -200 6840 1214 6896
rect 1270 6840 1275 6896
rect -200 6838 1275 6840
rect -200 6808 400 6838
rect 1209 6835 1275 6838
rect 8845 6626 8911 6629
rect 9600 6626 10200 6656
rect 8845 6624 10200 6626
rect 8845 6568 8850 6624
rect 8906 6568 10200 6624
rect 8845 6566 10200 6568
rect 8845 6563 8911 6566
rect 9600 6536 10200 6566
rect 596 6356 9432 6388
rect 596 6300 3776 6356
rect 3832 6300 3856 6356
rect 3912 6300 7776 6356
rect 7832 6300 7856 6356
rect 7912 6300 9432 6356
rect 596 6276 9432 6300
rect 596 6220 3776 6276
rect 3832 6220 3856 6276
rect 3912 6220 7776 6276
rect 7832 6220 7856 6276
rect 7912 6220 9432 6276
rect 596 6188 9432 6220
rect -200 6082 400 6112
rect 473 6082 539 6085
rect -200 6080 539 6082
rect -200 6024 478 6080
rect 534 6024 539 6080
rect -200 6022 539 6024
rect -200 5992 400 6022
rect 473 6019 539 6022
rect 596 5956 9432 5988
rect 596 5900 3376 5956
rect 3432 5900 3456 5956
rect 3512 5900 7376 5956
rect 7432 5900 7456 5956
rect 7512 5900 9432 5956
rect 596 5876 9432 5900
rect 596 5820 3376 5876
rect 3432 5820 3456 5876
rect 3512 5820 7376 5876
rect 7432 5820 7456 5876
rect 7512 5820 9432 5876
rect 596 5788 9432 5820
rect 9600 5813 10200 5840
rect 9581 5808 10200 5813
rect 9581 5752 9586 5808
rect 9642 5752 10200 5808
rect 9581 5747 10200 5752
rect 9600 5720 10200 5747
rect 596 5556 9432 5588
rect 596 5500 2976 5556
rect 3032 5500 3056 5556
rect 3112 5500 6976 5556
rect 7032 5500 7056 5556
rect 7112 5500 9432 5556
rect 596 5476 9432 5500
rect 596 5420 2976 5476
rect 3032 5420 3056 5476
rect 3112 5420 6976 5476
rect 7032 5420 7056 5476
rect 7112 5420 9432 5476
rect 596 5388 9432 5420
rect -200 5269 400 5296
rect -200 5264 447 5269
rect -200 5208 386 5264
rect 442 5208 447 5264
rect -200 5203 447 5208
rect -200 5176 400 5203
rect 596 5156 9432 5188
rect 596 5100 2576 5156
rect 2632 5100 2656 5156
rect 2712 5100 6576 5156
rect 6632 5100 6656 5156
rect 6712 5100 9432 5156
rect 596 5076 9432 5100
rect 596 5020 2576 5076
rect 2632 5020 2656 5076
rect 2712 5020 6576 5076
rect 6632 5020 6656 5076
rect 6712 5020 9432 5076
rect 596 4988 9432 5020
rect 9600 4997 10200 5024
rect 9581 4992 10200 4997
rect 9581 4936 9586 4992
rect 9642 4936 10200 4992
rect 9581 4931 10200 4936
rect 9600 4904 10200 4931
rect -200 4450 400 4480
rect 473 4450 539 4453
rect -200 4448 539 4450
rect -200 4392 478 4448
rect 534 4392 539 4448
rect -200 4390 539 4392
rect -200 4360 400 4390
rect 473 4387 539 4390
rect 8201 4178 8267 4181
rect 9600 4178 10200 4208
rect 8201 4176 10200 4178
rect 8201 4120 8206 4176
rect 8262 4120 10200 4176
rect 8201 4118 10200 4120
rect 8201 4115 8267 4118
rect 9600 4088 10200 4118
rect -200 3634 400 3664
rect 4245 3634 4311 3637
rect 4705 3634 4771 3637
rect -200 3632 4771 3634
rect -200 3576 4250 3632
rect 4306 3576 4710 3632
rect 4766 3576 4771 3632
rect -200 3574 4771 3576
rect -200 3544 400 3574
rect 4245 3571 4311 3574
rect 4705 3571 4771 3574
rect 5349 3498 5415 3501
rect 6453 3498 6519 3501
rect 5349 3496 6519 3498
rect 5349 3440 5354 3496
rect 5410 3440 6458 3496
rect 6514 3440 6519 3496
rect 5349 3438 6519 3440
rect 5349 3435 5415 3438
rect 6453 3435 6519 3438
rect 8385 3362 8451 3365
rect 9600 3362 10200 3392
rect 8385 3360 10200 3362
rect 8385 3304 8390 3360
rect 8446 3304 10200 3360
rect 8385 3302 10200 3304
rect 8385 3299 8451 3302
rect 9600 3272 10200 3302
rect -200 2818 400 2848
rect 933 2818 999 2821
rect -200 2816 999 2818
rect -200 2760 938 2816
rect 994 2760 999 2816
rect -200 2758 999 2760
rect -200 2728 400 2758
rect 933 2755 999 2758
rect 381 2546 447 2549
rect 1945 2546 2011 2549
rect 381 2544 2011 2546
rect 381 2488 386 2544
rect 442 2488 1950 2544
rect 2006 2488 2011 2544
rect 381 2486 2011 2488
rect 381 2483 447 2486
rect 1945 2483 2011 2486
rect 5625 2546 5691 2549
rect 9600 2546 10200 2576
rect 5625 2544 10200 2546
rect 5625 2488 5630 2544
rect 5686 2488 10200 2544
rect 5625 2486 10200 2488
rect 5625 2483 5691 2486
rect 9600 2456 10200 2486
rect 596 2356 9432 2388
rect 596 2300 932 2356
rect 988 2300 1012 2356
rect 1068 2300 3776 2356
rect 3832 2300 3856 2356
rect 3912 2300 7776 2356
rect 7832 2300 7856 2356
rect 7912 2300 9432 2356
rect 596 2276 9432 2300
rect 596 2220 932 2276
rect 988 2220 1012 2276
rect 1068 2220 3776 2276
rect 3832 2220 3856 2276
rect 3912 2220 7776 2276
rect 7832 2220 7856 2276
rect 7912 2220 9432 2276
rect 596 2188 9432 2220
rect -200 2005 400 2032
rect -200 2000 447 2005
rect -200 1944 386 2000
rect 442 1944 447 2000
rect -200 1939 447 1944
rect 596 1956 9432 1988
rect -200 1912 400 1939
rect 596 1900 1532 1956
rect 1588 1900 1612 1956
rect 1668 1900 7376 1956
rect 7432 1900 7456 1956
rect 7512 1900 9432 1956
rect 596 1876 9432 1900
rect 596 1820 1532 1876
rect 1588 1820 1612 1876
rect 1668 1820 7376 1876
rect 7432 1820 7456 1876
rect 7512 1820 9432 1876
rect 596 1788 9432 1820
rect 9600 1733 10200 1760
rect 9581 1728 10200 1733
rect 9581 1672 9586 1728
rect 9642 1672 10200 1728
rect 9581 1667 10200 1672
rect 9600 1640 10200 1667
rect 596 1556 9432 1588
rect 596 1500 6976 1556
rect 7032 1500 7056 1556
rect 7112 1500 9432 1556
rect 596 1476 9432 1500
rect 596 1420 6976 1476
rect 7032 1420 7056 1476
rect 7112 1420 9432 1476
rect 596 1388 9432 1420
rect 596 1156 9432 1188
rect 596 1100 6576 1156
rect 6632 1100 6656 1156
rect 6712 1100 9432 1156
rect 596 1076 9432 1100
rect 596 1020 6576 1076
rect 6632 1020 6656 1076
rect 6712 1020 9432 1076
rect 596 988 9432 1020
rect 9029 914 9095 917
rect 9600 914 10200 944
rect 9029 912 10200 914
rect 9029 856 9034 912
rect 9090 856 10200 912
rect 9029 854 10200 856
rect 9029 851 9095 854
rect 9600 824 10200 854
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1562557784
transform -1 0 6900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1562557784
transform -1 0 3588 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _059_
timestamp 21601
transform -1 0 8924 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _060_
timestamp 21601
transform 1 0 8556 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _061_
timestamp 21601
transform -1 0 7912 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _062_
timestamp 21601
transform 1 0 6072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _063_
timestamp 21601
transform -1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _064_
timestamp 21601
transform 1 0 6808 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _065_
timestamp 21601
transform -1 0 5796 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _066_
timestamp 21601
transform -1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _067_
timestamp 21601
transform -1 0 6348 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _068_
timestamp 21601
transform 1 0 3496 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _069_
timestamp 21601
transform -1 0 8924 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _070_
timestamp 21601
transform 1 0 6808 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _071_
timestamp 21601
transform -1 0 5704 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _072_
timestamp 21601
transform -1 0 2944 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _073_
timestamp 21601
transform -1 0 1840 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 21601
transform -1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _075_
timestamp 21601
transform -1 0 1564 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _076_
timestamp 21601
transform -1 0 3220 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _077_
timestamp 21601
transform -1 0 4324 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _078_
timestamp 21601
transform -1 0 6348 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _079_
timestamp 21601
transform 1 0 8464 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _080_
timestamp 21601
transform -1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _081_
timestamp 21601
transform 1 0 3496 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _082_
timestamp 21601
transform -1 0 8924 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _083_
timestamp 21601
transform -1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _084_
timestamp 21601
transform 1 0 8648 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _085_
timestamp 21601
transform -1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _086_
timestamp 21601
transform 1 0 5612 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _087_
timestamp 21601
transform 1 0 8464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _088_
timestamp 21601
transform -1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _089_
timestamp 21601
transform 1 0 7912 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _090_
timestamp 21601
transform 1 0 8464 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1562557784
transform -1 0 7544 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1562557784
transform 1 0 6072 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 1562557784
transform 1 0 5244 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1562557784
transform 1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1562557784
transform 1 0 5888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1562557784
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1562557784
transform -1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1562557784
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1562557784
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1562557784
transform 1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1562557784
transform 1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1562557784
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _103_
timestamp 1562557784
transform 1 0 1012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _104_
timestamp 21601
transform 1 0 1288 0 -1 8704
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _105_
timestamp 21601
transform 1 0 3404 0 1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _106_
timestamp 21601
transform 1 0 5980 0 1 2176
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _107_
timestamp 21601
transform 1 0 6348 0 -1 11968
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _108_
timestamp 21601
transform 1 0 3220 0 -1 13056
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _109_
timestamp 21601
transform 1 0 4692 0 1 11968
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 21601
transform 1 0 6532 0 -1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 21601
transform -1 0 7636 0 -1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 21601
transform 1 0 6532 0 -1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 21601
transform 1 0 4508 0 1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 21601
transform 1 0 6164 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 21601
transform 1 0 6532 0 -1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _116_
timestamp 21601
transform 1 0 6532 0 -1 13056
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_1  _117_
timestamp 21601
transform 1 0 920 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _118_
timestamp 21601
transform 1 0 920 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _119_
timestamp 21601
transform 1 0 1932 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp 21601
transform -1 0 3220 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _121_
timestamp 21601
transform 1 0 2760 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _122_
timestamp 21601
transform -1 0 5060 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _123_
timestamp 21601
transform 1 0 3864 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _124_
timestamp 21601
transform 1 0 4784 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _125_
timestamp 21601
transform 1 0 3772 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _126_
timestamp 21601
transform -1 0 5796 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _127_
timestamp 21601
transform -1 0 6716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 21601
transform 1 0 4876 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 21601
transform 1 0 5888 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 21601
transform -1 0 6808 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 21601
transform -1 0 5152 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _132_
timestamp 21601
transform 1 0 3956 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfbbn_2  _133_
timestamp 21601
transform 1 0 6348 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_1  _134_
timestamp 21601
transform -1 0 2760 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp 21601
transform -1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[0\]
timestamp 21601
transform -1 0 1932 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[1\]
timestamp 21601
transform -1 0 1932 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[2\]
timestamp 21601
transform -1 0 1932 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 21601
transform 1 0 6072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout40
timestamp 21601
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 21601
transform 1 0 5520 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 21601
transform -1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 21601
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23
timestamp 21601
transform 1 0 2760 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 21601
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 21601
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 21601
transform 1 0 3588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp 21601
transform 1 0 3864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp 21601
transform 1 0 4140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp 21601
transform 1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp 21601
transform 1 0 4692 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 21601
transform 1 0 4968 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49
timestamp 21601
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52
timestamp 21601
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55
timestamp 21601
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 21601
transform 1 0 5980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77
timestamp 21601
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80
timestamp 21601
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_83
timestamp 21601
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_86
timestamp 21601
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_23
timestamp 21601
transform 1 0 2760 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_26
timestamp 21601
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_29
timestamp 21601
transform 1 0 3312 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 21601
transform 1 0 6716 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 21601
transform 1 0 7544 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_77
timestamp 21601
transform 1 0 7728 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_80
timestamp 21601
transform 1 0 8004 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_83
timestamp 21601
transform 1 0 8280 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_86
timestamp 21601
transform 1 0 8556 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 21601
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_31
timestamp 21601
transform 1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_34
timestamp 21601
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp 21601
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_40
timestamp 21601
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 21601
transform 1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 21601
transform 1 0 5888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 21601
transform 1 0 9016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_23
timestamp 21601
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_26
timestamp 21601
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_29
timestamp 21601
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 21601
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 21601
transform 1 0 920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp 21601
transform 1 0 1196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp 21601
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp 21601
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp 21601
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp 21601
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_21
timestamp 21601
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp 21601
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 21601
transform 1 0 3128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 21601
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp 21601
transform 1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_35
timestamp 21601
transform 1 0 3864 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_80
timestamp 21601
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 21601
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 21601
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp 21601
transform 1 0 1196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp 21601
transform 1 0 1472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp 21601
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 21601
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp 21601
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp 21601
transform 1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp 21601
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 21601
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp 21601
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_33
timestamp 21601
transform 1 0 3680 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_54
timestamp 21601
transform 1 0 5612 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 21601
transform 1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 21601
transform 1 0 6440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 21601
transform 1 0 920 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_10
timestamp 21601
transform 1 0 1564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_17
timestamp 21601
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_20
timestamp 21601
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_23
timestamp 21601
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 21601
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 21601
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp 21601
transform 1 0 3588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp 21601
transform 1 0 3864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 21601
transform 1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 21601
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_23
timestamp 21601
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_26
timestamp 21601
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_29
timestamp 21601
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_32
timestamp 21601
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_35
timestamp 21601
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_38
timestamp 21601
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_41
timestamp 21601
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_44
timestamp 21601
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_47
timestamp 21601
transform 1 0 4968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 21601
transform 1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_19
timestamp 21601
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_22
timestamp 21601
transform 1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 21601
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 21601
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 21601
transform 1 0 3588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp 21601
transform 1 0 3864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp 21601
transform 1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 21601
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_44
timestamp 21601
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 21601
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp 21601
transform 1 0 1196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp 21601
transform 1 0 1472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_12
timestamp 21601
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp 21601
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp 21601
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp 21601
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_24
timestamp 21601
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 21601
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp 21601
transform 1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_33
timestamp 21601
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 21601
transform 1 0 5704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 21601
transform 1 0 5888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 21601
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp 21601
transform 1 0 1196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp 21601
transform 1 0 1472 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp 21601
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp 21601
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp 21601
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp 21601
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_24
timestamp 21601
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 21601
transform 1 0 3128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 21601
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 21601
transform 1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_35
timestamp 21601
transform 1 0 3864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 21601
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 21601
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_80
timestamp 21601
transform 1 0 8004 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 21601
transform 1 0 8280 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 21601
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_9
timestamp 21601
transform 1 0 1472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_12
timestamp 21601
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 21601
transform 1 0 2024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_25
timestamp 21601
transform 1 0 2944 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_48
timestamp 21601
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_91
timestamp 21601
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 21601
transform 1 0 920 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_22
timestamp 21601
transform 1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 21601
transform 1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 21601
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 21601
transform 1 0 3588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_35
timestamp 21601
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_45
timestamp 21601
transform 1 0 4784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_48
timestamp 21601
transform 1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_51
timestamp 21601
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 21601
transform 1 0 6808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 21601
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 21601
transform 1 0 920 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_40
timestamp 21601
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_43
timestamp 21601
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_46
timestamp 21601
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_49
timestamp 21601
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_52
timestamp 21601
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 21601
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 21601
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 21601
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 21601
transform 1 0 2392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_32
timestamp 21601
transform 1 0 3588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_43
timestamp 21601
transform 1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_46
timestamp 21601
transform 1 0 4876 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_72
timestamp 21601
transform 1 0 7268 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 21601
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_23
timestamp 21601
transform 1 0 2760 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_57
timestamp 21601
transform 1 0 5888 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 21601
transform 1 0 8924 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 21601
transform 1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_49
timestamp 21601
transform 1 0 5152 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 21601
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 21601
transform 1 0 5704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 21601
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_14
timestamp 21601
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 21601
transform 1 0 3312 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_58
timestamp 21601
transform 1 0 5980 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 21601
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 21601
transform 1 0 4600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 21601
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 21601
transform 1 0 920 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 21601
transform 1 0 3312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 21601
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 21601
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_19
timestamp 21601
transform 1 0 2392 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 21601
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 21601
transform 1 0 920 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 21601
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 21601
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 21601
transform 1 0 920 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 21601
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  gpio_control_block_44
timestamp 1562557784
transform 1 0 6440 0 -1 8704
box -38 -48 314 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 600 0 1 1252
box 0 0 1 1
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 21601
transform -1 0 3220 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 21601
transform -1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 21601
transform 1 0 1748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 21601
transform -1 0 5428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 21601
transform 1 0 1012 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 21601
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 21601
transform 1 0 1012 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 21601
transform -1 0 4692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 21601
transform 1 0 1748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 21601
transform -1 0 4324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 21601
transform -1 0 4692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 21601
transform -1 0 6624 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 21601
transform 1 0 4140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 21601
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 21601
transform -1 0 3220 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 21601
transform 1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 21601
transform -1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 21601
transform 1 0 4048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 21601
transform 1 0 5888 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 21601
transform 1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 21601
transform -1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 21601
transform 1 0 6716 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 21601
transform 1 0 6164 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 21601
transform 1 0 5152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 21601
transform 1 0 4784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 21601
transform -1 0 2944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 21601
transform -1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 21601
transform 1 0 5060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 21601
transform -1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 21601
transform 1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 21601
transform 1 0 2852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 21601
transform -1 0 3680 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 21601
transform -1 0 4600 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 21601
transform -1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 21601
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 21601
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 21601
transform 1 0 8740 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 21601
transform -1 0 6440 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 21601
transform -1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 21601
transform 1 0 3128 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 21601
transform 1 0 3312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 21601
transform -1 0 2392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 21601
transform -1 0 1472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 21601
transform -1 0 1196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 21601
transform -1 0 9108 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 21601
transform -1 0 1196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 21601
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 21601
transform -1 0 1196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 21601
transform 1 0 920 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 21601
transform 1 0 6164 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 21601
transform -1 0 8372 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 21601
transform -1 0 8372 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 21601
transform -1 0 8372 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 21601
transform -1 0 5060 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 21601
transform -1 0 8372 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 21601
transform 1 0 6900 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 21601
transform -1 0 9108 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 21601
transform -1 0 6900 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 21601
transform 1 0 7636 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 21601
transform 1 0 6900 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 21601
transform 1 0 4324 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output34
timestamp 21601
transform 1 0 6164 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output35
timestamp 21601
transform -1 0 4876 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output36
timestamp 21601
transform -1 0 8372 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output37
timestamp 21601
transform 1 0 920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 21601
transform -1 0 2392 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Left_3
timestamp 21601
transform 1 0 2484 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Right_27
timestamp 21601
transform -1 0 9384 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Left_0
timestamp 21601
transform 1 0 2484 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Right_4
timestamp 21601
transform -1 0 9384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Left_1
timestamp 21601
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Right_5
timestamp 21601
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Left_2
timestamp 21601
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Right_6
timestamp 21601
transform -1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_28
timestamp 21601
transform 1 0 644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_7
timestamp 21601
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_29
timestamp 21601
transform 1 0 644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_8
timestamp 21601
transform -1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_30
timestamp 21601
transform 1 0 644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_9
timestamp 21601
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_31
timestamp 21601
transform 1 0 644 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_10
timestamp 21601
transform -1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_32
timestamp 21601
transform 1 0 644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_11
timestamp 21601
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_33
timestamp 21601
transform 1 0 644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_12
timestamp 21601
transform -1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_34
timestamp 21601
transform 1 0 644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_13
timestamp 21601
transform -1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_35
timestamp 21601
transform 1 0 644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_14
timestamp 21601
transform -1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_36
timestamp 21601
transform 1 0 644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_15
timestamp 21601
transform -1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_37
timestamp 21601
transform 1 0 644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_16
timestamp 21601
transform -1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_38
timestamp 21601
transform 1 0 644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_17
timestamp 21601
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_39
timestamp 21601
transform 1 0 644 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_18
timestamp 21601
transform -1 0 9384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_40
timestamp 21601
transform 1 0 644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_19
timestamp 21601
transform -1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_41
timestamp 21601
transform 1 0 644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_20
timestamp 21601
transform -1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_42
timestamp 21601
transform 1 0 644 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_21
timestamp 21601
transform -1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_43
timestamp 21601
transform 1 0 644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_22
timestamp 21601
transform -1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_44
timestamp 21601
transform 1 0 644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_23
timestamp 21601
transform -1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_45
timestamp 21601
transform 1 0 644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_24
timestamp 21601
transform -1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_46
timestamp 21601
transform 1 0 644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_25
timestamp 21601
transform -1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_47
timestamp 21601
transform 1 0 644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_26
timestamp 21601
transform -1 0 9384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_2_84
timestamp 21601
transform 1 0 5060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_2_85
timestamp 21601
transform 1 0 7636 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_2_48
timestamp 21601
transform 1 0 7636 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_2_49
timestamp 21601
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_2_50
timestamp 21601
transform 1 0 7636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_51
timestamp 21601
transform 1 0 3220 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_52
timestamp 21601
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_53
timestamp 21601
transform 1 0 8372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_54
timestamp 21601
transform 1 0 5796 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp 21601
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_56
timestamp 21601
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_57
timestamp 21601
transform 1 0 5796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_58
timestamp 21601
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_59
timestamp 21601
transform 1 0 8372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_60
timestamp 21601
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_61
timestamp 21601
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_62
timestamp 21601
transform 1 0 8372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_63
timestamp 21601
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_64
timestamp 21601
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_65
timestamp 21601
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_66
timestamp 21601
transform 1 0 5796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_67
timestamp 21601
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_68
timestamp 21601
transform 1 0 8372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_69
timestamp 21601
transform 1 0 5796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_70
timestamp 21601
transform 1 0 3220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_71
timestamp 21601
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_72
timestamp 21601
transform 1 0 5796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_73
timestamp 21601
transform 1 0 3220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_74
timestamp 21601
transform 1 0 8372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_75
timestamp 21601
transform 1 0 5796 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_76
timestamp 21601
transform 1 0 3220 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_77
timestamp 21601
transform 1 0 8372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_78
timestamp 21601
transform 1 0 5796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_79
timestamp 21601
transform 1 0 3220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_80
timestamp 21601
transform 1 0 8372 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_81
timestamp 21601
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_82
timestamp 21601
transform 1 0 5796 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_83
timestamp 21601
transform 1 0 8372 0 -1 14144
box -38 -48 130 592
<< labels >>
flabel metal2 s 5078 14400 5134 15000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 7838 14400 7894 15000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 8114 14400 8170 15000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 8390 14400 8446 15000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 8666 14400 8722 15000 0 FreeSans 224 90 0 0 gpio_defaults[13]
port 4 nsew signal input
flabel metal2 s 8942 14400 8998 15000 0 FreeSans 224 90 0 0 gpio_defaults[14]
port 5 nsew signal input
flabel metal2 s 9218 14400 9274 15000 0 FreeSans 224 90 0 0 gpio_defaults[15]
port 6 nsew signal input
flabel metal2 s 5354 14400 5410 15000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 7 nsew signal input
flabel metal2 s 5630 14400 5686 15000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 8 nsew signal input
flabel metal2 s 5906 14400 5962 15000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 9 nsew signal input
flabel metal2 s 6182 14400 6238 15000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 10 nsew signal input
flabel metal2 s 6458 14400 6514 15000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 11 nsew signal input
flabel metal2 s 6734 14400 6790 15000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 12 nsew signal input
flabel metal2 s 7010 14400 7066 15000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 13 nsew signal input
flabel metal2 s 7286 14400 7342 15000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 14 nsew signal input
flabel metal2 s 7562 14400 7618 15000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 15 nsew signal input
flabel metal3 s -200 5176 400 5296 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 16 nsew signal output
flabel metal3 s -200 6808 400 6928 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 17 nsew signal input
flabel metal3 s -200 5992 400 6112 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 18 nsew signal input
flabel metal3 s 9600 3272 10200 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 19 nsew signal output
flabel metal3 s 9600 5720 10200 5840 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 20 nsew signal output
flabel metal3 s 9600 7352 10200 7472 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 21 nsew signal output
flabel metal3 s 9600 4088 10200 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 22 nsew signal output
flabel metal3 s 9600 2456 10200 2576 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 23 nsew signal output
flabel metal3 s 9600 9800 10200 9920 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 24 nsew signal output
flabel metal3 s 9600 10616 10200 10736 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 25 nsew signal output
flabel metal3 s 9600 8984 10200 9104 0 FreeSans 480 0 0 0 pad_gpio_hys_trim
port 26 nsew signal output
flabel metal3 s 9600 13064 10200 13184 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 27 nsew signal output
flabel metal3 s 9600 824 10200 944 0 FreeSans 480 0 0 0 pad_gpio_in
port 28 nsew signal input
flabel metal3 s 9600 6536 10200 6656 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 29 nsew signal output
flabel metal3 s 9600 11432 10200 11552 0 FreeSans 480 0 0 0 pad_gpio_out
port 30 nsew signal output
flabel metal3 s 9600 13880 10200 14000 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 31 nsew signal output
flabel metal3 s 9600 4904 10200 5024 0 FreeSans 480 0 0 0 pad_gpio_slew_ctl[0]
port 32 nsew signal output
flabel metal3 s 9600 8168 10200 8288 0 FreeSans 480 0 0 0 pad_gpio_slew_ctl[1]
port 33 nsew signal output
flabel metal3 s 9600 1640 10200 1760 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 34 nsew signal output
flabel metal3 s 9600 12248 10200 12368 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 35 nsew signal output
flabel metal3 s -200 1912 400 2032 0 FreeSans 480 0 0 0 resetn
port 36 nsew signal input
flabel metal3 s -200 10072 400 10192 0 FreeSans 480 0 0 0 resetn_out
port 37 nsew signal output
flabel metal3 s -200 2728 400 2848 0 FreeSans 480 0 0 0 serial_clock
port 38 nsew signal input
flabel metal3 s -200 10888 400 11008 0 FreeSans 480 0 0 0 serial_clock_out
port 39 nsew signal output
flabel metal3 s -200 4360 400 4480 0 FreeSans 480 0 0 0 serial_data_in
port 40 nsew signal input
flabel metal3 s -200 12520 400 12640 0 FreeSans 480 0 0 0 serial_data_out
port 41 nsew signal output
flabel metal3 s -200 3544 400 3664 0 FreeSans 480 0 0 0 serial_load
port 42 nsew signal input
flabel metal3 s -200 11704 400 11824 0 FreeSans 480 0 0 0 serial_load_out
port 43 nsew signal output
flabel metal3 s -200 9256 400 9376 0 FreeSans 480 0 0 0 user_gpio_in
port 44 nsew signal output
flabel metal3 s -200 8440 400 8560 0 FreeSans 480 0 0 0 user_gpio_oeb
port 45 nsew signal input
flabel metal3 s -200 7624 400 7744 0 FreeSans 480 0 0 0 user_gpio_out
port 46 nsew signal input
flabel metal2 s 2544 4094 2744 14192 0 FreeSans 896 90 0 0 vccd
port 47 nsew power bidirectional
flabel metal2 s 6544 988 6744 14192 0 FreeSans 896 90 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 988 9432 1188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 4988 9432 5188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 8988 9432 9188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 12988 9432 13188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal2 s 3344 4094 3544 14192 0 FreeSans 896 90 0 0 vccd1
port 48 nsew power bidirectional
flabel metal2 s 7344 1040 7544 14192 0 FreeSans 896 90 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 1788 9432 1988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 5788 9432 5988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 9788 9432 9988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 13788 9432 13988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal2 s 2944 4094 3144 14192 0 FreeSans 896 90 0 0 vssd
port 49 nsew ground bidirectional
flabel metal2 s 6944 1040 7144 14192 0 FreeSans 896 90 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 1388 9432 1588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 5388 9432 5588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 9388 9432 9588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 13388 9432 13588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal2 s 3744 1040 3944 14192 0 FreeSans 896 90 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal2 s 7744 1040 7944 14192 0 FreeSans 896 90 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal3 s 596 2188 9432 2388 0 FreeSans 960 0 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal3 s 596 6188 9432 6388 0 FreeSans 960 0 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal3 s 596 10188 9432 10388 0 FreeSans 960 0 0 0 vssd1
port 50 nsew ground bidirectional
rlabel metal1 5934 2720 5934 2720 0 vccd
rlabel via2 1640 1928 1640 1928 0 vccd1
rlabel metal1 5934 2176 5934 2176 0 vssd
rlabel via2 1040 2328 1040 2328 0 vssd1
rlabel metal1 3542 8466 3542 8466 0 _000_
rlabel metal2 2438 8670 2438 8670 0 _001_
rlabel metal1 5290 11152 5290 11152 0 _002_
rlabel metal1 5106 10778 5106 10778 0 _003_
rlabel metal1 8004 2414 8004 2414 0 _004_
rlabel metal1 6946 1734 6946 1734 0 _005_
rlabel metal2 8234 12444 8234 12444 0 _006_
rlabel metal1 8195 11798 8195 11798 0 _007_
rlabel metal2 5106 13022 5106 13022 0 _008_
rlabel metal1 4048 12342 4048 12342 0 _009_
rlabel metal1 7038 12206 7038 12206 0 _010_
rlabel metal2 6118 12376 6118 12376 0 _011_
rlabel metal1 8464 3706 8464 3706 0 _012_
rlabel metal1 8287 4182 8287 4182 0 _013_
rlabel metal2 9062 2618 9062 2618 0 _014_
rlabel metal1 7820 2618 7820 2618 0 _015_
rlabel metal2 8510 10812 8510 10812 0 _016_
rlabel metal1 8372 10166 8372 10166 0 _017_
rlabel metal2 6394 7242 6394 7242 0 _018_
rlabel metal2 5566 6936 5566 6936 0 _019_
rlabel metal2 8050 7548 8050 7548 0 _020_
rlabel metal1 7452 8806 7452 8806 0 _021_
rlabel metal1 8464 5882 8464 5882 0 _022_
rlabel metal1 8287 6358 8287 6358 0 _023_
rlabel metal2 8372 12818 8372 12818 0 _024_
rlabel metal1 6854 12954 6854 12954 0 _025_
rlabel metal2 8878 9350 8878 9350 0 _026_
rlabel metal2 7682 9384 7682 9384 0 _027_
rlabel metal1 6624 10234 6624 10234 0 _028_
rlabel metal1 7544 2074 7544 2074 0 _029_
rlabel metal1 6302 9486 6302 9486 0 _030_
rlabel metal1 6302 12750 6302 12750 0 _031_
rlabel metal1 6486 6222 6486 6222 0 _032_
rlabel metal1 6118 7310 6118 7310 0 _033_
rlabel metal1 4462 6766 4462 6766 0 _034_
rlabel metal1 7360 3706 7360 3706 0 _035_
rlabel metal1 3910 11322 3910 11322 0 _036_
rlabel metal1 2254 12410 2254 12410 0 _037_
rlabel metal1 6394 11798 6394 11798 0 _038_
rlabel metal1 5474 2482 5474 2482 0 _039_
rlabel metal1 3358 11186 3358 11186 0 _040_
rlabel metal1 1242 8398 1242 8398 0 _041_
rlabel metal1 3634 11526 3634 11526 0 _042_
rlabel metal1 1150 13974 1150 13974 0 gpio_defaults[0]
rlabel metal1 4278 13940 4278 13940 0 gpio_defaults[10]
rlabel metal1 6578 13804 6578 13804 0 gpio_defaults[11]
rlabel metal2 3266 14110 3266 14110 0 gpio_defaults[12]
rlabel metal2 9016 12716 9016 12716 0 gpio_defaults[13]
rlabel metal2 5382 12580 5382 12580 0 gpio_defaults[15]
rlabel metal1 7774 12206 7774 12206 0 gpio_defaults[2]
rlabel metal1 3404 13362 3404 13362 0 gpio_defaults[3]
rlabel metal1 2323 13294 2323 13294 0 gpio_defaults[4]
rlabel metal2 1150 13804 1150 13804 0 gpio_defaults[5]
rlabel metal1 4738 12274 4738 12274 0 gpio_defaults[6]
rlabel metal1 1886 13804 1886 13804 0 gpio_defaults[7]
rlabel metal2 4646 13838 4646 13838 0 gpio_defaults[8]
rlabel metal1 6302 13362 6302 13362 0 gpio_defaults[9]
rlabel metal1 1801 1530 1801 1530 0 gpio_logic1
rlabel metal1 7544 5678 7544 5678 0 gpio_slew_ctl
rlabel metal1 1656 7922 1656 7922 0 mgmt_ena
rlabel metal3 360 5236 360 5236 0 mgmt_gpio_in
rlabel metal3 774 6868 774 6868 0 mgmt_gpio_oeb
rlabel metal3 406 6052 406 6052 0 mgmt_gpio_out
rlabel metal1 3542 9078 3542 9078 0 net1
rlabel metal2 5658 8058 5658 8058 0 net10
rlabel viali 6946 8942 6946 8942 0 net11
rlabel metal1 4002 8500 4002 8500 0 net12
rlabel metal1 4370 13770 4370 13770 0 net13
rlabel metal2 3266 11645 3266 11645 0 net14
rlabel metal2 1426 7599 1426 7599 0 net15
rlabel metal2 1150 7140 1150 7140 0 net16
rlabel metal2 1334 3536 1334 3536 0 net17
rlabel metal1 1196 3978 1196 3978 0 net18
rlabel metal2 1426 7922 1426 7922 0 net19
rlabel metal1 8970 3502 8970 3502 0 net2
rlabel metal1 1150 7480 1150 7480 0 net20
rlabel metal2 1150 5236 1150 5236 0 net21
rlabel metal1 7314 1326 7314 1326 0 net22
rlabel metal2 8326 5882 8326 5882 0 net23
rlabel metal1 8468 7514 8468 7514 0 net24
rlabel metal1 8652 4250 8652 4250 0 net25
rlabel metal1 5099 3026 5099 3026 0 net26
rlabel metal1 8372 10030 8372 10030 0 net27
rlabel metal1 6946 11084 6946 11084 0 net28
rlabel via1 8974 12614 8974 12614 0 net29
rlabel metal2 2852 8908 2852 8908 0 net3
rlabel viali 7134 12274 7134 12274 0 net30
rlabel metal1 5756 12614 5756 12614 0 net31
rlabel metal3 6164 11628 6164 11628 0 net32
rlabel metal1 1794 7752 1794 7752 0 net33
rlabel metal2 6394 5508 6394 5508 0 net34
rlabel metal1 4738 2006 4738 2006 0 net35
rlabel metal1 8698 11866 8698 11866 0 net36
rlabel metal2 966 12342 966 12342 0 net37
rlabel metal2 2254 5780 2254 5780 0 net38
rlabel metal1 5113 3434 5113 3434 0 net39
rlabel metal1 8832 11050 8832 11050 0 net4
rlabel metal2 6210 5882 6210 5882 0 net40
rlabel metal1 5290 13328 5290 13328 0 net41
rlabel metal1 1557 12138 1557 12138 0 net42
rlabel metal2 2346 6290 2346 6290 0 net43
rlabel metal3 8426 8228 8426 8228 0 net44
rlabel metal1 2392 13226 2392 13226 0 net45
rlabel metal1 7498 12410 7498 12410 0 net46
rlabel metal1 2116 13158 2116 13158 0 net47
rlabel metal2 2162 11169 2162 11169 0 net48
rlabel via1 4186 13957 4186 13957 0 net49
rlabel viali 7773 8942 7773 8942 0 net5
rlabel metal1 3450 9588 3450 9588 0 net50
rlabel metal1 1656 13158 1656 13158 0 net51
rlabel metal1 3956 8942 3956 8942 0 net52
rlabel viali 3174 9555 3174 9555 0 net53
rlabel viali 3726 9555 3726 9555 0 net54
rlabel metal2 4002 13702 4002 13702 0 net55
rlabel metal1 2851 9538 2851 9538 0 net56
rlabel metal1 5244 2006 5244 2006 0 net57
rlabel metal1 2990 12614 2990 12614 0 net58
rlabel metal1 2392 10234 2392 10234 0 net59
rlabel metal1 6026 11594 6026 11594 0 net6
rlabel metal2 4278 10030 4278 10030 0 net60
rlabel metal2 7222 3298 7222 3298 0 net61
rlabel metal2 4922 7276 4922 7276 0 net62
rlabel metal1 6072 10098 6072 10098 0 net63
rlabel metal1 6440 7310 6440 7310 0 net64
rlabel metal1 4002 11186 4002 11186 0 net65
rlabel metal1 6210 3944 6210 3944 0 net66
rlabel metal2 6854 12036 6854 12036 0 net67
rlabel metal2 5474 3026 5474 3026 0 net68
rlabel metal1 5152 11526 5152 11526 0 net69
rlabel metal1 6256 11730 6256 11730 0 net7
rlabel metal2 1702 8976 1702 8976 0 net70
rlabel metal1 6348 8874 6348 8874 0 net71
rlabel metal1 6440 11662 6440 11662 0 net72
rlabel metal1 3588 13226 3588 13226 0 net8
rlabel viali 6209 12818 6209 12818 0 net9
rlabel metal3 9024 3332 9024 3332 0 pad_gpio_ana_en
rlabel metal1 8740 5746 8740 5746 0 pad_gpio_ana_pol
rlabel metal3 9024 7412 9024 7412 0 pad_gpio_ana_sel
rlabel metal3 8932 4148 8932 4148 0 pad_gpio_dm[0]
rlabel metal2 5658 2737 5658 2737 0 pad_gpio_dm[1]
rlabel via2 9622 9860 9622 9860 0 pad_gpio_dm[2]
rlabel metal3 8886 10676 8886 10676 0 pad_gpio_holdover
rlabel metal1 9108 8398 9108 8398 0 pad_gpio_hys_trim
rlabel via2 9622 13124 9622 13124 0 pad_gpio_ib_mode_sel
rlabel metal2 9062 1105 9062 1105 0 pad_gpio_in
rlabel metal3 9254 6596 9254 6596 0 pad_gpio_inenb
rlabel metal3 9392 11492 9392 11492 0 pad_gpio_out
rlabel via2 9622 13940 9622 13940 0 pad_gpio_outenb
rlabel via2 9622 4964 9622 4964 0 pad_gpio_slew_ctl[0]
rlabel via2 9622 1700 9622 1700 0 pad_gpio_slow_sel
rlabel metal3 9070 12308 9070 12308 0 pad_gpio_vtrip_sel
rlabel metal3 1196 2516 1196 2516 0 resetn
rlabel metal3 406 10132 406 10132 0 resetn_out
rlabel metal2 966 3961 966 3961 0 serial_clock
rlabel metal3 682 10948 682 10948 0 serial_clock_out
rlabel metal3 406 4420 406 4420 0 serial_data_in
rlabel metal3 866 12580 866 12580 0 serial_data_out
rlabel metal1 1150 8466 1150 8466 0 serial_load
rlabel metal3 360 11764 360 11764 0 serial_load_out
rlabel metal1 2576 5134 2576 5134 0 shift_register\[0\]
rlabel metal1 4278 4692 4278 4692 0 shift_register\[10\]
rlabel metal1 7498 1802 7498 1802 0 shift_register\[11\]
rlabel metal1 7774 6766 7774 6766 0 shift_register\[12\]
rlabel metal1 5474 9146 5474 9146 0 shift_register\[13\]
rlabel metal1 3312 10166 3312 10166 0 shift_register\[14\]
rlabel metal2 2438 11764 2438 11764 0 shift_register\[15\]
rlabel metal1 2346 9486 2346 9486 0 shift_register\[1\]
rlabel metal1 3933 10506 3933 10506 0 shift_register\[2\]
rlabel metal1 2024 12750 2024 12750 0 shift_register\[3\]
rlabel metal1 4692 11662 4692 11662 0 shift_register\[4\]
rlabel metal2 3266 7684 3266 7684 0 shift_register\[5\]
rlabel metal1 5888 6426 5888 6426 0 shift_register\[6\]
rlabel metal1 6716 5882 6716 5882 0 shift_register\[7\]
rlabel metal1 5428 2414 5428 2414 0 shift_register\[8\]
rlabel metal1 4554 3706 4554 3706 0 shift_register\[9\]
rlabel metal3 360 9316 360 9316 0 user_gpio_in
rlabel metal1 3174 8908 3174 8908 0 user_gpio_oeb
rlabel metal3 636 7684 636 7684 0 user_gpio_out
<< properties >>
string FIXED_BBOX 0 0 10000 14800
<< end >>
