VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO mgmt_protect
  CLASS BLOCK ;
  FOREIGN mgmt_protect ;
  ORIGIN 0.000 0.000 ;
  SIZE 220.000 BY 60.000 ;
  PIN frigate_HCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 15.270 0.000 15.550 2.000 ;
    END
  END frigate_HCLK
  PIN frigate_HRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 2.000 ;
    END
  END frigate_HRESETn
  PIN mprj_AHB_Ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 161.550 0.000 161.830 2.000 ;
    END
  END mprj_AHB_Ena
  PIN mprj_HADDR_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 24.930 0.000 25.210 2.000 ;
    END
  END mprj_HADDR_core[0]
  PIN mprj_HADDR_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 2.000 ;
    END
  END mprj_HADDR_core[10]
  PIN mprj_HADDR_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 40.110 0.000 40.390 2.000 ;
    END
  END mprj_HADDR_core[11]
  PIN mprj_HADDR_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 2.000 ;
    END
  END mprj_HADDR_core[12]
  PIN mprj_HADDR_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 42.870 0.000 43.150 2.000 ;
    END
  END mprj_HADDR_core[13]
  PIN mprj_HADDR_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 2.000 ;
    END
  END mprj_HADDR_core[14]
  PIN mprj_HADDR_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.630 0.000 45.910 2.000 ;
    END
  END mprj_HADDR_core[15]
  PIN mprj_HADDR_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 2.000 ;
    END
  END mprj_HADDR_core[16]
  PIN mprj_HADDR_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 2.000 ;
    END
  END mprj_HADDR_core[17]
  PIN mprj_HADDR_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 0.000 50.050 2.000 ;
    END
  END mprj_HADDR_core[18]
  PIN mprj_HADDR_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.150 0.000 51.430 2.000 ;
    END
  END mprj_HADDR_core[19]
  PIN mprj_HADDR_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 2.000 ;
    END
  END mprj_HADDR_core[1]
  PIN mprj_HADDR_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 52.530 0.000 52.810 2.000 ;
    END
  END mprj_HADDR_core[20]
  PIN mprj_HADDR_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 53.910 0.000 54.190 2.000 ;
    END
  END mprj_HADDR_core[21]
  PIN mprj_HADDR_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 2.000 ;
    END
  END mprj_HADDR_core[22]
  PIN mprj_HADDR_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 56.670 0.000 56.950 2.000 ;
    END
  END mprj_HADDR_core[23]
  PIN mprj_HADDR_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 2.000 ;
    END
  END mprj_HADDR_core[24]
  PIN mprj_HADDR_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 2.000 ;
    END
  END mprj_HADDR_core[25]
  PIN mprj_HADDR_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 60.810 0.000 61.090 2.000 ;
    END
  END mprj_HADDR_core[26]
  PIN mprj_HADDR_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 2.000 ;
    END
  END mprj_HADDR_core[27]
  PIN mprj_HADDR_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 63.570 0.000 63.850 2.000 ;
    END
  END mprj_HADDR_core[28]
  PIN mprj_HADDR_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 64.950 0.000 65.230 2.000 ;
    END
  END mprj_HADDR_core[29]
  PIN mprj_HADDR_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 2.000 ;
    END
  END mprj_HADDR_core[2]
  PIN mprj_HADDR_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 2.000 ;
    END
  END mprj_HADDR_core[30]
  PIN mprj_HADDR_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 2.000 ;
    END
  END mprj_HADDR_core[31]
  PIN mprj_HADDR_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 2.000 ;
    END
  END mprj_HADDR_core[3]
  PIN mprj_HADDR_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 2.000 ;
    END
  END mprj_HADDR_core[4]
  PIN mprj_HADDR_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 2.000 ;
    END
  END mprj_HADDR_core[5]
  PIN mprj_HADDR_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 33.210 0.000 33.490 2.000 ;
    END
  END mprj_HADDR_core[6]
  PIN mprj_HADDR_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 2.000 ;
    END
  END mprj_HADDR_core[7]
  PIN mprj_HADDR_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.970 0.000 36.250 2.000 ;
    END
  END mprj_HADDR_core[8]
  PIN mprj_HADDR_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 37.350 0.000 37.630 2.000 ;
    END
  END mprj_HADDR_core[9]
  PIN mprj_HADDR_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 36.430 58.000 36.710 60.000 ;
    END
  END mprj_HADDR_user[0]
  PIN mprj_HADDR_user[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 50.230 58.000 50.510 60.000 ;
    END
  END mprj_HADDR_user[10]
  PIN mprj_HADDR_user[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 58.000 51.890 60.000 ;
    END
  END mprj_HADDR_user[11]
  PIN mprj_HADDR_user[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 52.990 58.000 53.270 60.000 ;
    END
  END mprj_HADDR_user[12]
  PIN mprj_HADDR_user[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 54.370 58.000 54.650 60.000 ;
    END
  END mprj_HADDR_user[13]
  PIN mprj_HADDR_user[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 55.750 58.000 56.030 60.000 ;
    END
  END mprj_HADDR_user[14]
  PIN mprj_HADDR_user[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 57.130 58.000 57.410 60.000 ;
    END
  END mprj_HADDR_user[15]
  PIN mprj_HADDR_user[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 58.510 58.000 58.790 60.000 ;
    END
  END mprj_HADDR_user[16]
  PIN mprj_HADDR_user[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 59.890 58.000 60.170 60.000 ;
    END
  END mprj_HADDR_user[17]
  PIN mprj_HADDR_user[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 61.270 58.000 61.550 60.000 ;
    END
  END mprj_HADDR_user[18]
  PIN mprj_HADDR_user[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 62.650 58.000 62.930 60.000 ;
    END
  END mprj_HADDR_user[19]
  PIN mprj_HADDR_user[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 37.810 58.000 38.090 60.000 ;
    END
  END mprj_HADDR_user[1]
  PIN mprj_HADDR_user[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 64.030 58.000 64.310 60.000 ;
    END
  END mprj_HADDR_user[20]
  PIN mprj_HADDR_user[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 65.410 58.000 65.690 60.000 ;
    END
  END mprj_HADDR_user[21]
  PIN mprj_HADDR_user[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 66.790 58.000 67.070 60.000 ;
    END
  END mprj_HADDR_user[22]
  PIN mprj_HADDR_user[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 68.170 58.000 68.450 60.000 ;
    END
  END mprj_HADDR_user[23]
  PIN mprj_HADDR_user[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 69.550 58.000 69.830 60.000 ;
    END
  END mprj_HADDR_user[24]
  PIN mprj_HADDR_user[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 70.930 58.000 71.210 60.000 ;
    END
  END mprj_HADDR_user[25]
  PIN mprj_HADDR_user[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 72.310 58.000 72.590 60.000 ;
    END
  END mprj_HADDR_user[26]
  PIN mprj_HADDR_user[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 73.690 58.000 73.970 60.000 ;
    END
  END mprj_HADDR_user[27]
  PIN mprj_HADDR_user[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 75.070 58.000 75.350 60.000 ;
    END
  END mprj_HADDR_user[28]
  PIN mprj_HADDR_user[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 76.450 58.000 76.730 60.000 ;
    END
  END mprj_HADDR_user[29]
  PIN mprj_HADDR_user[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 39.190 58.000 39.470 60.000 ;
    END
  END mprj_HADDR_user[2]
  PIN mprj_HADDR_user[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 77.830 58.000 78.110 60.000 ;
    END
  END mprj_HADDR_user[30]
  PIN mprj_HADDR_user[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 79.210 58.000 79.490 60.000 ;
    END
  END mprj_HADDR_user[31]
  PIN mprj_HADDR_user[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 40.570 58.000 40.850 60.000 ;
    END
  END mprj_HADDR_user[3]
  PIN mprj_HADDR_user[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 41.950 58.000 42.230 60.000 ;
    END
  END mprj_HADDR_user[4]
  PIN mprj_HADDR_user[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 43.330 58.000 43.610 60.000 ;
    END
  END mprj_HADDR_user[5]
  PIN mprj_HADDR_user[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 44.710 58.000 44.990 60.000 ;
    END
  END mprj_HADDR_user[6]
  PIN mprj_HADDR_user[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 46.090 58.000 46.370 60.000 ;
    END
  END mprj_HADDR_user[7]
  PIN mprj_HADDR_user[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 47.470 58.000 47.750 60.000 ;
    END
  END mprj_HADDR_user[8]
  PIN mprj_HADDR_user[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 48.850 58.000 49.130 60.000 ;
    END
  END mprj_HADDR_user[9]
  PIN mprj_HRDATA_core[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 2.000 ;
    END
  END mprj_HRDATA_core[0]
  PIN mprj_HRDATA_core[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 2.000 ;
    END
  END mprj_HRDATA_core[10]
  PIN mprj_HRDATA_core[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 2.000 ;
    END
  END mprj_HRDATA_core[11]
  PIN mprj_HRDATA_core[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 2.000 ;
    END
  END mprj_HRDATA_core[12]
  PIN mprj_HRDATA_core[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 133.950 0.000 134.230 2.000 ;
    END
  END mprj_HRDATA_core[13]
  PIN mprj_HRDATA_core[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 2.000 ;
    END
  END mprj_HRDATA_core[14]
  PIN mprj_HRDATA_core[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 136.710 0.000 136.990 2.000 ;
    END
  END mprj_HRDATA_core[15]
  PIN mprj_HRDATA_core[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 138.090 0.000 138.370 2.000 ;
    END
  END mprj_HRDATA_core[16]
  PIN mprj_HRDATA_core[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 139.470 0.000 139.750 2.000 ;
    END
  END mprj_HRDATA_core[17]
  PIN mprj_HRDATA_core[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 2.000 ;
    END
  END mprj_HRDATA_core[18]
  PIN mprj_HRDATA_core[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 2.000 ;
    END
  END mprj_HRDATA_core[19]
  PIN mprj_HRDATA_core[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 2.000 ;
    END
  END mprj_HRDATA_core[1]
  PIN mprj_HRDATA_core[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 2.000 ;
    END
  END mprj_HRDATA_core[20]
  PIN mprj_HRDATA_core[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 2.000 ;
    END
  END mprj_HRDATA_core[21]
  PIN mprj_HRDATA_core[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 146.370 0.000 146.650 2.000 ;
    END
  END mprj_HRDATA_core[22]
  PIN mprj_HRDATA_core[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 147.750 0.000 148.030 2.000 ;
    END
  END mprj_HRDATA_core[23]
  PIN mprj_HRDATA_core[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 149.130 0.000 149.410 2.000 ;
    END
  END mprj_HRDATA_core[24]
  PIN mprj_HRDATA_core[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 2.000 ;
    END
  END mprj_HRDATA_core[25]
  PIN mprj_HRDATA_core[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 151.890 0.000 152.170 2.000 ;
    END
  END mprj_HRDATA_core[26]
  PIN mprj_HRDATA_core[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 153.270 0.000 153.550 2.000 ;
    END
  END mprj_HRDATA_core[27]
  PIN mprj_HRDATA_core[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 2.000 ;
    END
  END mprj_HRDATA_core[28]
  PIN mprj_HRDATA_core[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 156.030 0.000 156.310 2.000 ;
    END
  END mprj_HRDATA_core[29]
  PIN mprj_HRDATA_core[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 118.770 0.000 119.050 2.000 ;
    END
  END mprj_HRDATA_core[2]
  PIN mprj_HRDATA_core[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 2.000 ;
    END
  END mprj_HRDATA_core[30]
  PIN mprj_HRDATA_core[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 158.790 0.000 159.070 2.000 ;
    END
  END mprj_HRDATA_core[31]
  PIN mprj_HRDATA_core[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 120.150 0.000 120.430 2.000 ;
    END
  END mprj_HRDATA_core[3]
  PIN mprj_HRDATA_core[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 2.000 ;
    END
  END mprj_HRDATA_core[4]
  PIN mprj_HRDATA_core[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 2.000 ;
    END
  END mprj_HRDATA_core[5]
  PIN mprj_HRDATA_core[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 2.000 ;
    END
  END mprj_HRDATA_core[6]
  PIN mprj_HRDATA_core[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 2.000 ;
    END
  END mprj_HRDATA_core[7]
  PIN mprj_HRDATA_core[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 127.050 0.000 127.330 2.000 ;
    END
  END mprj_HRDATA_core[8]
  PIN mprj_HRDATA_core[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 128.430 0.000 128.710 2.000 ;
    END
  END mprj_HRDATA_core[9]
  PIN mprj_HRDATA_user[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 127.510 58.000 127.790 60.000 ;
    END
  END mprj_HRDATA_user[0]
  PIN mprj_HRDATA_user[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 141.310 58.000 141.590 60.000 ;
    END
  END mprj_HRDATA_user[10]
  PIN mprj_HRDATA_user[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 142.690 58.000 142.970 60.000 ;
    END
  END mprj_HRDATA_user[11]
  PIN mprj_HRDATA_user[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 144.070 58.000 144.350 60.000 ;
    END
  END mprj_HRDATA_user[12]
  PIN mprj_HRDATA_user[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 145.450 58.000 145.730 60.000 ;
    END
  END mprj_HRDATA_user[13]
  PIN mprj_HRDATA_user[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 146.830 58.000 147.110 60.000 ;
    END
  END mprj_HRDATA_user[14]
  PIN mprj_HRDATA_user[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 148.210 58.000 148.490 60.000 ;
    END
  END mprj_HRDATA_user[15]
  PIN mprj_HRDATA_user[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 149.590 58.000 149.870 60.000 ;
    END
  END mprj_HRDATA_user[16]
  PIN mprj_HRDATA_user[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 150.970 58.000 151.250 60.000 ;
    END
  END mprj_HRDATA_user[17]
  PIN mprj_HRDATA_user[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 152.350 58.000 152.630 60.000 ;
    END
  END mprj_HRDATA_user[18]
  PIN mprj_HRDATA_user[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 153.730 58.000 154.010 60.000 ;
    END
  END mprj_HRDATA_user[19]
  PIN mprj_HRDATA_user[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 128.890 58.000 129.170 60.000 ;
    END
  END mprj_HRDATA_user[1]
  PIN mprj_HRDATA_user[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 155.110 58.000 155.390 60.000 ;
    END
  END mprj_HRDATA_user[20]
  PIN mprj_HRDATA_user[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 156.490 58.000 156.770 60.000 ;
    END
  END mprj_HRDATA_user[21]
  PIN mprj_HRDATA_user[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 157.870 58.000 158.150 60.000 ;
    END
  END mprj_HRDATA_user[22]
  PIN mprj_HRDATA_user[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 159.250 58.000 159.530 60.000 ;
    END
  END mprj_HRDATA_user[23]
  PIN mprj_HRDATA_user[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 160.630 58.000 160.910 60.000 ;
    END
  END mprj_HRDATA_user[24]
  PIN mprj_HRDATA_user[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.010 58.000 162.290 60.000 ;
    END
  END mprj_HRDATA_user[25]
  PIN mprj_HRDATA_user[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 163.390 58.000 163.670 60.000 ;
    END
  END mprj_HRDATA_user[26]
  PIN mprj_HRDATA_user[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 164.770 58.000 165.050 60.000 ;
    END
  END mprj_HRDATA_user[27]
  PIN mprj_HRDATA_user[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 166.150 58.000 166.430 60.000 ;
    END
  END mprj_HRDATA_user[28]
  PIN mprj_HRDATA_user[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 167.530 58.000 167.810 60.000 ;
    END
  END mprj_HRDATA_user[29]
  PIN mprj_HRDATA_user[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 130.270 58.000 130.550 60.000 ;
    END
  END mprj_HRDATA_user[2]
  PIN mprj_HRDATA_user[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 168.910 58.000 169.190 60.000 ;
    END
  END mprj_HRDATA_user[30]
  PIN mprj_HRDATA_user[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 170.290 58.000 170.570 60.000 ;
    END
  END mprj_HRDATA_user[31]
  PIN mprj_HRDATA_user[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 131.650 58.000 131.930 60.000 ;
    END
  END mprj_HRDATA_user[3]
  PIN mprj_HRDATA_user[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 133.030 58.000 133.310 60.000 ;
    END
  END mprj_HRDATA_user[4]
  PIN mprj_HRDATA_user[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 134.410 58.000 134.690 60.000 ;
    END
  END mprj_HRDATA_user[5]
  PIN mprj_HRDATA_user[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 135.790 58.000 136.070 60.000 ;
    END
  END mprj_HRDATA_user[6]
  PIN mprj_HRDATA_user[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 137.170 58.000 137.450 60.000 ;
    END
  END mprj_HRDATA_user[7]
  PIN mprj_HRDATA_user[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 138.550 58.000 138.830 60.000 ;
    END
  END mprj_HRDATA_user[8]
  PIN mprj_HRDATA_user[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 139.930 58.000 140.210 60.000 ;
    END
  END mprj_HRDATA_user[9]
  PIN mprj_HREADYOUT_core
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 2.000 ;
    END
  END mprj_HREADYOUT_core
  PIN mprj_HREADYOUT_user
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 171.670 58.000 171.950 60.000 ;
    END
  END mprj_HREADYOUT_user
  PIN mprj_HREADY_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 18.030 0.000 18.310 2.000 ;
    END
  END mprj_HREADY_core
  PIN mprj_HREADY_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 29.530 58.000 29.810 60.000 ;
    END
  END mprj_HREADY_user
  PIN mprj_HSEL_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 2.000 ;
    END
  END mprj_HSEL_core
  PIN mprj_HSEL_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 28.150 58.000 28.430 60.000 ;
    END
  END mprj_HSEL_user
  PIN mprj_HSIZE_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.790 0.000 21.070 2.000 ;
    END
  END mprj_HSIZE_core[0]
  PIN mprj_HSIZE_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 22.170 0.000 22.450 2.000 ;
    END
  END mprj_HSIZE_core[1]
  PIN mprj_HSIZE_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 23.550 0.000 23.830 2.000 ;
    END
  END mprj_HSIZE_core[2]
  PIN mprj_HSIZE_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 58.000 32.570 60.000 ;
    END
  END mprj_HSIZE_user[0]
  PIN mprj_HSIZE_user[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 33.670 58.000 33.950 60.000 ;
    END
  END mprj_HSIZE_user[1]
  PIN mprj_HSIZE_user[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 35.050 58.000 35.330 60.000 ;
    END
  END mprj_HSIZE_user[2]
  PIN mprj_HTRANS_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 113.250 0.000 113.530 2.000 ;
    END
  END mprj_HTRANS_core[0]
  PIN mprj_HTRANS_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 2.000 ;
    END
  END mprj_HTRANS_core[1]
  PIN mprj_HTRANS_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 124.750 58.000 125.030 60.000 ;
    END
  END mprj_HTRANS_user[0]
  PIN mprj_HTRANS_user[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 126.130 58.000 126.410 60.000 ;
    END
  END mprj_HTRANS_user[1]
  PIN mprj_HWDATA_core[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 2.000 ;
    END
  END mprj_HWDATA_core[0]
  PIN mprj_HWDATA_core[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 82.890 0.000 83.170 2.000 ;
    END
  END mprj_HWDATA_core[10]
  PIN mprj_HWDATA_core[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.270 0.000 84.550 2.000 ;
    END
  END mprj_HWDATA_core[11]
  PIN mprj_HWDATA_core[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 85.650 0.000 85.930 2.000 ;
    END
  END mprj_HWDATA_core[12]
  PIN mprj_HWDATA_core[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 2.000 ;
    END
  END mprj_HWDATA_core[13]
  PIN mprj_HWDATA_core[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 2.000 ;
    END
  END mprj_HWDATA_core[14]
  PIN mprj_HWDATA_core[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 2.000 ;
    END
  END mprj_HWDATA_core[15]
  PIN mprj_HWDATA_core[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 2.000 ;
    END
  END mprj_HWDATA_core[16]
  PIN mprj_HWDATA_core[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 92.550 0.000 92.830 2.000 ;
    END
  END mprj_HWDATA_core[17]
  PIN mprj_HWDATA_core[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 93.930 0.000 94.210 2.000 ;
    END
  END mprj_HWDATA_core[18]
  PIN mprj_HWDATA_core[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 95.310 0.000 95.590 2.000 ;
    END
  END mprj_HWDATA_core[19]
  PIN mprj_HWDATA_core[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.470 0.000 70.750 2.000 ;
    END
  END mprj_HWDATA_core[1]
  PIN mprj_HWDATA_core[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 2.000 ;
    END
  END mprj_HWDATA_core[20]
  PIN mprj_HWDATA_core[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 2.000 ;
    END
  END mprj_HWDATA_core[21]
  PIN mprj_HWDATA_core[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 2.000 ;
    END
  END mprj_HWDATA_core[22]
  PIN mprj_HWDATA_core[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 100.830 0.000 101.110 2.000 ;
    END
  END mprj_HWDATA_core[23]
  PIN mprj_HWDATA_core[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 2.000 ;
    END
  END mprj_HWDATA_core[24]
  PIN mprj_HWDATA_core[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 2.000 ;
    END
  END mprj_HWDATA_core[25]
  PIN mprj_HWDATA_core[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 104.970 0.000 105.250 2.000 ;
    END
  END mprj_HWDATA_core[26]
  PIN mprj_HWDATA_core[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 2.000 ;
    END
  END mprj_HWDATA_core[27]
  PIN mprj_HWDATA_core[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 107.730 0.000 108.010 2.000 ;
    END
  END mprj_HWDATA_core[28]
  PIN mprj_HWDATA_core[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.110 0.000 109.390 2.000 ;
    END
  END mprj_HWDATA_core[29]
  PIN mprj_HWDATA_core[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 2.000 ;
    END
  END mprj_HWDATA_core[2]
  PIN mprj_HWDATA_core[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 2.000 ;
    END
  END mprj_HWDATA_core[30]
  PIN mprj_HWDATA_core[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 111.870 0.000 112.150 2.000 ;
    END
  END mprj_HWDATA_core[31]
  PIN mprj_HWDATA_core[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 73.230 0.000 73.510 2.000 ;
    END
  END mprj_HWDATA_core[3]
  PIN mprj_HWDATA_core[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 2.000 ;
    END
  END mprj_HWDATA_core[4]
  PIN mprj_HWDATA_core[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 2.000 ;
    END
  END mprj_HWDATA_core[5]
  PIN mprj_HWDATA_core[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 2.000 ;
    END
  END mprj_HWDATA_core[6]
  PIN mprj_HWDATA_core[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 2.000 ;
    END
  END mprj_HWDATA_core[7]
  PIN mprj_HWDATA_core[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 80.130 0.000 80.410 2.000 ;
    END
  END mprj_HWDATA_core[8]
  PIN mprj_HWDATA_core[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.510 0.000 81.790 2.000 ;
    END
  END mprj_HWDATA_core[9]
  PIN mprj_HWDATA_user[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 80.590 58.000 80.870 60.000 ;
    END
  END mprj_HWDATA_user[0]
  PIN mprj_HWDATA_user[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 94.390 58.000 94.670 60.000 ;
    END
  END mprj_HWDATA_user[10]
  PIN mprj_HWDATA_user[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 95.770 58.000 96.050 60.000 ;
    END
  END mprj_HWDATA_user[11]
  PIN mprj_HWDATA_user[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 97.150 58.000 97.430 60.000 ;
    END
  END mprj_HWDATA_user[12]
  PIN mprj_HWDATA_user[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 98.530 58.000 98.810 60.000 ;
    END
  END mprj_HWDATA_user[13]
  PIN mprj_HWDATA_user[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 99.910 58.000 100.190 60.000 ;
    END
  END mprj_HWDATA_user[14]
  PIN mprj_HWDATA_user[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 101.290 58.000 101.570 60.000 ;
    END
  END mprj_HWDATA_user[15]
  PIN mprj_HWDATA_user[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 102.670 58.000 102.950 60.000 ;
    END
  END mprj_HWDATA_user[16]
  PIN mprj_HWDATA_user[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 104.050 58.000 104.330 60.000 ;
    END
  END mprj_HWDATA_user[17]
  PIN mprj_HWDATA_user[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 105.430 58.000 105.710 60.000 ;
    END
  END mprj_HWDATA_user[18]
  PIN mprj_HWDATA_user[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 106.810 58.000 107.090 60.000 ;
    END
  END mprj_HWDATA_user[19]
  PIN mprj_HWDATA_user[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 81.970 58.000 82.250 60.000 ;
    END
  END mprj_HWDATA_user[1]
  PIN mprj_HWDATA_user[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 108.190 58.000 108.470 60.000 ;
    END
  END mprj_HWDATA_user[20]
  PIN mprj_HWDATA_user[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 109.570 58.000 109.850 60.000 ;
    END
  END mprj_HWDATA_user[21]
  PIN mprj_HWDATA_user[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 110.950 58.000 111.230 60.000 ;
    END
  END mprj_HWDATA_user[22]
  PIN mprj_HWDATA_user[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 112.330 58.000 112.610 60.000 ;
    END
  END mprj_HWDATA_user[23]
  PIN mprj_HWDATA_user[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 113.710 58.000 113.990 60.000 ;
    END
  END mprj_HWDATA_user[24]
  PIN mprj_HWDATA_user[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 115.090 58.000 115.370 60.000 ;
    END
  END mprj_HWDATA_user[25]
  PIN mprj_HWDATA_user[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 116.470 58.000 116.750 60.000 ;
    END
  END mprj_HWDATA_user[26]
  PIN mprj_HWDATA_user[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 117.850 58.000 118.130 60.000 ;
    END
  END mprj_HWDATA_user[27]
  PIN mprj_HWDATA_user[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 119.230 58.000 119.510 60.000 ;
    END
  END mprj_HWDATA_user[28]
  PIN mprj_HWDATA_user[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 120.610 58.000 120.890 60.000 ;
    END
  END mprj_HWDATA_user[29]
  PIN mprj_HWDATA_user[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 83.350 58.000 83.630 60.000 ;
    END
  END mprj_HWDATA_user[2]
  PIN mprj_HWDATA_user[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 121.990 58.000 122.270 60.000 ;
    END
  END mprj_HWDATA_user[30]
  PIN mprj_HWDATA_user[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 123.370 58.000 123.650 60.000 ;
    END
  END mprj_HWDATA_user[31]
  PIN mprj_HWDATA_user[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 84.730 58.000 85.010 60.000 ;
    END
  END mprj_HWDATA_user[3]
  PIN mprj_HWDATA_user[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 86.110 58.000 86.390 60.000 ;
    END
  END mprj_HWDATA_user[4]
  PIN mprj_HWDATA_user[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 87.490 58.000 87.770 60.000 ;
    END
  END mprj_HWDATA_user[5]
  PIN mprj_HWDATA_user[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 88.870 58.000 89.150 60.000 ;
    END
  END mprj_HWDATA_user[6]
  PIN mprj_HWDATA_user[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 58.000 90.530 60.000 ;
    END
  END mprj_HWDATA_user[7]
  PIN mprj_HWDATA_user[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 91.630 58.000 91.910 60.000 ;
    END
  END mprj_HWDATA_user[8]
  PIN mprj_HWDATA_user[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 93.010 58.000 93.290 60.000 ;
    END
  END mprj_HWDATA_user[9]
  PIN mprj_HWRITE_core
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 2.000 ;
    END
  END mprj_HWRITE_core
  PIN mprj_HWRITE_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 30.910 58.000 31.190 60.000 ;
    END
  END mprj_HWRITE_user
  PIN user_HCLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 25.390 58.000 25.670 60.000 ;
    END
  END user_HCLK
  PIN user_HRESETn
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 1.358700 ;
    PORT
      LAYER met2 ;
        RECT 26.770 58.000 27.050 60.000 ;
    END
  END user_HRESETn
  PIN user_irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.050 58.000 173.330 60.000 ;
    END
  END user_irq[0]
  PIN user_irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 186.850 58.000 187.130 60.000 ;
    END
  END user_irq[10]
  PIN user_irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 188.230 58.000 188.510 60.000 ;
    END
  END user_irq[11]
  PIN user_irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 189.610 58.000 189.890 60.000 ;
    END
  END user_irq[12]
  PIN user_irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 190.990 58.000 191.270 60.000 ;
    END
  END user_irq[13]
  PIN user_irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 192.370 58.000 192.650 60.000 ;
    END
  END user_irq[14]
  PIN user_irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 193.750 58.000 194.030 60.000 ;
    END
  END user_irq[15]
  PIN user_irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 174.430 58.000 174.710 60.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 175.810 58.000 176.090 60.000 ;
    END
  END user_irq[2]
  PIN user_irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 177.190 58.000 177.470 60.000 ;
    END
  END user_irq[3]
  PIN user_irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 178.570 58.000 178.850 60.000 ;
    END
  END user_irq[4]
  PIN user_irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 179.950 58.000 180.230 60.000 ;
    END
  END user_irq[5]
  PIN user_irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 181.330 58.000 181.610 60.000 ;
    END
  END user_irq[6]
  PIN user_irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 182.710 58.000 182.990 60.000 ;
    END
  END user_irq[7]
  PIN user_irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 184.090 58.000 184.370 60.000 ;
    END
  END user_irq[8]
  PIN user_irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 185.470 58.000 185.750 60.000 ;
    END
  END user_irq[9]
  PIN user_irq_core[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 2.000 ;
    END
  END user_irq_core[0]
  PIN user_irq_core[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 2.000 ;
    END
  END user_irq_core[10]
  PIN user_irq_core[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 2.000 ;
    END
  END user_irq_core[11]
  PIN user_irq_core[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 2.000 ;
    END
  END user_irq_core[12]
  PIN user_irq_core[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 2.000 ;
    END
  END user_irq_core[13]
  PIN user_irq_core[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 2.000 ;
    END
  END user_irq_core[14]
  PIN user_irq_core[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 205.710 0.000 205.990 2.000 ;
    END
  END user_irq_core[15]
  PIN user_irq_core[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 186.390 0.000 186.670 2.000 ;
    END
  END user_irq_core[1]
  PIN user_irq_core[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 2.000 ;
    END
  END user_irq_core[2]
  PIN user_irq_core[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 189.150 0.000 189.430 2.000 ;
    END
  END user_irq_core[3]
  PIN user_irq_core[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 190.530 0.000 190.810 2.000 ;
    END
  END user_irq_core[4]
  PIN user_irq_core[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 191.910 0.000 192.190 2.000 ;
    END
  END user_irq_core[5]
  PIN user_irq_core[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 193.290 0.000 193.570 2.000 ;
    END
  END user_irq_core[6]
  PIN user_irq_core[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 194.670 0.000 194.950 2.000 ;
    END
  END user_irq_core[7]
  PIN user_irq_core[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 196.050 0.000 196.330 2.000 ;
    END
  END user_irq_core[8]
  PIN user_irq_core[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.880200 ;
    PORT
      LAYER met2 ;
        RECT 197.430 0.000 197.710 2.000 ;
    END
  END user_irq_core[9]
  PIN user_irq_ena[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.930 0.000 163.210 2.000 ;
    END
  END user_irq_ena[0]
  PIN user_irq_ena[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 2.000 ;
    END
  END user_irq_ena[10]
  PIN user_irq_ena[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 178.110 0.000 178.390 2.000 ;
    END
  END user_irq_ena[11]
  PIN user_irq_ena[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 179.490 0.000 179.770 2.000 ;
    END
  END user_irq_ena[12]
  PIN user_irq_ena[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.870 0.000 181.150 2.000 ;
    END
  END user_irq_ena[13]
  PIN user_irq_ena[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 182.250 0.000 182.530 2.000 ;
    END
  END user_irq_ena[14]
  PIN user_irq_ena[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 2.000 ;
    END
  END user_irq_ena[15]
  PIN user_irq_ena[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 2.000 ;
    END
  END user_irq_ena[1]
  PIN user_irq_ena[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 2.000 ;
    END
  END user_irq_ena[2]
  PIN user_irq_ena[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 167.070 0.000 167.350 2.000 ;
    END
  END user_irq_ena[3]
  PIN user_irq_ena[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 168.450 0.000 168.730 2.000 ;
    END
  END user_irq_ena[4]
  PIN user_irq_ena[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 2.000 ;
    END
  END user_irq_ena[5]
  PIN user_irq_ena[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 171.210 0.000 171.490 2.000 ;
    END
  END user_irq_ena[6]
  PIN user_irq_ena[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 2.000 ;
    END
  END user_irq_ena[7]
  PIN user_irq_ena[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 2.000 ;
    END
  END user_irq_ena[8]
  PIN user_irq_ena[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 175.350 0.000 175.630 2.000 ;
    END
  END user_irq_ena[9]
  PIN vccd0
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 6.500 2.480 8.100 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 46.500 2.480 48.100 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 86.500 2.480 88.100 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.500 2.480 128.100 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.500 2.480 168.100 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 206.500 2.480 208.100 57.360 ;
    END
  END vccd0
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 92.900 2.480 94.500 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 132.900 2.480 134.500 57.360 ;
    END
  END vccd1
  PIN vssd0
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 9.700 2.480 11.300 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 49.700 2.480 51.300 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 89.700 2.480 91.300 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.700 2.480 131.300 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 169.700 2.480 171.300 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 209.700 2.480 211.300 57.360 ;
    END
  END vssd0
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 96.100 2.480 97.700 57.360 ;
    END
    PORT
      LAYER met4 ;
        RECT 136.100 2.480 137.700 57.360 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 2.110 2.635 217.770 57.205 ;
      LAYER li1 ;
        RECT 2.300 2.635 217.580 57.205 ;
      LAYER met1 ;
        RECT 2.300 0.040 217.580 58.100 ;
      LAYER met2 ;
        RECT 6.530 57.720 25.110 58.130 ;
        RECT 25.950 57.720 26.490 58.130 ;
        RECT 27.330 57.720 27.870 58.130 ;
        RECT 28.710 57.720 29.250 58.130 ;
        RECT 30.090 57.720 30.630 58.130 ;
        RECT 31.470 57.720 32.010 58.130 ;
        RECT 32.850 57.720 33.390 58.130 ;
        RECT 34.230 57.720 34.770 58.130 ;
        RECT 35.610 57.720 36.150 58.130 ;
        RECT 36.990 57.720 37.530 58.130 ;
        RECT 38.370 57.720 38.910 58.130 ;
        RECT 39.750 57.720 40.290 58.130 ;
        RECT 41.130 57.720 41.670 58.130 ;
        RECT 42.510 57.720 43.050 58.130 ;
        RECT 43.890 57.720 44.430 58.130 ;
        RECT 45.270 57.720 45.810 58.130 ;
        RECT 46.650 57.720 47.190 58.130 ;
        RECT 48.030 57.720 48.570 58.130 ;
        RECT 49.410 57.720 49.950 58.130 ;
        RECT 50.790 57.720 51.330 58.130 ;
        RECT 52.170 57.720 52.710 58.130 ;
        RECT 53.550 57.720 54.090 58.130 ;
        RECT 54.930 57.720 55.470 58.130 ;
        RECT 56.310 57.720 56.850 58.130 ;
        RECT 57.690 57.720 58.230 58.130 ;
        RECT 59.070 57.720 59.610 58.130 ;
        RECT 60.450 57.720 60.990 58.130 ;
        RECT 61.830 57.720 62.370 58.130 ;
        RECT 63.210 57.720 63.750 58.130 ;
        RECT 64.590 57.720 65.130 58.130 ;
        RECT 65.970 57.720 66.510 58.130 ;
        RECT 67.350 57.720 67.890 58.130 ;
        RECT 68.730 57.720 69.270 58.130 ;
        RECT 70.110 57.720 70.650 58.130 ;
        RECT 71.490 57.720 72.030 58.130 ;
        RECT 72.870 57.720 73.410 58.130 ;
        RECT 74.250 57.720 74.790 58.130 ;
        RECT 75.630 57.720 76.170 58.130 ;
        RECT 77.010 57.720 77.550 58.130 ;
        RECT 78.390 57.720 78.930 58.130 ;
        RECT 79.770 57.720 80.310 58.130 ;
        RECT 81.150 57.720 81.690 58.130 ;
        RECT 82.530 57.720 83.070 58.130 ;
        RECT 83.910 57.720 84.450 58.130 ;
        RECT 85.290 57.720 85.830 58.130 ;
        RECT 86.670 57.720 87.210 58.130 ;
        RECT 88.050 57.720 88.590 58.130 ;
        RECT 89.430 57.720 89.970 58.130 ;
        RECT 90.810 57.720 91.350 58.130 ;
        RECT 92.190 57.720 92.730 58.130 ;
        RECT 93.570 57.720 94.110 58.130 ;
        RECT 94.950 57.720 95.490 58.130 ;
        RECT 96.330 57.720 96.870 58.130 ;
        RECT 97.710 57.720 98.250 58.130 ;
        RECT 99.090 57.720 99.630 58.130 ;
        RECT 100.470 57.720 101.010 58.130 ;
        RECT 101.850 57.720 102.390 58.130 ;
        RECT 103.230 57.720 103.770 58.130 ;
        RECT 104.610 57.720 105.150 58.130 ;
        RECT 105.990 57.720 106.530 58.130 ;
        RECT 107.370 57.720 107.910 58.130 ;
        RECT 108.750 57.720 109.290 58.130 ;
        RECT 110.130 57.720 110.670 58.130 ;
        RECT 111.510 57.720 112.050 58.130 ;
        RECT 112.890 57.720 113.430 58.130 ;
        RECT 114.270 57.720 114.810 58.130 ;
        RECT 115.650 57.720 116.190 58.130 ;
        RECT 117.030 57.720 117.570 58.130 ;
        RECT 118.410 57.720 118.950 58.130 ;
        RECT 119.790 57.720 120.330 58.130 ;
        RECT 121.170 57.720 121.710 58.130 ;
        RECT 122.550 57.720 123.090 58.130 ;
        RECT 123.930 57.720 124.470 58.130 ;
        RECT 125.310 57.720 125.850 58.130 ;
        RECT 126.690 57.720 127.230 58.130 ;
        RECT 128.070 57.720 128.610 58.130 ;
        RECT 129.450 57.720 129.990 58.130 ;
        RECT 130.830 57.720 131.370 58.130 ;
        RECT 132.210 57.720 132.750 58.130 ;
        RECT 133.590 57.720 134.130 58.130 ;
        RECT 134.970 57.720 135.510 58.130 ;
        RECT 136.350 57.720 136.890 58.130 ;
        RECT 137.730 57.720 138.270 58.130 ;
        RECT 139.110 57.720 139.650 58.130 ;
        RECT 140.490 57.720 141.030 58.130 ;
        RECT 141.870 57.720 142.410 58.130 ;
        RECT 143.250 57.720 143.790 58.130 ;
        RECT 144.630 57.720 145.170 58.130 ;
        RECT 146.010 57.720 146.550 58.130 ;
        RECT 147.390 57.720 147.930 58.130 ;
        RECT 148.770 57.720 149.310 58.130 ;
        RECT 150.150 57.720 150.690 58.130 ;
        RECT 151.530 57.720 152.070 58.130 ;
        RECT 152.910 57.720 153.450 58.130 ;
        RECT 154.290 57.720 154.830 58.130 ;
        RECT 155.670 57.720 156.210 58.130 ;
        RECT 157.050 57.720 157.590 58.130 ;
        RECT 158.430 57.720 158.970 58.130 ;
        RECT 159.810 57.720 160.350 58.130 ;
        RECT 161.190 57.720 161.730 58.130 ;
        RECT 162.570 57.720 163.110 58.130 ;
        RECT 163.950 57.720 164.490 58.130 ;
        RECT 165.330 57.720 165.870 58.130 ;
        RECT 166.710 57.720 167.250 58.130 ;
        RECT 168.090 57.720 168.630 58.130 ;
        RECT 169.470 57.720 170.010 58.130 ;
        RECT 170.850 57.720 171.390 58.130 ;
        RECT 172.230 57.720 172.770 58.130 ;
        RECT 173.610 57.720 174.150 58.130 ;
        RECT 174.990 57.720 175.530 58.130 ;
        RECT 176.370 57.720 176.910 58.130 ;
        RECT 177.750 57.720 178.290 58.130 ;
        RECT 179.130 57.720 179.670 58.130 ;
        RECT 180.510 57.720 181.050 58.130 ;
        RECT 181.890 57.720 182.430 58.130 ;
        RECT 183.270 57.720 183.810 58.130 ;
        RECT 184.650 57.720 185.190 58.130 ;
        RECT 186.030 57.720 186.570 58.130 ;
        RECT 187.410 57.720 187.950 58.130 ;
        RECT 188.790 57.720 189.330 58.130 ;
        RECT 190.170 57.720 190.710 58.130 ;
        RECT 191.550 57.720 192.090 58.130 ;
        RECT 192.930 57.720 193.470 58.130 ;
        RECT 194.310 57.720 211.970 58.130 ;
        RECT 6.530 2.280 211.970 57.720 ;
        RECT 6.530 0.010 13.610 2.280 ;
        RECT 14.450 0.010 14.990 2.280 ;
        RECT 15.830 0.010 16.370 2.280 ;
        RECT 17.210 0.010 17.750 2.280 ;
        RECT 18.590 0.010 19.130 2.280 ;
        RECT 19.970 0.010 20.510 2.280 ;
        RECT 21.350 0.010 21.890 2.280 ;
        RECT 22.730 0.010 23.270 2.280 ;
        RECT 24.110 0.010 24.650 2.280 ;
        RECT 25.490 0.010 26.030 2.280 ;
        RECT 26.870 0.010 27.410 2.280 ;
        RECT 28.250 0.010 28.790 2.280 ;
        RECT 29.630 0.010 30.170 2.280 ;
        RECT 31.010 0.010 31.550 2.280 ;
        RECT 32.390 0.010 32.930 2.280 ;
        RECT 33.770 0.010 34.310 2.280 ;
        RECT 35.150 0.010 35.690 2.280 ;
        RECT 36.530 0.010 37.070 2.280 ;
        RECT 37.910 0.010 38.450 2.280 ;
        RECT 39.290 0.010 39.830 2.280 ;
        RECT 40.670 0.010 41.210 2.280 ;
        RECT 42.050 0.010 42.590 2.280 ;
        RECT 43.430 0.010 43.970 2.280 ;
        RECT 44.810 0.010 45.350 2.280 ;
        RECT 46.190 0.010 46.730 2.280 ;
        RECT 47.570 0.010 48.110 2.280 ;
        RECT 48.950 0.010 49.490 2.280 ;
        RECT 50.330 0.010 50.870 2.280 ;
        RECT 51.710 0.010 52.250 2.280 ;
        RECT 53.090 0.010 53.630 2.280 ;
        RECT 54.470 0.010 55.010 2.280 ;
        RECT 55.850 0.010 56.390 2.280 ;
        RECT 57.230 0.010 57.770 2.280 ;
        RECT 58.610 0.010 59.150 2.280 ;
        RECT 59.990 0.010 60.530 2.280 ;
        RECT 61.370 0.010 61.910 2.280 ;
        RECT 62.750 0.010 63.290 2.280 ;
        RECT 64.130 0.010 64.670 2.280 ;
        RECT 65.510 0.010 66.050 2.280 ;
        RECT 66.890 0.010 67.430 2.280 ;
        RECT 68.270 0.010 68.810 2.280 ;
        RECT 69.650 0.010 70.190 2.280 ;
        RECT 71.030 0.010 71.570 2.280 ;
        RECT 72.410 0.010 72.950 2.280 ;
        RECT 73.790 0.010 74.330 2.280 ;
        RECT 75.170 0.010 75.710 2.280 ;
        RECT 76.550 0.010 77.090 2.280 ;
        RECT 77.930 0.010 78.470 2.280 ;
        RECT 79.310 0.010 79.850 2.280 ;
        RECT 80.690 0.010 81.230 2.280 ;
        RECT 82.070 0.010 82.610 2.280 ;
        RECT 83.450 0.010 83.990 2.280 ;
        RECT 84.830 0.010 85.370 2.280 ;
        RECT 86.210 0.010 86.750 2.280 ;
        RECT 87.590 0.010 88.130 2.280 ;
        RECT 88.970 0.010 89.510 2.280 ;
        RECT 90.350 0.010 90.890 2.280 ;
        RECT 91.730 0.010 92.270 2.280 ;
        RECT 93.110 0.010 93.650 2.280 ;
        RECT 94.490 0.010 95.030 2.280 ;
        RECT 95.870 0.010 96.410 2.280 ;
        RECT 97.250 0.010 97.790 2.280 ;
        RECT 98.630 0.010 99.170 2.280 ;
        RECT 100.010 0.010 100.550 2.280 ;
        RECT 101.390 0.010 101.930 2.280 ;
        RECT 102.770 0.010 103.310 2.280 ;
        RECT 104.150 0.010 104.690 2.280 ;
        RECT 105.530 0.010 106.070 2.280 ;
        RECT 106.910 0.010 107.450 2.280 ;
        RECT 108.290 0.010 108.830 2.280 ;
        RECT 109.670 0.010 110.210 2.280 ;
        RECT 111.050 0.010 111.590 2.280 ;
        RECT 112.430 0.010 112.970 2.280 ;
        RECT 113.810 0.010 114.350 2.280 ;
        RECT 115.190 0.010 115.730 2.280 ;
        RECT 116.570 0.010 117.110 2.280 ;
        RECT 117.950 0.010 118.490 2.280 ;
        RECT 119.330 0.010 119.870 2.280 ;
        RECT 120.710 0.010 121.250 2.280 ;
        RECT 122.090 0.010 122.630 2.280 ;
        RECT 123.470 0.010 124.010 2.280 ;
        RECT 124.850 0.010 125.390 2.280 ;
        RECT 126.230 0.010 126.770 2.280 ;
        RECT 127.610 0.010 128.150 2.280 ;
        RECT 128.990 0.010 129.530 2.280 ;
        RECT 130.370 0.010 130.910 2.280 ;
        RECT 131.750 0.010 132.290 2.280 ;
        RECT 133.130 0.010 133.670 2.280 ;
        RECT 134.510 0.010 135.050 2.280 ;
        RECT 135.890 0.010 136.430 2.280 ;
        RECT 137.270 0.010 137.810 2.280 ;
        RECT 138.650 0.010 139.190 2.280 ;
        RECT 140.030 0.010 140.570 2.280 ;
        RECT 141.410 0.010 141.950 2.280 ;
        RECT 142.790 0.010 143.330 2.280 ;
        RECT 144.170 0.010 144.710 2.280 ;
        RECT 145.550 0.010 146.090 2.280 ;
        RECT 146.930 0.010 147.470 2.280 ;
        RECT 148.310 0.010 148.850 2.280 ;
        RECT 149.690 0.010 150.230 2.280 ;
        RECT 151.070 0.010 151.610 2.280 ;
        RECT 152.450 0.010 152.990 2.280 ;
        RECT 153.830 0.010 154.370 2.280 ;
        RECT 155.210 0.010 155.750 2.280 ;
        RECT 156.590 0.010 157.130 2.280 ;
        RECT 157.970 0.010 158.510 2.280 ;
        RECT 159.350 0.010 159.890 2.280 ;
        RECT 160.730 0.010 161.270 2.280 ;
        RECT 162.110 0.010 162.650 2.280 ;
        RECT 163.490 0.010 164.030 2.280 ;
        RECT 164.870 0.010 165.410 2.280 ;
        RECT 166.250 0.010 166.790 2.280 ;
        RECT 167.630 0.010 168.170 2.280 ;
        RECT 169.010 0.010 169.550 2.280 ;
        RECT 170.390 0.010 170.930 2.280 ;
        RECT 171.770 0.010 172.310 2.280 ;
        RECT 173.150 0.010 173.690 2.280 ;
        RECT 174.530 0.010 175.070 2.280 ;
        RECT 175.910 0.010 176.450 2.280 ;
        RECT 177.290 0.010 177.830 2.280 ;
        RECT 178.670 0.010 179.210 2.280 ;
        RECT 180.050 0.010 180.590 2.280 ;
        RECT 181.430 0.010 181.970 2.280 ;
        RECT 182.810 0.010 183.350 2.280 ;
        RECT 184.190 0.010 184.730 2.280 ;
        RECT 185.570 0.010 186.110 2.280 ;
        RECT 186.950 0.010 187.490 2.280 ;
        RECT 188.330 0.010 188.870 2.280 ;
        RECT 189.710 0.010 190.250 2.280 ;
        RECT 191.090 0.010 191.630 2.280 ;
        RECT 192.470 0.010 193.010 2.280 ;
        RECT 193.850 0.010 194.390 2.280 ;
        RECT 195.230 0.010 195.770 2.280 ;
        RECT 196.610 0.010 197.150 2.280 ;
        RECT 197.990 0.010 198.530 2.280 ;
        RECT 199.370 0.010 199.910 2.280 ;
        RECT 200.750 0.010 201.290 2.280 ;
        RECT 202.130 0.010 202.670 2.280 ;
        RECT 203.510 0.010 204.050 2.280 ;
        RECT 204.890 0.010 205.430 2.280 ;
        RECT 206.270 0.010 211.970 2.280 ;
      LAYER met3 ;
        RECT 6.510 2.555 211.995 57.285 ;
      LAYER met4 ;
        RECT 49.055 3.575 49.300 48.785 ;
        RECT 51.700 3.575 86.100 48.785 ;
        RECT 88.500 3.575 89.300 48.785 ;
        RECT 91.700 3.575 92.500 48.785 ;
        RECT 94.900 3.575 95.700 48.785 ;
        RECT 98.100 3.575 126.100 48.785 ;
        RECT 128.500 3.575 129.300 48.785 ;
        RECT 131.700 3.575 132.500 48.785 ;
        RECT 134.900 3.575 135.700 48.785 ;
        RECT 138.100 3.575 166.100 48.785 ;
        RECT 168.500 3.575 169.300 48.785 ;
        RECT 171.700 3.575 194.745 48.785 ;
  END
END mgmt_protect
END LIBRARY

