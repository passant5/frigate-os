VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gpio_control_block_mgmt_monitor
  CLASS BLOCK ;
  FOREIGN gpio_control_block_mgmt_monitor ;
  ORIGIN 0.000 0.000 ;
  SIZE 50.000 BY 74.000 ;
  PIN gpio_defaults[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 25.390 72.000 25.670 75.000 ;
    END
  END gpio_defaults[0]
  PIN gpio_defaults[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 39.190 72.000 39.470 75.000 ;
    END
  END gpio_defaults[10]
  PIN gpio_defaults[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 40.570 72.000 40.850 75.000 ;
    END
  END gpio_defaults[11]
  PIN gpio_defaults[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 72.000 42.230 75.000 ;
    END
  END gpio_defaults[12]
  PIN gpio_defaults[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 43.330 72.000 43.610 75.000 ;
    END
  END gpio_defaults[13]
  PIN gpio_defaults[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 72.000 44.990 75.000 ;
    END
  END gpio_defaults[14]
  PIN gpio_defaults[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 46.090 72.000 46.370 75.000 ;
    END
  END gpio_defaults[15]
  PIN gpio_defaults[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.770 72.000 27.050 75.000 ;
    END
  END gpio_defaults[1]
  PIN gpio_defaults[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 28.150 72.000 28.430 75.000 ;
    END
  END gpio_defaults[2]
  PIN gpio_defaults[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 29.530 72.000 29.810 75.000 ;
    END
  END gpio_defaults[3]
  PIN gpio_defaults[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 30.910 72.000 31.190 75.000 ;
    END
  END gpio_defaults[4]
  PIN gpio_defaults[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 32.290 72.000 32.570 75.000 ;
    END
  END gpio_defaults[5]
  PIN gpio_defaults[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 33.670 72.000 33.950 75.000 ;
    END
  END gpio_defaults[6]
  PIN gpio_defaults[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 35.050 72.000 35.330 75.000 ;
    END
  END gpio_defaults[7]
  PIN gpio_defaults[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 36.430 72.000 36.710 75.000 ;
    END
  END gpio_defaults[8]
  PIN gpio_defaults[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 37.810 72.000 38.090 75.000 ;
    END
  END gpio_defaults[9]
  PIN mgmt_gpio_in
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -1.000 25.880 2.000 26.480 ;
    END
  END mgmt_gpio_in
  PIN mgmt_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -1.000 34.040 2.000 34.640 ;
    END
  END mgmt_gpio_oeb
  PIN mgmt_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -1.000 29.960 2.000 30.560 ;
    END
  END mgmt_gpio_out
  PIN pad_gpio_ana_en
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 16.360 51.000 16.960 ;
    END
  END pad_gpio_ana_en
  PIN pad_gpio_ana_pol
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 28.600 51.000 29.200 ;
    END
  END pad_gpio_ana_pol
  PIN pad_gpio_ana_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 36.760 51.000 37.360 ;
    END
  END pad_gpio_ana_sel
  PIN pad_gpio_dm[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 20.440 51.000 21.040 ;
    END
  END pad_gpio_dm[0]
  PIN pad_gpio_dm[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 12.280 51.000 12.880 ;
    END
  END pad_gpio_dm[1]
  PIN pad_gpio_dm[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 49.000 51.000 49.600 ;
    END
  END pad_gpio_dm[2]
  PIN pad_gpio_holdover
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 53.080 51.000 53.680 ;
    END
  END pad_gpio_holdover
  PIN pad_gpio_hys_trim
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 44.920 51.000 45.520 ;
    END
  END pad_gpio_hys_trim
  PIN pad_gpio_ib_mode_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 65.320 51.000 65.920 ;
    END
  END pad_gpio_ib_mode_sel
  PIN pad_gpio_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT 48.000 4.120 51.000 4.720 ;
    END
  END pad_gpio_in
  PIN pad_gpio_inenb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 32.680 51.000 33.280 ;
    END
  END pad_gpio_inenb
  PIN pad_gpio_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 57.160 51.000 57.760 ;
    END
  END pad_gpio_out
  PIN pad_gpio_outenb
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 69.400 51.000 70.000 ;
    END
  END pad_gpio_outenb
  PIN pad_gpio_slew_ctl[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 24.520 51.000 25.120 ;
    END
  END pad_gpio_slew_ctl[0]
  PIN pad_gpio_slew_ctl[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 48.000 40.840 51.000 41.440 ;
    END
  END pad_gpio_slew_ctl[1]
  PIN pad_gpio_slow_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 8.200 51.000 8.800 ;
    END
  END pad_gpio_slow_sel
  PIN pad_gpio_vtrip_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT 48.000 61.240 51.000 61.840 ;
    END
  END pad_gpio_vtrip_sel
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639000 ;
    PORT
      LAYER met3 ;
        RECT -1.000 9.560 2.000 10.160 ;
    END
  END resetn
  PIN resetn_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT -1.000 50.360 2.000 50.960 ;
    END
  END resetn_out
  PIN serial_clock
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.465000 ;
    PORT
      LAYER met3 ;
        RECT -1.000 13.640 2.000 14.240 ;
    END
  END serial_clock
  PIN serial_clock_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT -1.000 54.440 2.000 55.040 ;
    END
  END serial_clock_out
  PIN serial_data_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -1.000 21.800 2.000 22.400 ;
    END
  END serial_data_in
  PIN serial_data_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -1.000 62.600 2.000 63.200 ;
    END
  END serial_data_out
  PIN serial_load
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.356000 ;
    PORT
      LAYER met3 ;
        RECT -1.000 17.720 2.000 18.320 ;
    END
  END serial_load
  PIN serial_load_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.590400 ;
    PORT
      LAYER met3 ;
        RECT -1.000 58.520 2.000 59.120 ;
    END
  END serial_load_out
  PIN user_gpio_in
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met3 ;
        RECT -1.000 46.280 2.000 46.880 ;
    END
  END user_gpio_in
  PIN user_gpio_oeb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -1.000 42.200 2.000 42.800 ;
    END
  END user_gpio_oeb
  PIN user_gpio_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met3 ;
        RECT -1.000 38.120 2.000 38.720 ;
    END
  END user_gpio_out
  PIN vccd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 12.720 20.470 13.720 70.960 ;
    END
    PORT
      LAYER met2 ;
        RECT 32.720 4.940 33.720 70.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 4.940 47.160 5.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 24.940 47.160 25.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 44.940 47.160 45.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 64.940 47.160 65.940 ;
    END
  END vccd
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 16.720 20.470 17.720 70.960 ;
    END
    PORT
      LAYER met2 ;
        RECT 36.720 5.200 37.720 70.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 8.940 47.160 9.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 28.940 47.160 29.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 48.940 47.160 49.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 68.940 47.160 69.940 ;
    END
  END vccd1
  PIN vssd
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 14.720 20.470 15.720 70.960 ;
    END
    PORT
      LAYER met2 ;
        RECT 34.720 5.200 35.720 70.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 6.940 47.160 7.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 26.940 47.160 27.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 46.940 47.160 47.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 66.940 47.160 67.940 ;
    END
  END vssd
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 18.720 5.200 19.720 70.960 ;
    END
    PORT
      LAYER met2 ;
        RECT 38.720 5.200 39.720 70.960 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 10.940 47.160 11.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 30.940 47.160 31.940 ;
    END
    PORT
      LAYER met3 ;
        RECT 2.980 50.940 47.160 51.940 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 2.810 5.355 47.110 70.805 ;
      LAYER li1 ;
        RECT 3.000 5.355 46.920 70.805 ;
      LAYER met1 ;
        RECT 1.910 5.200 48.230 71.700 ;
      LAYER met2 ;
        RECT 1.930 71.720 25.110 72.490 ;
        RECT 25.950 71.720 26.490 72.490 ;
        RECT 27.330 71.720 27.870 72.490 ;
        RECT 28.710 71.720 29.250 72.490 ;
        RECT 30.090 71.720 30.630 72.490 ;
        RECT 31.470 71.720 32.010 72.490 ;
        RECT 32.850 71.720 33.390 72.490 ;
        RECT 34.230 71.720 34.770 72.490 ;
        RECT 35.610 71.720 36.150 72.490 ;
        RECT 36.990 71.720 37.530 72.490 ;
        RECT 38.370 71.720 38.910 72.490 ;
        RECT 39.750 71.720 40.290 72.490 ;
        RECT 41.130 71.720 41.670 72.490 ;
        RECT 42.510 71.720 43.050 72.490 ;
        RECT 43.890 71.720 44.430 72.490 ;
        RECT 45.270 71.720 45.810 72.490 ;
        RECT 46.650 71.720 48.210 72.490 ;
        RECT 1.930 71.240 48.210 71.720 ;
        RECT 1.930 20.190 12.440 71.240 ;
        RECT 14.000 20.190 14.440 71.240 ;
        RECT 16.000 20.190 16.440 71.240 ;
        RECT 18.000 20.190 18.440 71.240 ;
        RECT 1.930 4.920 18.440 20.190 ;
        RECT 20.000 4.920 32.440 71.240 ;
        RECT 1.930 4.660 32.440 4.920 ;
        RECT 34.000 4.920 34.440 71.240 ;
        RECT 36.000 4.920 36.440 71.240 ;
        RECT 38.000 4.920 38.440 71.240 ;
        RECT 40.000 4.920 48.210 71.240 ;
        RECT 34.000 4.660 48.210 4.920 ;
        RECT 1.930 4.235 48.210 4.660 ;
      LAYER met3 ;
        RECT 1.905 68.540 2.580 69.865 ;
        RECT 47.560 69.000 47.600 69.865 ;
        RECT 47.560 68.540 48.000 69.000 ;
        RECT 1.905 68.340 48.000 68.540 ;
        RECT 1.905 66.540 2.580 68.340 ;
        RECT 47.560 66.540 48.000 68.340 ;
        RECT 1.905 66.340 48.000 66.540 ;
        RECT 1.905 64.540 2.580 66.340 ;
        RECT 47.560 66.320 48.000 66.340 ;
        RECT 47.560 64.920 47.600 66.320 ;
        RECT 47.560 64.540 48.000 64.920 ;
        RECT 1.905 63.600 48.000 64.540 ;
        RECT 2.400 62.240 48.000 63.600 ;
        RECT 2.400 62.200 47.600 62.240 ;
        RECT 1.905 60.840 47.600 62.200 ;
        RECT 1.905 59.520 48.000 60.840 ;
        RECT 2.400 58.160 48.000 59.520 ;
        RECT 2.400 58.120 47.600 58.160 ;
        RECT 1.905 56.760 47.600 58.120 ;
        RECT 1.905 55.440 48.000 56.760 ;
        RECT 2.400 54.080 48.000 55.440 ;
        RECT 2.400 54.040 47.600 54.080 ;
        RECT 1.905 52.680 47.600 54.040 ;
        RECT 1.905 52.340 48.000 52.680 ;
        RECT 1.905 51.360 2.580 52.340 ;
        RECT 2.400 50.540 2.580 51.360 ;
        RECT 47.560 50.540 48.000 52.340 ;
        RECT 2.400 50.340 48.000 50.540 ;
        RECT 2.400 49.960 2.580 50.340 ;
        RECT 1.905 48.540 2.580 49.960 ;
        RECT 47.560 50.000 48.000 50.340 ;
        RECT 47.560 48.600 47.600 50.000 ;
        RECT 47.560 48.540 48.000 48.600 ;
        RECT 1.905 48.340 48.000 48.540 ;
        RECT 1.905 47.280 2.580 48.340 ;
        RECT 2.400 46.540 2.580 47.280 ;
        RECT 47.560 46.540 48.000 48.340 ;
        RECT 2.400 46.340 48.000 46.540 ;
        RECT 2.400 45.880 2.580 46.340 ;
        RECT 1.905 44.540 2.580 45.880 ;
        RECT 47.560 45.920 48.000 46.340 ;
        RECT 47.560 44.540 47.600 45.920 ;
        RECT 1.905 44.520 47.600 44.540 ;
        RECT 1.905 43.200 48.000 44.520 ;
        RECT 2.400 41.840 48.000 43.200 ;
        RECT 2.400 41.800 47.600 41.840 ;
        RECT 1.905 40.440 47.600 41.800 ;
        RECT 1.905 39.120 48.000 40.440 ;
        RECT 2.400 37.760 48.000 39.120 ;
        RECT 2.400 37.720 47.600 37.760 ;
        RECT 1.905 36.360 47.600 37.720 ;
        RECT 1.905 35.040 48.000 36.360 ;
        RECT 2.400 33.680 48.000 35.040 ;
        RECT 2.400 33.640 47.600 33.680 ;
        RECT 1.905 32.340 47.600 33.640 ;
        RECT 1.905 30.960 2.580 32.340 ;
        RECT 2.400 30.540 2.580 30.960 ;
        RECT 47.560 32.280 47.600 32.340 ;
        RECT 47.560 30.540 48.000 32.280 ;
        RECT 2.400 30.340 48.000 30.540 ;
        RECT 2.400 29.560 2.580 30.340 ;
        RECT 1.905 28.540 2.580 29.560 ;
        RECT 47.560 29.600 48.000 30.340 ;
        RECT 47.560 28.540 47.600 29.600 ;
        RECT 1.905 28.340 47.600 28.540 ;
        RECT 1.905 26.880 2.580 28.340 ;
        RECT 2.400 26.540 2.580 26.880 ;
        RECT 47.560 28.200 47.600 28.340 ;
        RECT 47.560 26.540 48.000 28.200 ;
        RECT 2.400 26.340 48.000 26.540 ;
        RECT 2.400 25.480 2.580 26.340 ;
        RECT 1.905 24.540 2.580 25.480 ;
        RECT 47.560 25.520 48.000 26.340 ;
        RECT 47.560 24.540 47.600 25.520 ;
        RECT 1.905 24.120 47.600 24.540 ;
        RECT 1.905 22.800 48.000 24.120 ;
        RECT 2.400 21.440 48.000 22.800 ;
        RECT 2.400 21.400 47.600 21.440 ;
        RECT 1.905 20.040 47.600 21.400 ;
        RECT 1.905 18.720 48.000 20.040 ;
        RECT 2.400 17.360 48.000 18.720 ;
        RECT 2.400 17.320 47.600 17.360 ;
        RECT 1.905 15.960 47.600 17.320 ;
        RECT 1.905 14.640 48.000 15.960 ;
        RECT 2.400 13.280 48.000 14.640 ;
        RECT 2.400 13.240 47.600 13.280 ;
        RECT 1.905 12.340 47.600 13.240 ;
        RECT 1.905 10.560 2.580 12.340 ;
        RECT 2.400 10.540 2.580 10.560 ;
        RECT 47.560 11.880 47.600 12.340 ;
        RECT 47.560 10.540 48.000 11.880 ;
        RECT 2.400 10.340 48.000 10.540 ;
        RECT 2.400 9.160 2.580 10.340 ;
        RECT 1.905 8.540 2.580 9.160 ;
        RECT 47.560 9.200 48.000 10.340 ;
        RECT 47.560 8.540 47.600 9.200 ;
        RECT 1.905 8.340 47.600 8.540 ;
        RECT 1.905 6.540 2.580 8.340 ;
        RECT 47.560 7.800 47.600 8.340 ;
        RECT 47.560 6.540 48.000 7.800 ;
        RECT 1.905 6.340 48.000 6.540 ;
        RECT 1.905 4.540 2.580 6.340 ;
        RECT 47.560 5.120 48.000 6.340 ;
        RECT 47.560 4.540 47.600 5.120 ;
        RECT 1.905 4.255 47.600 4.540 ;
  END
END gpio_control_block_mgmt_monitor
END LIBRARY

