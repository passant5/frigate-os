module manual_power_connections ();
endmodule