magic
tech sky130A
magscale 1 2
timestamp 1750041009
<< viali >>
rect 24501 11305 24535 11339
rect 26709 11305 26743 11339
rect 27077 11305 27111 11339
rect 29009 11305 29043 11339
rect 30113 11305 30147 11339
rect 30297 11305 30331 11339
rect 31217 11305 31251 11339
rect 33701 11305 33735 11339
rect 33885 11305 33919 11339
rect 34161 11305 34195 11339
rect 29193 11237 29227 11271
rect 31769 11237 31803 11271
rect 24133 11169 24167 11203
rect 24317 11169 24351 11203
rect 25513 11169 25547 11203
rect 25697 11169 25731 11203
rect 25881 11169 25915 11203
rect 26065 11169 26099 11203
rect 26341 11169 26375 11203
rect 26525 11169 26559 11203
rect 27813 11169 27847 11203
rect 27997 11169 28031 11203
rect 28089 11169 28123 11203
rect 28273 11169 28307 11203
rect 28549 11169 28583 11203
rect 28733 11169 28767 11203
rect 29469 11169 29503 11203
rect 29653 11169 29687 11203
rect 29745 11169 29779 11203
rect 29929 11169 29963 11203
rect 30389 11169 30423 11203
rect 30573 11169 30607 11203
rect 30665 11169 30699 11203
rect 30849 11169 30883 11203
rect 31493 11169 31527 11203
rect 31677 11169 31711 11203
rect 32321 11169 32355 11203
rect 32496 11167 32530 11201
rect 32597 11169 32631 11203
rect 32781 11169 32815 11203
rect 32873 11169 32907 11203
rect 33057 11169 33091 11203
rect 33149 11169 33183 11203
rect 33333 11169 33367 11203
rect 26893 11101 26927 11135
rect 28457 11101 28491 11135
rect 31033 11101 31067 11135
rect 33517 11101 33551 11135
rect 25605 11033 25639 11067
rect 30757 11033 30791 11067
rect 31585 11033 31619 11067
rect 32413 11033 32447 11067
rect 32965 11033 32999 11067
rect 24225 10965 24259 10999
rect 25973 10965 26007 10999
rect 26433 10965 26467 10999
rect 27905 10965 27939 10999
rect 28181 10965 28215 10999
rect 28641 10965 28675 10999
rect 29561 10965 29595 10999
rect 29837 10965 29871 10999
rect 30481 10965 30515 10999
rect 32689 10965 32723 10999
rect 33241 10965 33275 10999
rect 24685 10761 24719 10795
rect 27905 10761 27939 10795
rect 32321 10761 32355 10795
rect 25421 10693 25455 10727
rect 25605 10625 25639 10659
rect 24317 10557 24351 10591
rect 24501 10557 24535 10591
rect 24777 10557 24811 10591
rect 24961 10557 24995 10591
rect 25053 10557 25087 10591
rect 25237 10557 25271 10591
rect 27537 10557 27571 10591
rect 27721 10557 27755 10591
rect 31953 10557 31987 10591
rect 32137 10557 32171 10591
rect 32045 10489 32079 10523
rect 24501 10421 24535 10455
rect 24869 10421 24903 10455
rect 25145 10421 25179 10455
rect 27721 10421 27755 10455
rect 14749 10217 14783 10251
rect 16681 10217 16715 10251
rect 17325 10217 17359 10251
rect 18245 10217 18279 10251
rect 20821 10217 20855 10251
rect 21281 10217 21315 10251
rect 24961 10217 24995 10251
rect 27813 10217 27847 10251
rect 28181 10217 28215 10251
rect 31309 10217 31343 10251
rect 32045 10217 32079 10251
rect 14657 10149 14691 10183
rect 17969 10149 18003 10183
rect 19901 10149 19935 10183
rect 30021 10149 30055 10183
rect 31033 10149 31067 10183
rect 20545 10081 20579 10115
rect 24593 10081 24627 10115
rect 24777 10081 24811 10115
rect 26893 10081 26927 10115
rect 27077 10081 27111 10115
rect 27169 10081 27203 10115
rect 27353 10081 27387 10115
rect 27468 10081 27502 10115
rect 27629 10081 27663 10115
rect 28917 10071 28951 10105
rect 29101 10081 29135 10115
rect 29193 10081 29227 10115
rect 29377 10081 29411 10115
rect 29929 10081 29963 10115
rect 30113 10081 30147 10115
rect 30665 10081 30699 10115
rect 30849 10081 30883 10115
rect 30941 10081 30975 10115
rect 31125 10081 31159 10115
rect 31677 10081 31711 10115
rect 31861 10081 31895 10115
rect 27997 10013 28031 10047
rect 29561 10013 29595 10047
rect 17509 9945 17543 9979
rect 20361 9945 20395 9979
rect 30297 9945 30331 9979
rect 31769 9945 31803 9979
rect 13921 9877 13955 9911
rect 14473 9877 14507 9911
rect 16129 9877 16163 9911
rect 16405 9877 16439 9911
rect 16865 9877 16899 9911
rect 17049 9877 17083 9911
rect 17785 9877 17819 9911
rect 19073 9877 19107 9911
rect 19441 9877 19475 9911
rect 19717 9877 19751 9911
rect 20729 9877 20763 9911
rect 24685 9877 24719 9911
rect 26985 9877 27019 9911
rect 27261 9877 27295 9911
rect 27537 9877 27571 9911
rect 29009 9877 29043 9911
rect 29285 9877 29319 9911
rect 29745 9877 29779 9911
rect 30757 9877 30791 9911
rect 31585 9877 31619 9911
rect 16313 9673 16347 9707
rect 16957 9673 16991 9707
rect 13185 9605 13219 9639
rect 15025 9605 15059 9639
rect 15945 9605 15979 9639
rect 18429 9605 18463 9639
rect 19165 9605 19199 9639
rect 20177 9605 20211 9639
rect 22661 9605 22695 9639
rect 23213 9605 23247 9639
rect 24317 9605 24351 9639
rect 25513 9605 25547 9639
rect 28549 9605 28583 9639
rect 13553 9537 13587 9571
rect 14013 9537 14047 9571
rect 14565 9537 14599 9571
rect 15393 9537 15427 9571
rect 18061 9537 18095 9571
rect 19533 9537 19567 9571
rect 20085 9537 20119 9571
rect 20637 9537 20671 9571
rect 21189 9537 21223 9571
rect 21373 9537 21407 9571
rect 21925 9537 21959 9571
rect 23949 9537 23983 9571
rect 24593 9537 24627 9571
rect 14105 9469 14139 9503
rect 16037 9469 16071 9503
rect 16129 9469 16163 9503
rect 17141 9469 17175 9503
rect 17233 9469 17267 9503
rect 17509 9469 17543 9503
rect 17601 9469 17635 9503
rect 18889 9469 18923 9503
rect 19625 9469 19659 9503
rect 20729 9469 20763 9503
rect 22109 9469 22143 9503
rect 23857 9469 23891 9503
rect 28181 9469 28215 9503
rect 28365 9469 28399 9503
rect 14749 9401 14783 9435
rect 15577 9401 15611 9435
rect 22569 9401 22603 9435
rect 25421 9401 25455 9435
rect 13829 9333 13863 9367
rect 15209 9333 15243 9367
rect 15761 9333 15795 9367
rect 17417 9333 17451 9367
rect 18153 9333 18187 9367
rect 18613 9333 18647 9367
rect 19073 9333 19107 9367
rect 19441 9333 19475 9367
rect 20453 9333 20487 9367
rect 21465 9333 21499 9367
rect 21741 9333 21775 9367
rect 23489 9333 23523 9367
rect 24133 9333 24167 9367
rect 24777 9333 24811 9367
rect 28365 9333 28399 9367
rect 11621 9129 11655 9163
rect 16129 9129 16163 9163
rect 27077 9129 27111 9163
rect 10517 9061 10551 9095
rect 11437 9061 11471 9095
rect 13001 9061 13035 9095
rect 14473 9061 14507 9095
rect 15117 9061 15151 9095
rect 17785 9061 17819 9095
rect 18429 9061 18463 9095
rect 18521 9061 18555 9095
rect 19717 9061 19751 9095
rect 20361 9061 20395 9095
rect 21005 9061 21039 9095
rect 21833 9061 21867 9095
rect 21925 9061 21959 9095
rect 23213 9061 23247 9095
rect 23949 9061 23983 9095
rect 24869 9061 24903 9095
rect 10885 8993 10919 9027
rect 10977 8993 11011 9027
rect 12449 8993 12483 9027
rect 12561 8993 12595 9027
rect 13737 8993 13771 9027
rect 13829 8993 13863 9027
rect 13921 8993 13955 9027
rect 14013 8993 14047 9027
rect 14657 8993 14691 9027
rect 15209 8993 15243 9027
rect 15669 8993 15703 9027
rect 17049 8993 17083 9027
rect 17233 8993 17267 9027
rect 17325 8993 17359 9027
rect 17969 8993 18003 9027
rect 18981 8993 19015 9027
rect 19165 8993 19199 9027
rect 19257 8993 19291 9027
rect 19901 8993 19935 9027
rect 20453 8993 20487 9027
rect 20545 8993 20579 9027
rect 21281 8993 21315 9027
rect 21373 8993 21407 9027
rect 22385 8993 22419 9027
rect 22661 8993 22695 9027
rect 22753 8993 22787 9027
rect 23765 8993 23799 9027
rect 23857 8993 23891 9027
rect 24409 8993 24443 9027
rect 25329 8993 25363 9027
rect 25421 8993 25455 9027
rect 25932 8993 25966 9027
rect 26065 8993 26099 9027
rect 26709 8993 26743 9027
rect 26893 8993 26927 9027
rect 11805 8925 11839 8959
rect 14565 8925 14599 8959
rect 15761 8925 15795 8959
rect 17141 8925 17175 8959
rect 17877 8925 17911 8959
rect 19073 8925 19107 8959
rect 19809 8925 19843 8959
rect 22477 8925 22511 8959
rect 24501 8925 24535 8959
rect 24685 8925 24719 8959
rect 25513 8925 25547 8959
rect 26525 8925 26559 8959
rect 10333 8857 10367 8891
rect 16313 8857 16347 8891
rect 10609 8789 10643 8823
rect 11897 8789 11931 8823
rect 12081 8789 12115 8823
rect 12265 8789 12299 8823
rect 13185 8789 13219 8823
rect 13553 8789 13587 8823
rect 16405 8789 16439 8823
rect 16865 8789 16899 8823
rect 23581 8789 23615 8823
rect 26341 8789 26375 8823
rect 26801 8789 26835 8823
rect 6469 8585 6503 8619
rect 7573 8585 7607 8619
rect 8401 8585 8435 8619
rect 9229 8585 9263 8619
rect 10057 8585 10091 8619
rect 10977 8585 11011 8619
rect 11989 8585 12023 8619
rect 12357 8585 12391 8619
rect 14289 8585 14323 8619
rect 16313 8585 16347 8619
rect 16865 8585 16899 8619
rect 17417 8585 17451 8619
rect 18061 8585 18095 8619
rect 18981 8585 19015 8619
rect 19625 8585 19659 8619
rect 21005 8585 21039 8619
rect 21557 8585 21591 8619
rect 22845 8585 22879 8619
rect 26617 8585 26651 8619
rect 27169 8585 27203 8619
rect 9781 8517 9815 8551
rect 13737 8517 13771 8551
rect 17049 8517 17083 8551
rect 10149 8449 10183 8483
rect 10701 8449 10735 8483
rect 11069 8449 11103 8483
rect 11621 8449 11655 8483
rect 11805 8449 11839 8483
rect 13277 8449 13311 8483
rect 13921 8449 13955 8483
rect 14555 8449 14589 8483
rect 14657 8449 14691 8483
rect 15209 8449 15243 8483
rect 15301 8449 15335 8483
rect 15853 8449 15887 8483
rect 17693 8449 17727 8483
rect 18705 8449 18739 8483
rect 19349 8449 19383 8483
rect 20545 8449 20579 8483
rect 21925 8449 21959 8483
rect 22477 8449 22511 8483
rect 23213 8449 23247 8483
rect 24317 8449 24351 8483
rect 26065 8449 26099 8483
rect 7665 8381 7699 8415
rect 9321 8381 9355 8415
rect 9689 8381 9723 8415
rect 10609 8381 10643 8415
rect 11161 8381 11195 8415
rect 12541 8381 12575 8415
rect 12633 8381 12667 8415
rect 12725 8381 12759 8415
rect 12817 8381 12851 8415
rect 14473 8381 14507 8415
rect 14749 8381 14783 8415
rect 15393 8381 15427 8415
rect 16497 8381 16531 8415
rect 16589 8381 16623 8415
rect 17601 8381 17635 8415
rect 18245 8381 18279 8415
rect 18337 8381 18371 8415
rect 18797 8381 18831 8415
rect 19441 8381 19475 8415
rect 20453 8381 20487 8415
rect 20729 8381 20763 8415
rect 21741 8381 21775 8415
rect 21833 8381 21867 8415
rect 22017 8381 22051 8415
rect 23029 8381 23063 8415
rect 23121 8381 23155 8415
rect 24225 8381 24259 8415
rect 24869 8381 24903 8415
rect 24961 8381 24995 8415
rect 25053 8381 25087 8415
rect 25513 8381 25547 8415
rect 25605 8381 25639 8415
rect 26801 8381 26835 8415
rect 26893 8381 26927 8415
rect 6653 8313 6687 8347
rect 8585 8313 8619 8347
rect 13461 8313 13495 8347
rect 19993 8313 20027 8347
rect 23397 8313 23431 8347
rect 23765 8313 23799 8347
rect 24409 8313 24443 8347
rect 25881 8313 25915 8347
rect 26985 8313 27019 8347
rect 5549 8245 5583 8279
rect 5825 8245 5859 8279
rect 25697 8245 25731 8279
rect 4445 8041 4479 8075
rect 5549 8041 5583 8075
rect 6745 8041 6779 8075
rect 7481 8041 7515 8075
rect 9137 8041 9171 8075
rect 10977 8041 11011 8075
rect 6285 7973 6319 8007
rect 7389 7973 7423 8007
rect 8217 7973 8251 8007
rect 9045 7973 9079 8007
rect 9321 7973 9355 8007
rect 5181 7905 5215 7939
rect 5825 7905 5859 7939
rect 6929 7905 6963 7939
rect 7757 7905 7791 7939
rect 8585 7905 8619 7939
rect 9781 7905 9815 7939
rect 9873 7905 9907 7939
rect 10057 7905 10091 7939
rect 10241 7905 10275 7939
rect 5273 7837 5307 7871
rect 5733 7837 5767 7871
rect 6837 7837 6871 7871
rect 7665 7837 7699 7871
rect 8493 7837 8527 7871
rect 10149 7837 10183 7871
rect 10701 7837 10735 7871
rect 4169 7701 4203 7735
rect 4629 7701 4663 7735
rect 4997 7701 5031 7735
rect 6469 7701 6503 7735
rect 8309 7701 8343 7735
rect 11161 7701 11195 7735
rect 4629 7497 4663 7531
rect 5917 7497 5951 7531
rect 8585 7497 8619 7531
rect 8953 7497 8987 7531
rect 10977 7497 11011 7531
rect 3709 7361 3743 7395
rect 4261 7361 4295 7395
rect 4905 7361 4939 7395
rect 4997 7361 5031 7395
rect 5549 7361 5583 7395
rect 6837 7361 6871 7395
rect 7481 7361 7515 7395
rect 7573 7361 7607 7395
rect 8125 7361 8159 7395
rect 9229 7361 9263 7395
rect 9873 7361 9907 7395
rect 9965 7361 9999 7395
rect 11253 7361 11287 7395
rect 32781 7361 32815 7395
rect 33333 7361 33367 7395
rect 3801 7293 3835 7327
rect 4813 7293 4847 7327
rect 5089 7293 5123 7327
rect 6101 7293 6135 7327
rect 6193 7293 6227 7327
rect 6285 7293 6319 7327
rect 6377 7293 6411 7327
rect 6929 7293 6963 7327
rect 7021 7293 7055 7327
rect 7665 7293 7699 7327
rect 9137 7293 9171 7327
rect 9321 7293 9355 7327
rect 9413 7293 9447 7327
rect 10057 7293 10091 7327
rect 10517 7293 10551 7327
rect 11161 7293 11195 7327
rect 32873 7293 32907 7327
rect 33425 7293 33459 7327
rect 3525 7157 3559 7191
rect 8309 7157 8343 7191
rect 4537 6953 4571 6987
rect 6009 6953 6043 6987
rect 4997 6817 5031 6851
rect 5457 6817 5491 6851
rect 6377 6817 6411 6851
rect 6837 6817 6871 6851
rect 7021 6817 7055 6851
rect 7205 6817 7239 6851
rect 7665 6817 7699 6851
rect 8677 6817 8711 6851
rect 8769 6817 8803 6851
rect 8953 6817 8987 6851
rect 9505 6817 9539 6851
rect 9597 6817 9631 6851
rect 10261 6817 10295 6851
rect 11161 6817 11195 6851
rect 32873 6817 32907 6851
rect 32965 6817 32999 6851
rect 33425 6817 33459 6851
rect 33977 6817 34011 6851
rect 34621 6817 34655 6851
rect 34805 6817 34839 6851
rect 4353 6749 4387 6783
rect 4905 6749 4939 6783
rect 5733 6749 5767 6783
rect 6285 6749 6319 6783
rect 7113 6749 7147 6783
rect 8861 6749 8895 6783
rect 10057 6749 10091 6783
rect 10149 6749 10183 6783
rect 10701 6749 10735 6783
rect 10977 6749 11011 6783
rect 33517 6749 33551 6783
rect 34345 6749 34379 6783
rect 4721 6681 4755 6715
rect 6101 6681 6135 6715
rect 4169 6613 4203 6647
rect 7849 6613 7883 6647
rect 8125 6613 8159 6647
rect 8493 6613 8527 6647
rect 9137 6613 9171 6647
rect 5641 6409 5675 6443
rect 7849 6409 7883 6443
rect 8401 6409 8435 6443
rect 9505 6273 9539 6307
rect 10333 6273 10367 6307
rect 10701 6273 10735 6307
rect 11253 6273 11287 6307
rect 33057 6273 33091 6307
rect 34621 6273 34655 6307
rect 8953 6205 8987 6239
rect 9045 6205 9079 6239
rect 9781 6205 9815 6239
rect 9873 6205 9907 6239
rect 10793 6205 10827 6239
rect 33149 6205 33183 6239
rect 33609 6205 33643 6239
rect 34253 6205 34287 6239
rect 34897 6205 34931 6239
rect 35173 6205 35207 6239
rect 35633 6205 35667 6239
rect 7389 6137 7423 6171
rect 8493 6137 8527 6171
rect 10609 6137 10643 6171
rect 6929 6069 6963 6103
rect 8677 6069 8711 6103
rect 9689 6069 9723 6103
rect 32873 6069 32907 6103
rect 35725 6069 35759 6103
rect 36001 6069 36035 6103
rect 9781 5865 9815 5899
rect 10241 5865 10275 5899
rect 10517 5865 10551 5899
rect 11253 5865 11287 5899
rect 9597 5797 9631 5831
rect 9873 5593 9907 5627
rect 9321 5525 9355 5559
rect 33149 5185 33183 5219
rect 33333 5117 33367 5151
rect 36001 5117 36035 5151
rect 32965 5049 32999 5083
rect 32781 4981 32815 5015
rect 33977 4981 34011 5015
rect 36093 4981 36127 5015
rect 36369 4981 36403 5015
rect 32781 4641 32815 4675
rect 33149 4641 33183 4675
rect 33241 4641 33275 4675
rect 33701 4641 33735 4675
rect 34529 4641 34563 4675
rect 35173 4641 35207 4675
rect 35357 4641 35391 4675
rect 33793 4573 33827 4607
rect 34897 4573 34931 4607
rect 32873 4505 32907 4539
rect 33977 4437 34011 4471
rect 34345 4437 34379 4471
rect 35633 4437 35667 4471
rect 34345 4233 34379 4267
rect 37105 4233 37139 4267
rect 34529 4165 34563 4199
rect 36001 4165 36035 4199
rect 34897 4097 34931 4131
rect 36185 4097 36219 4131
rect 36461 4097 36495 4131
rect 32781 4029 32815 4063
rect 33057 4029 33091 4063
rect 33425 4029 33459 4063
rect 33517 4029 33551 4063
rect 34069 4029 34103 4063
rect 35633 4029 35667 4063
rect 35909 4029 35943 4063
rect 32873 3961 32907 3995
rect 33977 3961 34011 3995
rect 36553 3961 36587 3995
rect 37013 3961 37047 3995
rect 33149 3893 33183 3927
rect 34161 3893 34195 3927
rect 34713 3893 34747 3927
rect 35173 3893 35207 3927
rect 35449 3893 35483 3927
rect 36737 3893 36771 3927
rect 34345 3689 34379 3723
rect 37933 3689 37967 3723
rect 36829 3621 36863 3655
rect 32965 3553 32999 3587
rect 34253 3553 34287 3587
rect 34529 3553 34563 3587
rect 34805 3553 34839 3587
rect 35357 3553 35391 3587
rect 35725 3553 35759 3587
rect 36369 3553 36403 3587
rect 36921 3553 36955 3587
rect 37013 3553 37047 3587
rect 38117 3553 38151 3587
rect 33977 3485 34011 3519
rect 35633 3485 35667 3519
rect 36277 3485 36311 3519
rect 37473 3485 37507 3519
rect 37749 3417 37783 3451
rect 34621 3349 34655 3383
rect 34897 3349 34931 3383
rect 35909 3349 35943 3383
rect 31033 3145 31067 3179
rect 33793 3145 33827 3179
rect 36737 3145 36771 3179
rect 38669 3077 38703 3111
rect 29837 3009 29871 3043
rect 30757 3009 30791 3043
rect 34529 3009 34563 3043
rect 37473 3009 37507 3043
rect 38485 3009 38519 3043
rect 27721 2941 27755 2975
rect 28457 2941 28491 2975
rect 28733 2941 28767 2975
rect 30297 2941 30331 2975
rect 30389 2941 30423 2975
rect 30665 2941 30699 2975
rect 30941 2941 30975 2975
rect 32689 2941 32723 2975
rect 32965 2941 32999 2975
rect 33241 2941 33275 2975
rect 33517 2941 33551 2975
rect 34253 2941 34287 2975
rect 35541 2941 35575 2975
rect 35633 2941 35667 2975
rect 36185 2941 36219 2975
rect 36645 2941 36679 2975
rect 37197 2941 37231 2975
rect 37565 2941 37599 2975
rect 38025 2941 38059 2975
rect 38301 2941 38335 2975
rect 26065 2873 26099 2907
rect 26525 2873 26559 2907
rect 27813 2873 27847 2907
rect 28365 2873 28399 2907
rect 30481 2873 30515 2907
rect 31769 2873 31803 2907
rect 33057 2873 33091 2907
rect 33609 2873 33643 2907
rect 36093 2873 36127 2907
rect 25973 2805 26007 2839
rect 27997 2805 28031 2839
rect 28641 2805 28675 2839
rect 31217 2805 31251 2839
rect 33333 2805 33367 2839
rect 36277 2805 36311 2839
rect 38117 2805 38151 2839
rect 38853 2805 38887 2839
rect 38945 2601 38979 2635
rect 39865 2601 39899 2635
rect 26525 2533 26559 2567
rect 30205 2533 30239 2567
rect 35633 2533 35667 2567
rect 25605 2465 25639 2499
rect 27721 2465 27755 2499
rect 29009 2465 29043 2499
rect 29285 2465 29319 2499
rect 30757 2465 30791 2499
rect 31033 2465 31067 2499
rect 31493 2465 31527 2499
rect 33057 2465 33091 2499
rect 34621 2465 34655 2499
rect 35909 2465 35943 2499
rect 36001 2465 36035 2499
rect 36461 2465 36495 2499
rect 36645 2465 36679 2499
rect 37289 2465 37323 2499
rect 37473 2465 37507 2499
rect 38117 2465 38151 2499
rect 38301 2465 38335 2499
rect 38393 2465 38427 2499
rect 24593 2397 24627 2431
rect 25881 2397 25915 2431
rect 27997 2397 28031 2431
rect 31953 2397 31987 2431
rect 33425 2397 33459 2431
rect 37013 2397 37047 2431
rect 37841 2397 37875 2431
rect 38853 2397 38887 2431
rect 39497 2329 39531 2363
rect 40233 2329 40267 2363
rect 26065 2261 26099 2295
rect 30849 2261 30883 2295
rect 31125 2261 31159 2295
rect 39129 2261 39163 2295
rect 39313 2261 39347 2295
rect 39681 2261 39715 2295
rect 40049 2261 40083 2295
rect 40509 2261 40543 2295
rect 28365 2057 28399 2091
rect 39589 2057 39623 2091
rect 39865 2057 39899 2091
rect 40877 2057 40911 2091
rect 39313 1989 39347 2023
rect 40141 1989 40175 2023
rect 25789 1921 25823 1955
rect 33057 1921 33091 1955
rect 33333 1921 33367 1955
rect 34621 1921 34655 1955
rect 36001 1921 36035 1955
rect 37381 1921 37415 1955
rect 38209 1921 38243 1955
rect 25053 1853 25087 1887
rect 25513 1853 25547 1887
rect 26801 1853 26835 1887
rect 28273 1853 28307 1887
rect 28549 1853 28583 1887
rect 30297 1853 30331 1887
rect 30389 1853 30423 1887
rect 31861 1853 31895 1887
rect 33425 1853 33459 1887
rect 33885 1853 33919 1887
rect 34069 1853 34103 1887
rect 35541 1853 35575 1887
rect 37013 1853 37047 1887
rect 37749 1853 37783 1887
rect 37841 1853 37875 1887
rect 38577 1853 38611 1887
rect 38669 1855 38703 1889
rect 39221 1853 39255 1887
rect 39497 1853 39531 1887
rect 39773 1853 39807 1887
rect 40049 1853 40083 1887
rect 41061 1853 41095 1887
rect 24041 1785 24075 1819
rect 27905 1785 27939 1819
rect 29101 1785 29135 1819
rect 31401 1785 31435 1819
rect 40509 1785 40543 1819
rect 28641 1717 28675 1751
rect 38761 1717 38795 1751
rect 38945 1717 38979 1751
rect 40325 1717 40359 1751
rect 40693 1717 40727 1751
rect 41245 1717 41279 1751
rect 25145 1513 25179 1547
rect 25973 1513 26007 1547
rect 41245 1513 41279 1547
rect 25605 1445 25639 1479
rect 28733 1445 28767 1479
rect 35357 1445 35391 1479
rect 40877 1445 40911 1479
rect 23581 1377 23615 1411
rect 25237 1377 25271 1411
rect 25697 1377 25731 1411
rect 26065 1377 26099 1411
rect 26341 1377 26375 1411
rect 27445 1377 27479 1411
rect 27997 1377 28031 1411
rect 29285 1377 29319 1411
rect 30849 1377 30883 1411
rect 31493 1377 31527 1411
rect 32965 1377 32999 1411
rect 34437 1377 34471 1411
rect 36001 1377 36035 1411
rect 36645 1377 36679 1411
rect 37197 1377 37231 1411
rect 37473 1377 37507 1411
rect 38025 1377 38059 1411
rect 38301 1377 38335 1411
rect 39037 1377 39071 1411
rect 39129 1377 39163 1411
rect 39865 1377 39899 1411
rect 40049 1377 40083 1411
rect 40509 1377 40543 1411
rect 40785 1377 40819 1411
rect 24041 1309 24075 1343
rect 29745 1309 29779 1343
rect 30757 1309 30791 1343
rect 31309 1309 31343 1343
rect 32689 1309 32723 1343
rect 33425 1309 33459 1343
rect 35909 1309 35943 1343
rect 36461 1309 36495 1343
rect 37841 1309 37875 1343
rect 38669 1309 38703 1343
rect 39497 1309 39531 1343
rect 40325 1309 40359 1343
rect 41797 1309 41831 1343
rect 23397 1241 23431 1275
rect 42165 1241 42199 1275
rect 25329 1173 25363 1207
rect 36737 1173 36771 1207
rect 41061 1173 41095 1207
rect 41429 1173 41463 1207
rect 41981 1173 42015 1207
rect 23213 969 23247 1003
rect 25329 969 25363 1003
rect 25881 969 25915 1003
rect 27905 969 27939 1003
rect 28181 969 28215 1003
rect 30757 969 30791 1003
rect 31217 969 31251 1003
rect 33057 969 33091 1003
rect 36369 969 36403 1003
rect 41337 969 41371 1003
rect 41797 969 41831 1003
rect 26065 901 26099 935
rect 30481 901 30515 935
rect 40233 901 40267 935
rect 23029 833 23063 867
rect 24225 833 24259 867
rect 26801 833 26835 867
rect 33333 833 33367 867
rect 33885 833 33919 867
rect 35909 833 35943 867
rect 39773 833 39807 867
rect 41061 833 41095 867
rect 23305 765 23339 799
rect 23581 765 23615 799
rect 23765 765 23799 799
rect 25237 765 25271 799
rect 25513 765 25547 799
rect 25789 765 25823 799
rect 26341 765 26375 799
rect 27813 765 27847 799
rect 28089 765 28123 799
rect 28365 765 28399 799
rect 28457 765 28491 799
rect 28917 765 28951 799
rect 30389 765 30423 799
rect 30665 765 30699 799
rect 30941 765 30975 799
rect 31033 765 31067 799
rect 31493 765 31527 799
rect 32965 765 32999 799
rect 33425 765 33459 799
rect 34069 765 34103 799
rect 35541 765 35575 799
rect 36277 765 36311 799
rect 36645 765 36679 799
rect 38117 765 38151 799
rect 38485 765 38519 799
rect 38669 765 38703 799
rect 39221 765 39255 799
rect 39313 765 39347 799
rect 39865 765 39899 799
rect 40141 765 40175 799
rect 40417 765 40451 799
rect 40509 765 40543 799
rect 40693 765 40727 799
rect 40961 767 40995 801
rect 41245 765 41279 799
rect 42165 765 42199 799
rect 42349 765 42383 799
rect 23489 697 23523 731
rect 28641 697 28675 731
rect 29837 697 29871 731
rect 32689 697 32723 731
rect 35265 697 35299 731
rect 37565 697 37599 731
rect 42533 697 42567 731
rect 25605 629 25639 663
rect 38945 629 38979 663
rect 39957 629 39991 663
rect 40785 629 40819 663
rect 41521 629 41555 663
rect 41981 629 42015 663
<< metal1 >>
rect 31754 11568 31760 11620
rect 31812 11608 31818 11620
rect 32674 11608 32680 11620
rect 31812 11580 32680 11608
rect 31812 11568 31818 11580
rect 32674 11568 32680 11580
rect 32732 11568 32738 11620
rect 10042 11500 10048 11552
rect 10100 11540 10106 11552
rect 10410 11540 10416 11552
rect 10100 11512 10416 11540
rect 10100 11500 10106 11512
rect 10410 11500 10416 11512
rect 10468 11500 10474 11552
rect 18046 11500 18052 11552
rect 18104 11540 18110 11552
rect 18690 11540 18696 11552
rect 18104 11512 18696 11540
rect 18104 11500 18110 11512
rect 18690 11500 18696 11512
rect 18748 11500 18754 11552
rect 25866 11500 25872 11552
rect 25924 11540 25930 11552
rect 26050 11540 26056 11552
rect 25924 11512 26056 11540
rect 25924 11500 25930 11512
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 30098 11500 30104 11552
rect 30156 11540 30162 11552
rect 30742 11540 30748 11552
rect 30156 11512 30748 11540
rect 30156 11500 30162 11512
rect 30742 11500 30748 11512
rect 30800 11500 30806 11552
rect 31386 11500 31392 11552
rect 31444 11540 31450 11552
rect 32122 11540 32128 11552
rect 31444 11512 32128 11540
rect 31444 11500 31450 11512
rect 32122 11500 32128 11512
rect 32180 11500 32186 11552
rect 32214 11500 32220 11552
rect 32272 11540 32278 11552
rect 33502 11540 33508 11552
rect 32272 11512 33508 11540
rect 32272 11500 32278 11512
rect 33502 11500 33508 11512
rect 33560 11500 33566 11552
rect 460 11450 43516 11472
rect 460 11398 1946 11450
rect 1998 11398 2010 11450
rect 2062 11398 2074 11450
rect 2126 11398 2138 11450
rect 2190 11398 2202 11450
rect 2254 11398 9946 11450
rect 9998 11398 10010 11450
rect 10062 11398 10074 11450
rect 10126 11398 10138 11450
rect 10190 11398 10202 11450
rect 10254 11398 17946 11450
rect 17998 11398 18010 11450
rect 18062 11398 18074 11450
rect 18126 11398 18138 11450
rect 18190 11398 18202 11450
rect 18254 11398 25946 11450
rect 25998 11398 26010 11450
rect 26062 11398 26074 11450
rect 26126 11398 26138 11450
rect 26190 11398 26202 11450
rect 26254 11398 33946 11450
rect 33998 11398 34010 11450
rect 34062 11398 34074 11450
rect 34126 11398 34138 11450
rect 34190 11398 34202 11450
rect 34254 11398 41946 11450
rect 41998 11398 42010 11450
rect 42062 11398 42074 11450
rect 42126 11398 42138 11450
rect 42190 11398 42202 11450
rect 42254 11398 43516 11450
rect 460 11376 43516 11398
rect 24489 11339 24547 11345
rect 24489 11305 24501 11339
rect 24535 11336 24547 11339
rect 25498 11336 25504 11348
rect 24535 11308 25504 11336
rect 24535 11305 24547 11308
rect 24489 11299 24547 11305
rect 24504 11268 24532 11299
rect 25498 11296 25504 11308
rect 25556 11296 25562 11348
rect 26697 11339 26755 11345
rect 26697 11305 26709 11339
rect 26743 11336 26755 11339
rect 26878 11336 26884 11348
rect 26743 11308 26884 11336
rect 26743 11305 26755 11308
rect 26697 11299 26755 11305
rect 26712 11268 26740 11299
rect 26878 11296 26884 11308
rect 26936 11296 26942 11348
rect 27065 11339 27123 11345
rect 27065 11305 27077 11339
rect 27111 11336 27123 11339
rect 27430 11336 27436 11348
rect 27111 11308 27436 11336
rect 27111 11305 27123 11308
rect 27065 11299 27123 11305
rect 24136 11240 24532 11268
rect 25700 11240 26740 11268
rect 24136 11209 24164 11240
rect 24121 11203 24179 11209
rect 24121 11169 24133 11203
rect 24167 11169 24179 11203
rect 24121 11163 24179 11169
rect 24302 11160 24308 11212
rect 24360 11200 24366 11212
rect 25700 11209 25728 11240
rect 25501 11203 25559 11209
rect 25501 11200 25513 11203
rect 24360 11172 25513 11200
rect 24360 11160 24366 11172
rect 25501 11169 25513 11172
rect 25547 11169 25559 11203
rect 25501 11163 25559 11169
rect 25685 11203 25743 11209
rect 25685 11169 25697 11203
rect 25731 11169 25743 11203
rect 25685 11163 25743 11169
rect 25869 11203 25927 11209
rect 25869 11169 25881 11203
rect 25915 11200 25927 11203
rect 25958 11200 25964 11212
rect 25915 11172 25964 11200
rect 25915 11169 25927 11172
rect 25869 11163 25927 11169
rect 25516 11132 25544 11163
rect 25884 11132 25912 11163
rect 25958 11160 25964 11172
rect 26016 11160 26022 11212
rect 26053 11203 26111 11209
rect 26053 11169 26065 11203
rect 26099 11198 26111 11203
rect 26099 11170 26188 11198
rect 26099 11169 26111 11170
rect 26053 11163 26111 11169
rect 25516 11104 25912 11132
rect 26160 11132 26188 11170
rect 26234 11160 26240 11212
rect 26292 11200 26298 11212
rect 26329 11203 26387 11209
rect 26329 11200 26341 11203
rect 26292 11172 26341 11200
rect 26292 11160 26298 11172
rect 26329 11169 26341 11172
rect 26375 11169 26387 11203
rect 26329 11163 26387 11169
rect 26513 11203 26571 11209
rect 26513 11169 26525 11203
rect 26559 11200 26571 11203
rect 27080 11200 27108 11299
rect 27430 11296 27436 11308
rect 27488 11296 27494 11348
rect 28626 11336 28632 11348
rect 28092 11308 28632 11336
rect 28092 11268 28120 11308
rect 28626 11296 28632 11308
rect 28684 11296 28690 11348
rect 28997 11339 29055 11345
rect 28997 11305 29009 11339
rect 29043 11336 29055 11339
rect 29362 11336 29368 11348
rect 29043 11308 29368 11336
rect 29043 11305 29055 11308
rect 28997 11299 29055 11305
rect 29012 11268 29040 11299
rect 29362 11296 29368 11308
rect 29420 11296 29426 11348
rect 29914 11336 29920 11348
rect 29472 11308 29920 11336
rect 27816 11240 28120 11268
rect 26559 11172 27108 11200
rect 26559 11169 26571 11172
rect 26513 11163 26571 11169
rect 27522 11160 27528 11212
rect 27580 11200 27586 11212
rect 27816 11209 27844 11240
rect 28092 11209 28120 11240
rect 28460 11240 29040 11268
rect 29181 11271 29239 11277
rect 27801 11203 27859 11209
rect 27801 11200 27813 11203
rect 27580 11172 27813 11200
rect 27580 11160 27586 11172
rect 27801 11169 27813 11172
rect 27847 11169 27859 11203
rect 27801 11163 27859 11169
rect 27985 11203 28043 11209
rect 27985 11169 27997 11203
rect 28031 11169 28043 11203
rect 27985 11163 28043 11169
rect 28077 11203 28135 11209
rect 28077 11169 28089 11203
rect 28123 11169 28135 11203
rect 28077 11163 28135 11169
rect 28261 11203 28319 11209
rect 28261 11169 28273 11203
rect 28307 11190 28319 11203
rect 28460 11198 28488 11240
rect 29181 11237 29193 11271
rect 29227 11268 29239 11271
rect 29472 11268 29500 11308
rect 29914 11296 29920 11308
rect 29972 11296 29978 11348
rect 30098 11296 30104 11348
rect 30156 11296 30162 11348
rect 30285 11339 30343 11345
rect 30285 11305 30297 11339
rect 30331 11336 30343 11339
rect 30926 11336 30932 11348
rect 30331 11308 30932 11336
rect 30331 11305 30343 11308
rect 30285 11299 30343 11305
rect 30116 11268 30144 11296
rect 29227 11240 29500 11268
rect 29664 11240 30144 11268
rect 29227 11237 29239 11240
rect 29181 11231 29239 11237
rect 28368 11190 28488 11198
rect 28307 11170 28488 11190
rect 28537 11203 28595 11209
rect 28307 11169 28396 11170
rect 28261 11163 28396 11169
rect 28537 11169 28549 11203
rect 28583 11200 28595 11203
rect 28626 11200 28632 11212
rect 28583 11172 28632 11200
rect 28583 11169 28595 11172
rect 28537 11163 28595 11169
rect 26881 11135 26939 11141
rect 26881 11132 26893 11135
rect 26160 11104 26893 11132
rect 26881 11101 26893 11104
rect 26927 11132 26939 11135
rect 27154 11132 27160 11144
rect 26927 11104 27160 11132
rect 26927 11101 26939 11104
rect 26881 11095 26939 11101
rect 27154 11092 27160 11104
rect 27212 11092 27218 11144
rect 28000 11132 28028 11163
rect 28276 11162 28396 11163
rect 28626 11160 28632 11172
rect 28684 11160 28690 11212
rect 28721 11203 28779 11209
rect 28721 11169 28733 11203
rect 28767 11200 28779 11203
rect 29196 11200 29224 11231
rect 29664 11210 29692 11240
rect 29656 11209 29692 11210
rect 28767 11172 29224 11200
rect 29457 11203 29515 11209
rect 28767 11169 28779 11172
rect 28721 11163 28779 11169
rect 29457 11169 29469 11203
rect 29503 11169 29515 11203
rect 29457 11163 29515 11169
rect 29641 11203 29699 11209
rect 29641 11169 29653 11203
rect 29687 11169 29699 11203
rect 29641 11163 29699 11169
rect 29733 11203 29791 11209
rect 29733 11169 29745 11203
rect 29779 11169 29791 11203
rect 29733 11163 29791 11169
rect 29917 11203 29975 11209
rect 29917 11169 29929 11203
rect 29963 11200 29975 11203
rect 30300 11200 30328 11299
rect 30926 11296 30932 11308
rect 30984 11296 30990 11348
rect 31110 11296 31116 11348
rect 31168 11336 31174 11348
rect 31205 11339 31263 11345
rect 31205 11336 31217 11339
rect 31168 11308 31217 11336
rect 31168 11296 31174 11308
rect 31205 11305 31217 11308
rect 31251 11336 31263 11339
rect 31846 11336 31852 11348
rect 31251 11308 31852 11336
rect 31251 11305 31263 11308
rect 31205 11299 31263 11305
rect 31846 11296 31852 11308
rect 31904 11296 31910 11348
rect 32582 11336 32588 11348
rect 32324 11308 32588 11336
rect 31754 11268 31760 11280
rect 30392 11240 30696 11268
rect 30392 11209 30420 11240
rect 30668 11212 30696 11240
rect 31680 11240 31760 11268
rect 29963 11172 30328 11200
rect 30377 11203 30435 11209
rect 29963 11169 29975 11172
rect 29917 11163 29975 11169
rect 30377 11169 30389 11203
rect 30423 11169 30435 11203
rect 30377 11163 30435 11169
rect 30561 11203 30619 11209
rect 30561 11169 30573 11203
rect 30607 11169 30619 11203
rect 30561 11163 30619 11169
rect 28445 11135 28503 11141
rect 28445 11132 28457 11135
rect 28000 11104 28457 11132
rect 28445 11101 28457 11104
rect 28491 11132 28503 11135
rect 29086 11132 29092 11144
rect 28491 11104 29092 11132
rect 28491 11101 28503 11104
rect 28445 11095 28503 11101
rect 29086 11092 29092 11104
rect 29144 11092 29150 11144
rect 29472 11132 29500 11163
rect 29748 11132 29776 11163
rect 30392 11132 30420 11163
rect 29472 11104 30420 11132
rect 30576 11132 30604 11163
rect 30650 11160 30656 11212
rect 30708 11160 30714 11212
rect 30834 11160 30840 11212
rect 30892 11160 30898 11212
rect 31680 11209 31708 11240
rect 31754 11228 31760 11240
rect 31812 11228 31818 11280
rect 31481 11203 31539 11209
rect 31481 11169 31493 11203
rect 31527 11169 31539 11203
rect 31481 11163 31539 11169
rect 31665 11203 31723 11209
rect 31665 11169 31677 11203
rect 31711 11169 31723 11203
rect 31665 11163 31723 11169
rect 31021 11135 31079 11141
rect 31021 11132 31033 11135
rect 30576 11104 31033 11132
rect 25593 11067 25651 11073
rect 25593 11033 25605 11067
rect 25639 11064 25651 11067
rect 29178 11064 29184 11076
rect 25639 11036 29184 11064
rect 25639 11033 25651 11036
rect 25593 11027 25651 11033
rect 29178 11024 29184 11036
rect 29236 11024 29242 11076
rect 9122 10956 9128 11008
rect 9180 10996 9186 11008
rect 9490 10996 9496 11008
rect 9180 10968 9496 10996
rect 9180 10956 9186 10968
rect 9490 10956 9496 10968
rect 9548 10956 9554 11008
rect 17126 10956 17132 11008
rect 17184 10996 17190 11008
rect 17494 10996 17500 11008
rect 17184 10968 17500 10996
rect 17184 10956 17190 10968
rect 17494 10956 17500 10968
rect 17552 10956 17558 11008
rect 24210 10956 24216 11008
rect 24268 10956 24274 11008
rect 25222 10956 25228 11008
rect 25280 10996 25286 11008
rect 25961 10999 26019 11005
rect 25961 10996 25973 10999
rect 25280 10968 25973 10996
rect 25280 10956 25286 10968
rect 25961 10965 25973 10968
rect 26007 10965 26019 10999
rect 25961 10959 26019 10965
rect 26418 10956 26424 11008
rect 26476 10956 26482 11008
rect 27890 10956 27896 11008
rect 27948 10956 27954 11008
rect 28166 10956 28172 11008
rect 28224 10956 28230 11008
rect 28626 10956 28632 11008
rect 28684 10956 28690 11008
rect 28718 10956 28724 11008
rect 28776 10996 28782 11008
rect 29472 10996 29500 11104
rect 31021 11101 31033 11104
rect 31067 11132 31079 11135
rect 31496 11132 31524 11163
rect 32030 11160 32036 11212
rect 32088 11200 32094 11212
rect 32324 11209 32352 11308
rect 32582 11296 32588 11308
rect 32640 11296 32646 11348
rect 32766 11296 32772 11348
rect 32824 11336 32830 11348
rect 33689 11339 33747 11345
rect 33689 11336 33701 11339
rect 32824 11308 33701 11336
rect 32824 11296 32830 11308
rect 33689 11305 33701 11308
rect 33735 11336 33747 11339
rect 33778 11336 33784 11348
rect 33735 11308 33784 11336
rect 33735 11305 33747 11308
rect 33689 11299 33747 11305
rect 33778 11296 33784 11308
rect 33836 11296 33842 11348
rect 33870 11296 33876 11348
rect 33928 11296 33934 11348
rect 34149 11339 34207 11345
rect 34149 11305 34161 11339
rect 34195 11336 34207 11339
rect 34330 11336 34336 11348
rect 34195 11308 34336 11336
rect 34195 11305 34207 11308
rect 34149 11299 34207 11305
rect 33888 11268 33916 11296
rect 33068 11240 33916 11268
rect 32309 11203 32367 11209
rect 32309 11200 32321 11203
rect 32088 11172 32321 11200
rect 32088 11160 32094 11172
rect 32309 11169 32321 11172
rect 32355 11169 32367 11203
rect 32484 11201 32542 11207
rect 32484 11200 32496 11201
rect 32309 11163 32367 11169
rect 32416 11172 32496 11200
rect 32048 11132 32076 11160
rect 31067 11104 31340 11132
rect 31496 11104 32076 11132
rect 31067 11101 31079 11104
rect 31021 11095 31079 11101
rect 30745 11067 30803 11073
rect 30745 11033 30757 11067
rect 30791 11064 30803 11067
rect 31312 11064 31340 11104
rect 32214 11092 32220 11144
rect 32272 11132 32278 11144
rect 32416 11132 32444 11172
rect 32484 11167 32496 11172
rect 32530 11167 32542 11201
rect 32484 11161 32542 11167
rect 32582 11160 32588 11212
rect 32640 11160 32646 11212
rect 32766 11160 32772 11212
rect 32824 11160 32830 11212
rect 32858 11160 32864 11212
rect 32916 11198 32922 11212
rect 33068 11209 33096 11240
rect 33045 11203 33103 11209
rect 32916 11170 32996 11198
rect 32916 11160 32922 11170
rect 32272 11104 32444 11132
rect 32968 11132 32996 11170
rect 33045 11169 33057 11203
rect 33091 11169 33103 11203
rect 33045 11163 33103 11169
rect 33137 11203 33195 11209
rect 33137 11169 33149 11203
rect 33183 11169 33195 11203
rect 33137 11163 33195 11169
rect 33321 11203 33379 11209
rect 33321 11169 33333 11203
rect 33367 11200 33379 11203
rect 34164 11200 34192 11299
rect 34330 11296 34336 11308
rect 34388 11296 34394 11348
rect 33367 11172 34192 11200
rect 33367 11169 33379 11172
rect 33321 11163 33379 11169
rect 33158 11132 33186 11163
rect 32968 11104 33186 11132
rect 32272 11092 32278 11104
rect 33502 11092 33508 11144
rect 33560 11092 33566 11144
rect 31478 11064 31484 11076
rect 30791 11036 31248 11064
rect 31312 11036 31484 11064
rect 30791 11033 30803 11036
rect 30745 11027 30803 11033
rect 28776 10968 29500 10996
rect 28776 10956 28782 10968
rect 29546 10956 29552 11008
rect 29604 10956 29610 11008
rect 29822 10956 29828 11008
rect 29880 10956 29886 11008
rect 30466 10956 30472 11008
rect 30524 10956 30530 11008
rect 31220 10996 31248 11036
rect 31478 11024 31484 11036
rect 31536 11024 31542 11076
rect 31573 11067 31631 11073
rect 31573 11033 31585 11067
rect 31619 11064 31631 11067
rect 32401 11067 32459 11073
rect 31619 11036 31984 11064
rect 31619 11033 31631 11036
rect 31573 11027 31631 11033
rect 31956 11008 31984 11036
rect 32401 11033 32413 11067
rect 32447 11064 32459 11067
rect 32953 11067 33011 11073
rect 32447 11036 32904 11064
rect 32447 11033 32459 11036
rect 32401 11027 32459 11033
rect 31846 10996 31852 11008
rect 31220 10968 31852 10996
rect 31846 10956 31852 10968
rect 31904 10956 31910 11008
rect 31938 10956 31944 11008
rect 31996 10956 32002 11008
rect 32677 10999 32735 11005
rect 32677 10965 32689 10999
rect 32723 10996 32735 10999
rect 32766 10996 32772 11008
rect 32723 10968 32772 10996
rect 32723 10965 32735 10968
rect 32677 10959 32735 10965
rect 32766 10956 32772 10968
rect 32824 10956 32830 11008
rect 32876 10996 32904 11036
rect 32953 11033 32965 11067
rect 32999 11064 33011 11067
rect 33686 11064 33692 11076
rect 32999 11036 33692 11064
rect 32999 11033 33011 11036
rect 32953 11027 33011 11033
rect 33686 11024 33692 11036
rect 33744 11024 33750 11076
rect 33134 10996 33140 11008
rect 32876 10968 33140 10996
rect 33134 10956 33140 10968
rect 33192 10956 33198 11008
rect 33229 10999 33287 11005
rect 33229 10965 33241 10999
rect 33275 10996 33287 10999
rect 33778 10996 33784 11008
rect 33275 10968 33784 10996
rect 33275 10965 33287 10968
rect 33229 10959 33287 10965
rect 33778 10956 33784 10968
rect 33836 10956 33842 11008
rect 460 10906 43516 10928
rect 460 10854 1306 10906
rect 1358 10854 1370 10906
rect 1422 10854 1434 10906
rect 1486 10854 1498 10906
rect 1550 10854 1562 10906
rect 1614 10854 9306 10906
rect 9358 10854 9370 10906
rect 9422 10854 9434 10906
rect 9486 10854 9498 10906
rect 9550 10854 9562 10906
rect 9614 10854 17306 10906
rect 17358 10854 17370 10906
rect 17422 10854 17434 10906
rect 17486 10854 17498 10906
rect 17550 10854 17562 10906
rect 17614 10854 25306 10906
rect 25358 10854 25370 10906
rect 25422 10854 25434 10906
rect 25486 10854 25498 10906
rect 25550 10854 25562 10906
rect 25614 10854 33306 10906
rect 33358 10854 33370 10906
rect 33422 10854 33434 10906
rect 33486 10854 33498 10906
rect 33550 10854 33562 10906
rect 33614 10854 41306 10906
rect 41358 10854 41370 10906
rect 41422 10854 41434 10906
rect 41486 10854 41498 10906
rect 41550 10854 41562 10906
rect 41614 10854 43516 10906
rect 460 10832 43516 10854
rect 24673 10795 24731 10801
rect 24673 10761 24685 10795
rect 24719 10792 24731 10795
rect 25774 10792 25780 10804
rect 24719 10764 25780 10792
rect 24719 10761 24731 10764
rect 24673 10755 24731 10761
rect 24302 10548 24308 10600
rect 24360 10548 24366 10600
rect 24489 10591 24547 10597
rect 24489 10557 24501 10591
rect 24535 10588 24547 10591
rect 24688 10588 24716 10755
rect 25774 10752 25780 10764
rect 25832 10752 25838 10804
rect 27893 10795 27951 10801
rect 27893 10761 27905 10795
rect 27939 10792 27951 10795
rect 28810 10792 28816 10804
rect 27939 10764 28816 10792
rect 27939 10761 27951 10764
rect 27893 10755 27951 10761
rect 25409 10727 25467 10733
rect 25409 10693 25421 10727
rect 25455 10724 25467 10727
rect 26326 10724 26332 10736
rect 25455 10696 26332 10724
rect 25455 10693 25467 10696
rect 25409 10687 25467 10693
rect 25424 10656 25452 10687
rect 26326 10684 26332 10696
rect 26384 10684 26390 10736
rect 24964 10628 25452 10656
rect 25593 10659 25651 10665
rect 24964 10597 24992 10628
rect 25593 10625 25605 10659
rect 25639 10656 25651 10659
rect 26602 10656 26608 10668
rect 25639 10628 26608 10656
rect 25639 10625 25651 10628
rect 25593 10619 25651 10625
rect 24535 10560 24716 10588
rect 24765 10591 24823 10597
rect 24535 10557 24547 10560
rect 24489 10551 24547 10557
rect 24765 10557 24777 10591
rect 24811 10557 24823 10591
rect 24765 10551 24823 10557
rect 24949 10591 25007 10597
rect 24949 10557 24961 10591
rect 24995 10557 25007 10591
rect 24949 10551 25007 10557
rect 25041 10591 25099 10597
rect 25041 10557 25053 10591
rect 25087 10557 25099 10591
rect 25041 10551 25099 10557
rect 25225 10591 25283 10597
rect 25225 10557 25237 10591
rect 25271 10588 25283 10591
rect 25608 10588 25636 10619
rect 26602 10616 26608 10628
rect 26660 10616 26666 10668
rect 25271 10560 25636 10588
rect 25271 10557 25283 10560
rect 25225 10551 25283 10557
rect 24320 10520 24348 10548
rect 24780 10520 24808 10551
rect 25056 10520 25084 10551
rect 27154 10548 27160 10600
rect 27212 10588 27218 10600
rect 27522 10588 27528 10600
rect 27212 10560 27528 10588
rect 27212 10548 27218 10560
rect 27522 10548 27528 10560
rect 27580 10548 27586 10600
rect 27709 10591 27767 10597
rect 27709 10557 27721 10591
rect 27755 10588 27767 10591
rect 27908 10588 27936 10755
rect 28810 10752 28816 10764
rect 28868 10752 28874 10804
rect 30466 10752 30472 10804
rect 30524 10792 30530 10804
rect 32214 10792 32220 10804
rect 30524 10764 32220 10792
rect 30524 10752 30530 10764
rect 32214 10752 32220 10764
rect 32272 10752 32278 10804
rect 32309 10795 32367 10801
rect 32309 10761 32321 10795
rect 32355 10792 32367 10795
rect 33226 10792 33232 10804
rect 32355 10764 33232 10792
rect 32355 10761 32367 10764
rect 32309 10755 32367 10761
rect 29546 10684 29552 10736
rect 29604 10724 29610 10736
rect 31202 10724 31208 10736
rect 29604 10696 31208 10724
rect 29604 10684 29610 10696
rect 31202 10684 31208 10696
rect 31260 10684 31266 10736
rect 32030 10656 32036 10668
rect 31956 10628 32036 10656
rect 27755 10560 27936 10588
rect 27755 10557 27767 10560
rect 27709 10551 27767 10557
rect 30650 10548 30656 10600
rect 30708 10588 30714 10600
rect 31662 10588 31668 10600
rect 30708 10560 31668 10588
rect 30708 10548 30714 10560
rect 31662 10548 31668 10560
rect 31720 10588 31726 10600
rect 31956 10597 31984 10628
rect 32030 10616 32036 10628
rect 32088 10616 32094 10668
rect 31941 10591 31999 10597
rect 31941 10588 31953 10591
rect 31720 10560 31953 10588
rect 31720 10548 31726 10560
rect 31941 10557 31953 10560
rect 31987 10557 31999 10591
rect 31941 10551 31999 10557
rect 32125 10591 32183 10597
rect 32125 10557 32137 10591
rect 32171 10588 32183 10591
rect 32324 10588 32352 10755
rect 33226 10752 33232 10764
rect 33284 10752 33290 10804
rect 32171 10560 32352 10588
rect 32171 10557 32183 10560
rect 32125 10551 32183 10557
rect 24320 10492 25084 10520
rect 32033 10523 32091 10529
rect 32033 10489 32045 10523
rect 32079 10520 32091 10523
rect 33042 10520 33048 10532
rect 32079 10492 33048 10520
rect 32079 10489 32091 10492
rect 32033 10483 32091 10489
rect 33042 10480 33048 10492
rect 33100 10480 33106 10532
rect 24486 10412 24492 10464
rect 24544 10412 24550 10464
rect 24854 10412 24860 10464
rect 24912 10412 24918 10464
rect 25130 10412 25136 10464
rect 25188 10412 25194 10464
rect 27706 10412 27712 10464
rect 27764 10412 27770 10464
rect 30006 10412 30012 10464
rect 30064 10452 30070 10464
rect 33226 10452 33232 10464
rect 30064 10424 33232 10452
rect 30064 10412 30070 10424
rect 33226 10412 33232 10424
rect 33284 10412 33290 10464
rect 460 10362 43516 10384
rect 460 10310 1946 10362
rect 1998 10310 2010 10362
rect 2062 10310 2074 10362
rect 2126 10310 2138 10362
rect 2190 10310 2202 10362
rect 2254 10310 9946 10362
rect 9998 10310 10010 10362
rect 10062 10310 10074 10362
rect 10126 10310 10138 10362
rect 10190 10310 10202 10362
rect 10254 10310 17946 10362
rect 17998 10310 18010 10362
rect 18062 10310 18074 10362
rect 18126 10310 18138 10362
rect 18190 10310 18202 10362
rect 18254 10310 25946 10362
rect 25998 10310 26010 10362
rect 26062 10310 26074 10362
rect 26126 10310 26138 10362
rect 26190 10310 26202 10362
rect 26254 10310 33946 10362
rect 33998 10310 34010 10362
rect 34062 10310 34074 10362
rect 34126 10310 34138 10362
rect 34190 10310 34202 10362
rect 34254 10310 41946 10362
rect 41998 10310 42010 10362
rect 42062 10310 42074 10362
rect 42126 10310 42138 10362
rect 42190 10310 42202 10362
rect 42254 10310 43516 10362
rect 460 10288 43516 10310
rect 14734 10208 14740 10260
rect 14792 10208 14798 10260
rect 16666 10208 16672 10260
rect 16724 10208 16730 10260
rect 17218 10208 17224 10260
rect 17276 10248 17282 10260
rect 17313 10251 17371 10257
rect 17313 10248 17325 10251
rect 17276 10220 17325 10248
rect 17276 10208 17282 10220
rect 17313 10217 17325 10220
rect 17359 10217 17371 10251
rect 17313 10211 17371 10217
rect 18046 10208 18052 10260
rect 18104 10248 18110 10260
rect 18233 10251 18291 10257
rect 18233 10248 18245 10251
rect 18104 10220 18245 10248
rect 18104 10208 18110 10220
rect 18233 10217 18245 10220
rect 18279 10248 18291 10251
rect 18690 10248 18696 10260
rect 18279 10220 18696 10248
rect 18279 10217 18291 10220
rect 18233 10211 18291 10217
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 19978 10208 19984 10260
rect 20036 10248 20042 10260
rect 20809 10251 20867 10257
rect 20809 10248 20821 10251
rect 20036 10220 20821 10248
rect 20036 10208 20042 10220
rect 20809 10217 20821 10220
rect 20855 10217 20867 10251
rect 20809 10211 20867 10217
rect 20990 10208 20996 10260
rect 21048 10248 21054 10260
rect 21269 10251 21327 10257
rect 21269 10248 21281 10251
rect 21048 10220 21281 10248
rect 21048 10208 21054 10220
rect 21269 10217 21281 10220
rect 21315 10248 21327 10251
rect 21358 10248 21364 10260
rect 21315 10220 21364 10248
rect 21315 10217 21327 10220
rect 21269 10211 21327 10217
rect 21358 10208 21364 10220
rect 21416 10208 21422 10260
rect 24949 10251 25007 10257
rect 24949 10217 24961 10251
rect 24995 10248 25007 10251
rect 25866 10248 25872 10260
rect 24995 10220 25872 10248
rect 24995 10217 25007 10220
rect 24949 10211 25007 10217
rect 14458 10140 14464 10192
rect 14516 10180 14522 10192
rect 14645 10183 14703 10189
rect 14645 10180 14657 10183
rect 14516 10152 14657 10180
rect 14516 10140 14522 10152
rect 14645 10149 14657 10152
rect 14691 10180 14703 10183
rect 15010 10180 15016 10192
rect 14691 10152 15016 10180
rect 14691 10149 14703 10152
rect 14645 10143 14703 10149
rect 15010 10140 15016 10152
rect 15068 10140 15074 10192
rect 17770 10140 17776 10192
rect 17828 10180 17834 10192
rect 17957 10183 18015 10189
rect 17957 10180 17969 10183
rect 17828 10152 17969 10180
rect 17828 10140 17834 10152
rect 17957 10149 17969 10152
rect 18003 10180 18015 10183
rect 18598 10180 18604 10192
rect 18003 10152 18604 10180
rect 18003 10149 18015 10152
rect 17957 10143 18015 10149
rect 18598 10140 18604 10152
rect 18656 10140 18662 10192
rect 19794 10140 19800 10192
rect 19852 10180 19858 10192
rect 19889 10183 19947 10189
rect 19889 10180 19901 10183
rect 19852 10152 19901 10180
rect 19852 10140 19858 10152
rect 19889 10149 19901 10152
rect 19935 10180 19947 10183
rect 20438 10180 20444 10192
rect 19935 10152 20444 10180
rect 19935 10149 19947 10152
rect 19889 10143 19947 10149
rect 20438 10140 20444 10152
rect 20496 10140 20502 10192
rect 13446 10072 13452 10124
rect 13504 10112 13510 10124
rect 18782 10112 18788 10124
rect 13504 10084 18788 10112
rect 13504 10072 13510 10084
rect 18782 10072 18788 10084
rect 18840 10072 18846 10124
rect 20346 10072 20352 10124
rect 20404 10112 20410 10124
rect 20533 10115 20591 10121
rect 20533 10112 20545 10115
rect 20404 10084 20545 10112
rect 20404 10072 20410 10084
rect 20533 10081 20545 10084
rect 20579 10112 20591 10115
rect 20806 10112 20812 10124
rect 20579 10084 20812 10112
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 20806 10072 20812 10084
rect 20864 10072 20870 10124
rect 24302 10072 24308 10124
rect 24360 10112 24366 10124
rect 24581 10115 24639 10121
rect 24581 10112 24593 10115
rect 24360 10084 24593 10112
rect 24360 10072 24366 10084
rect 24581 10081 24593 10084
rect 24627 10081 24639 10115
rect 24581 10075 24639 10081
rect 24765 10115 24823 10121
rect 24765 10081 24777 10115
rect 24811 10112 24823 10115
rect 24964 10112 24992 10211
rect 25866 10208 25872 10220
rect 25924 10208 25930 10260
rect 27801 10251 27859 10257
rect 27801 10217 27813 10251
rect 27847 10248 27859 10251
rect 27982 10248 27988 10260
rect 27847 10220 27988 10248
rect 27847 10217 27859 10220
rect 27801 10211 27859 10217
rect 27816 10180 27844 10211
rect 27982 10208 27988 10220
rect 28040 10208 28046 10260
rect 28169 10251 28227 10257
rect 28169 10217 28181 10251
rect 28215 10248 28227 10251
rect 28534 10248 28540 10260
rect 28215 10220 28540 10248
rect 28215 10217 28227 10220
rect 28169 10211 28227 10217
rect 27080 10152 27844 10180
rect 24811 10084 24992 10112
rect 24811 10081 24823 10084
rect 24765 10075 24823 10081
rect 26326 10072 26332 10124
rect 26384 10112 26390 10124
rect 27080 10121 27108 10152
rect 26881 10115 26939 10121
rect 26881 10112 26893 10115
rect 26384 10084 26893 10112
rect 26384 10072 26390 10084
rect 26881 10081 26893 10084
rect 26927 10081 26939 10115
rect 26881 10075 26939 10081
rect 27065 10115 27123 10121
rect 27065 10081 27077 10115
rect 27111 10081 27123 10115
rect 27065 10075 27123 10081
rect 15654 10004 15660 10056
rect 15712 10044 15718 10056
rect 18230 10044 18236 10056
rect 15712 10016 18236 10044
rect 15712 10004 15718 10016
rect 18230 10004 18236 10016
rect 18288 10004 18294 10056
rect 26896 10044 26924 10075
rect 27154 10072 27160 10124
rect 27212 10072 27218 10124
rect 27338 10072 27344 10124
rect 27396 10072 27402 10124
rect 27456 10115 27514 10121
rect 27456 10081 27468 10115
rect 27502 10081 27514 10115
rect 27456 10075 27514 10081
rect 27617 10115 27675 10121
rect 27617 10081 27629 10115
rect 27663 10112 27675 10115
rect 28184 10112 28212 10211
rect 28534 10208 28540 10220
rect 28592 10208 28598 10260
rect 29932 10220 30696 10248
rect 29932 10180 29960 10220
rect 29012 10152 29960 10180
rect 29012 10122 29040 10152
rect 27663 10084 28212 10112
rect 28828 10105 29040 10122
rect 29196 10121 29224 10152
rect 29932 10121 29960 10152
rect 30006 10140 30012 10192
rect 30064 10140 30070 10192
rect 30668 10180 30696 10220
rect 30834 10208 30840 10260
rect 30892 10248 30898 10260
rect 31297 10251 31355 10257
rect 31297 10248 31309 10251
rect 30892 10220 31309 10248
rect 30892 10208 30898 10220
rect 31297 10217 31309 10220
rect 31343 10248 31355 10251
rect 31386 10248 31392 10260
rect 31343 10220 31392 10248
rect 31343 10217 31355 10220
rect 31297 10211 31355 10217
rect 31386 10208 31392 10220
rect 31444 10208 31450 10260
rect 32033 10251 32091 10257
rect 32033 10217 32045 10251
rect 32079 10248 32091 10251
rect 32950 10248 32956 10260
rect 32079 10220 32956 10248
rect 32079 10217 32091 10220
rect 32033 10211 32091 10217
rect 31021 10183 31079 10189
rect 30668 10152 30972 10180
rect 30668 10121 30696 10152
rect 27663 10081 27675 10084
rect 27617 10075 27675 10081
rect 27172 10044 27200 10072
rect 27471 10044 27499 10075
rect 28828 10074 28917 10105
rect 26896 10016 27499 10044
rect 27985 10047 28043 10053
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 17497 9979 17555 9985
rect 17497 9976 17509 9979
rect 16632 9948 17509 9976
rect 16632 9936 16638 9948
rect 17497 9945 17509 9948
rect 17543 9945 17555 9979
rect 17497 9939 17555 9945
rect 20349 9979 20407 9985
rect 20349 9945 20361 9979
rect 20395 9976 20407 9979
rect 20530 9976 20536 9988
rect 20395 9948 20536 9976
rect 20395 9945 20407 9948
rect 20349 9939 20407 9945
rect 20530 9936 20536 9948
rect 20588 9936 20594 9988
rect 27448 9976 27476 10016
rect 27985 10013 27997 10047
rect 28031 10044 28043 10047
rect 28258 10044 28264 10056
rect 28031 10016 28264 10044
rect 28031 10013 28043 10016
rect 27985 10007 28043 10013
rect 28258 10004 28264 10016
rect 28316 10004 28322 10056
rect 28828 10044 28856 10074
rect 28905 10071 28917 10074
rect 28951 10094 29040 10105
rect 29089 10115 29147 10121
rect 28951 10071 28963 10094
rect 29089 10081 29101 10115
rect 29135 10081 29147 10115
rect 29089 10075 29147 10081
rect 29181 10115 29239 10121
rect 29181 10081 29193 10115
rect 29227 10081 29239 10115
rect 29181 10075 29239 10081
rect 29365 10115 29423 10121
rect 29365 10081 29377 10115
rect 29411 10110 29423 10115
rect 29917 10115 29975 10121
rect 29411 10082 29500 10110
rect 29411 10081 29423 10082
rect 29365 10075 29423 10081
rect 28905 10065 28963 10071
rect 28460 10016 28856 10044
rect 28074 9976 28080 9988
rect 27448 9948 28080 9976
rect 28074 9936 28080 9948
rect 28132 9976 28138 9988
rect 28460 9976 28488 10016
rect 28132 9948 28488 9976
rect 29104 9976 29132 10075
rect 29472 9976 29500 10082
rect 29917 10081 29929 10115
rect 29963 10081 29975 10115
rect 29917 10075 29975 10081
rect 30101 10115 30159 10121
rect 30101 10081 30113 10115
rect 30147 10112 30159 10115
rect 30653 10115 30711 10121
rect 30147 10084 30328 10112
rect 30147 10081 30159 10084
rect 30101 10075 30159 10081
rect 29546 10004 29552 10056
rect 29604 10044 29610 10056
rect 30190 10044 30196 10056
rect 29604 10016 30196 10044
rect 29604 10004 29610 10016
rect 30190 10004 30196 10016
rect 30248 10004 30254 10056
rect 30300 9985 30328 10084
rect 30653 10081 30665 10115
rect 30699 10081 30711 10115
rect 30653 10075 30711 10081
rect 30834 10072 30840 10124
rect 30892 10072 30898 10124
rect 30944 10121 30972 10152
rect 31021 10149 31033 10183
rect 31067 10180 31079 10183
rect 32122 10180 32128 10192
rect 31067 10152 32128 10180
rect 31067 10149 31079 10152
rect 31021 10143 31079 10149
rect 32122 10140 32128 10152
rect 32180 10140 32186 10192
rect 30929 10115 30987 10121
rect 30929 10081 30941 10115
rect 30975 10081 30987 10115
rect 30929 10075 30987 10081
rect 31110 10072 31116 10124
rect 31168 10072 31174 10124
rect 31662 10072 31668 10124
rect 31720 10072 31726 10124
rect 31849 10115 31907 10121
rect 31849 10081 31861 10115
rect 31895 10112 31907 10115
rect 32416 10112 32444 10220
rect 32950 10208 32956 10220
rect 33008 10208 33014 10260
rect 31895 10084 32444 10112
rect 31895 10081 31907 10084
rect 31849 10075 31907 10081
rect 30285 9979 30343 9985
rect 29104 9948 29408 9976
rect 29472 9948 29776 9976
rect 28132 9936 28138 9948
rect 13909 9911 13967 9917
rect 13909 9877 13921 9911
rect 13955 9908 13967 9911
rect 14090 9908 14096 9920
rect 13955 9880 14096 9908
rect 13955 9877 13967 9880
rect 13909 9871 13967 9877
rect 14090 9868 14096 9880
rect 14148 9868 14154 9920
rect 14461 9911 14519 9917
rect 14461 9877 14473 9911
rect 14507 9908 14519 9911
rect 14642 9908 14648 9920
rect 14507 9880 14648 9908
rect 14507 9877 14519 9880
rect 14461 9871 14519 9877
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16206 9908 16212 9920
rect 16163 9880 16212 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16206 9868 16212 9880
rect 16264 9868 16270 9920
rect 16298 9868 16304 9920
rect 16356 9908 16362 9920
rect 16393 9911 16451 9917
rect 16393 9908 16405 9911
rect 16356 9880 16405 9908
rect 16356 9868 16362 9880
rect 16393 9877 16405 9880
rect 16439 9877 16451 9911
rect 16393 9871 16451 9877
rect 16850 9868 16856 9920
rect 16908 9868 16914 9920
rect 17034 9868 17040 9920
rect 17092 9868 17098 9920
rect 17773 9911 17831 9917
rect 17773 9877 17785 9911
rect 17819 9908 17831 9911
rect 17862 9908 17868 9920
rect 17819 9880 17868 9908
rect 17819 9877 17831 9880
rect 17773 9871 17831 9877
rect 17862 9868 17868 9880
rect 17920 9868 17926 9920
rect 19061 9911 19119 9917
rect 19061 9877 19073 9911
rect 19107 9908 19119 9911
rect 19242 9908 19248 9920
rect 19107 9880 19248 9908
rect 19107 9877 19119 9880
rect 19061 9871 19119 9877
rect 19242 9868 19248 9880
rect 19300 9868 19306 9920
rect 19429 9911 19487 9917
rect 19429 9877 19441 9911
rect 19475 9908 19487 9911
rect 19610 9908 19616 9920
rect 19475 9880 19616 9908
rect 19475 9877 19487 9880
rect 19429 9871 19487 9877
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 19705 9911 19763 9917
rect 19705 9877 19717 9911
rect 19751 9908 19763 9911
rect 19886 9908 19892 9920
rect 19751 9880 19892 9908
rect 19751 9877 19763 9880
rect 19705 9871 19763 9877
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 20714 9868 20720 9920
rect 20772 9868 20778 9920
rect 24670 9868 24676 9920
rect 24728 9868 24734 9920
rect 26970 9868 26976 9920
rect 27028 9868 27034 9920
rect 27246 9868 27252 9920
rect 27304 9868 27310 9920
rect 27525 9911 27583 9917
rect 27525 9877 27537 9911
rect 27571 9908 27583 9911
rect 27614 9908 27620 9920
rect 27571 9880 27620 9908
rect 27571 9877 27583 9880
rect 27525 9871 27583 9877
rect 27614 9868 27620 9880
rect 27672 9868 27678 9920
rect 28994 9868 29000 9920
rect 29052 9868 29058 9920
rect 29270 9868 29276 9920
rect 29328 9868 29334 9920
rect 29380 9908 29408 9948
rect 29546 9908 29552 9920
rect 29380 9880 29552 9908
rect 29546 9868 29552 9880
rect 29604 9868 29610 9920
rect 29748 9917 29776 9948
rect 30285 9945 30297 9979
rect 30331 9976 30343 9979
rect 31294 9976 31300 9988
rect 30331 9948 31300 9976
rect 30331 9945 30343 9948
rect 30285 9939 30343 9945
rect 31294 9936 31300 9948
rect 31352 9936 31358 9988
rect 31757 9979 31815 9985
rect 31757 9945 31769 9979
rect 31803 9976 31815 9979
rect 32674 9976 32680 9988
rect 31803 9948 32680 9976
rect 31803 9945 31815 9948
rect 31757 9939 31815 9945
rect 32674 9936 32680 9948
rect 32732 9936 32738 9988
rect 29733 9911 29791 9917
rect 29733 9877 29745 9911
rect 29779 9908 29791 9911
rect 30374 9908 30380 9920
rect 29779 9880 30380 9908
rect 29779 9877 29791 9880
rect 29733 9871 29791 9877
rect 30374 9868 30380 9880
rect 30432 9868 30438 9920
rect 30742 9868 30748 9920
rect 30800 9868 30806 9920
rect 31110 9868 31116 9920
rect 31168 9908 31174 9920
rect 31573 9911 31631 9917
rect 31573 9908 31585 9911
rect 31168 9880 31585 9908
rect 31168 9868 31174 9880
rect 31573 9877 31585 9880
rect 31619 9908 31631 9911
rect 32398 9908 32404 9920
rect 31619 9880 32404 9908
rect 31619 9877 31631 9880
rect 31573 9871 31631 9877
rect 32398 9868 32404 9880
rect 32456 9868 32462 9920
rect 460 9818 43516 9840
rect 460 9766 1306 9818
rect 1358 9766 1370 9818
rect 1422 9766 1434 9818
rect 1486 9766 1498 9818
rect 1550 9766 1562 9818
rect 1614 9766 9306 9818
rect 9358 9766 9370 9818
rect 9422 9766 9434 9818
rect 9486 9766 9498 9818
rect 9550 9766 9562 9818
rect 9614 9766 17306 9818
rect 17358 9766 17370 9818
rect 17422 9766 17434 9818
rect 17486 9766 17498 9818
rect 17550 9766 17562 9818
rect 17614 9766 25306 9818
rect 25358 9766 25370 9818
rect 25422 9766 25434 9818
rect 25486 9766 25498 9818
rect 25550 9766 25562 9818
rect 25614 9766 33306 9818
rect 33358 9766 33370 9818
rect 33422 9766 33434 9818
rect 33486 9766 33498 9818
rect 33550 9766 33562 9818
rect 33614 9766 41306 9818
rect 41358 9766 41370 9818
rect 41422 9766 41434 9818
rect 41486 9766 41498 9818
rect 41550 9766 41562 9818
rect 41614 9766 43516 9818
rect 460 9744 43516 9766
rect 14366 9704 14372 9716
rect 13832 9676 14372 9704
rect 12986 9596 12992 9648
rect 13044 9636 13050 9648
rect 13173 9639 13231 9645
rect 13173 9636 13185 9639
rect 13044 9608 13185 9636
rect 13044 9596 13050 9608
rect 13173 9605 13185 9608
rect 13219 9636 13231 9639
rect 13630 9636 13636 9648
rect 13219 9608 13636 9636
rect 13219 9605 13231 9608
rect 13173 9599 13231 9605
rect 13630 9596 13636 9608
rect 13688 9596 13694 9648
rect 13832 9580 13860 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 16301 9707 16359 9713
rect 14936 9676 15700 9704
rect 14936 9636 14964 9676
rect 13924 9608 14964 9636
rect 15013 9639 15071 9645
rect 11054 9528 11060 9580
rect 11112 9568 11118 9580
rect 13446 9568 13452 9580
rect 11112 9540 13452 9568
rect 11112 9528 11118 9540
rect 13446 9528 13452 9540
rect 13504 9528 13510 9580
rect 13541 9571 13599 9577
rect 13541 9537 13553 9571
rect 13587 9568 13599 9571
rect 13814 9568 13820 9580
rect 13587 9540 13820 9568
rect 13587 9537 13599 9540
rect 13541 9531 13599 9537
rect 13814 9528 13820 9540
rect 13872 9528 13878 9580
rect 8754 9460 8760 9512
rect 8812 9500 8818 9512
rect 13924 9500 13952 9608
rect 15013 9605 15025 9639
rect 15059 9636 15071 9639
rect 15562 9636 15568 9648
rect 15059 9608 15568 9636
rect 15059 9605 15071 9608
rect 15013 9599 15071 9605
rect 15562 9596 15568 9608
rect 15620 9596 15626 9648
rect 15672 9636 15700 9676
rect 16301 9673 16313 9707
rect 16347 9704 16359 9707
rect 16666 9704 16672 9716
rect 16347 9676 16672 9704
rect 16347 9673 16359 9676
rect 16301 9667 16359 9673
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 16945 9707 17003 9713
rect 16945 9673 16957 9707
rect 16991 9704 17003 9707
rect 17218 9704 17224 9716
rect 16991 9676 17224 9704
rect 16991 9673 17003 9676
rect 16945 9667 17003 9673
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17586 9664 17592 9716
rect 17644 9704 17650 9716
rect 17862 9704 17868 9716
rect 17644 9676 17868 9704
rect 17644 9664 17650 9676
rect 17862 9664 17868 9676
rect 17920 9664 17926 9716
rect 21542 9704 21548 9716
rect 19628 9676 21548 9704
rect 15746 9636 15752 9648
rect 15672 9608 15752 9636
rect 15746 9596 15752 9608
rect 15804 9596 15810 9648
rect 15933 9639 15991 9645
rect 15933 9605 15945 9639
rect 15979 9636 15991 9639
rect 16114 9636 16120 9648
rect 15979 9608 16120 9636
rect 15979 9605 15991 9608
rect 15933 9599 15991 9605
rect 16114 9596 16120 9608
rect 16172 9596 16178 9648
rect 16500 9608 18368 9636
rect 14001 9571 14059 9577
rect 14001 9537 14013 9571
rect 14047 9568 14059 9571
rect 14274 9568 14280 9580
rect 14047 9540 14280 9568
rect 14047 9537 14059 9540
rect 14001 9531 14059 9537
rect 14274 9528 14280 9540
rect 14332 9528 14338 9580
rect 14553 9571 14611 9577
rect 14553 9537 14565 9571
rect 14599 9568 14611 9571
rect 14734 9568 14740 9580
rect 14599 9540 14740 9568
rect 14599 9537 14611 9540
rect 14553 9531 14611 9537
rect 14734 9528 14740 9540
rect 14792 9528 14798 9580
rect 15194 9528 15200 9580
rect 15252 9568 15258 9580
rect 15381 9571 15439 9577
rect 15381 9568 15393 9571
rect 15252 9540 15393 9568
rect 15252 9528 15258 9540
rect 15381 9537 15393 9540
rect 15427 9568 15439 9571
rect 15838 9568 15844 9580
rect 15427 9540 15844 9568
rect 15427 9537 15439 9540
rect 15381 9531 15439 9537
rect 15838 9528 15844 9540
rect 15896 9528 15902 9580
rect 16500 9568 16528 9608
rect 15948 9540 16528 9568
rect 8812 9472 13952 9500
rect 8812 9460 8818 9472
rect 14090 9460 14096 9512
rect 14148 9460 14154 9512
rect 15948 9500 15976 9540
rect 16574 9528 16580 9580
rect 16632 9568 16638 9580
rect 16632 9540 17632 9568
rect 16632 9528 16638 9540
rect 14660 9472 15976 9500
rect 13262 9392 13268 9444
rect 13320 9432 13326 9444
rect 14660 9432 14688 9472
rect 16022 9460 16028 9512
rect 16080 9460 16086 9512
rect 16117 9503 16175 9509
rect 16117 9469 16129 9503
rect 16163 9500 16175 9503
rect 16206 9500 16212 9512
rect 16163 9472 16212 9500
rect 16163 9469 16175 9472
rect 16117 9463 16175 9469
rect 16206 9460 16212 9472
rect 16264 9460 16270 9512
rect 16666 9460 16672 9512
rect 16724 9500 16730 9512
rect 16850 9500 16856 9512
rect 16724 9472 16856 9500
rect 16724 9460 16730 9472
rect 16850 9460 16856 9472
rect 16908 9500 16914 9512
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 16908 9472 17141 9500
rect 16908 9460 16914 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 17221 9503 17279 9509
rect 17221 9469 17233 9503
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 13320 9404 14688 9432
rect 13320 9392 13326 9404
rect 14734 9392 14740 9444
rect 14792 9432 14798 9444
rect 15470 9432 15476 9444
rect 14792 9404 15476 9432
rect 14792 9392 14798 9404
rect 15470 9392 15476 9404
rect 15528 9392 15534 9444
rect 15565 9435 15623 9441
rect 15565 9401 15577 9435
rect 15611 9432 15623 9435
rect 16942 9432 16948 9444
rect 15611 9404 16948 9432
rect 15611 9401 15623 9404
rect 15565 9395 15623 9401
rect 16942 9392 16948 9404
rect 17000 9392 17006 9444
rect 17236 9432 17264 9463
rect 17494 9460 17500 9512
rect 17552 9460 17558 9512
rect 17604 9509 17632 9540
rect 18046 9528 18052 9580
rect 18104 9528 18110 9580
rect 18340 9568 18368 9608
rect 18414 9596 18420 9648
rect 18472 9636 18478 9648
rect 18874 9636 18880 9648
rect 18472 9608 18880 9636
rect 18472 9596 18478 9608
rect 18874 9596 18880 9608
rect 18932 9596 18938 9648
rect 19150 9596 19156 9648
rect 19208 9596 19214 9648
rect 19628 9636 19656 9676
rect 21542 9664 21548 9676
rect 21600 9664 21606 9716
rect 22112 9676 24440 9704
rect 19444 9608 19656 9636
rect 18690 9568 18696 9580
rect 18340 9540 18696 9568
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 19444 9568 19472 9608
rect 19702 9596 19708 9648
rect 19760 9636 19766 9648
rect 20165 9639 20223 9645
rect 20165 9636 20177 9639
rect 19760 9608 20177 9636
rect 19760 9596 19766 9608
rect 20165 9605 20177 9608
rect 20211 9605 20223 9639
rect 22112 9636 22140 9676
rect 20165 9599 20223 9605
rect 20640 9608 22140 9636
rect 18800 9540 19472 9568
rect 19521 9571 19579 9577
rect 17589 9503 17647 9509
rect 17589 9469 17601 9503
rect 17635 9469 17647 9503
rect 18800 9500 18828 9540
rect 19521 9537 19533 9571
rect 19567 9568 19579 9571
rect 19567 9540 19932 9568
rect 19567 9537 19579 9540
rect 19521 9531 19579 9537
rect 17589 9463 17647 9469
rect 18340 9472 18828 9500
rect 18877 9503 18935 9509
rect 18340 9432 18368 9472
rect 18877 9469 18889 9503
rect 18923 9500 18935 9503
rect 18966 9500 18972 9512
rect 18923 9472 18972 9500
rect 18923 9469 18935 9472
rect 18877 9463 18935 9469
rect 18966 9460 18972 9472
rect 19024 9500 19030 9512
rect 19426 9500 19432 9512
rect 19024 9472 19432 9500
rect 19024 9460 19030 9472
rect 19426 9460 19432 9472
rect 19484 9460 19490 9512
rect 19610 9460 19616 9512
rect 19668 9460 19674 9512
rect 19904 9500 19932 9540
rect 19978 9528 19984 9580
rect 20036 9568 20042 9580
rect 20640 9577 20668 9608
rect 22186 9596 22192 9648
rect 22244 9636 22250 9648
rect 22649 9639 22707 9645
rect 22649 9636 22661 9639
rect 22244 9608 22661 9636
rect 22244 9596 22250 9608
rect 22649 9605 22661 9608
rect 22695 9605 22707 9639
rect 22649 9599 22707 9605
rect 22738 9596 22744 9648
rect 22796 9636 22802 9648
rect 23201 9639 23259 9645
rect 23201 9636 23213 9639
rect 22796 9608 23213 9636
rect 22796 9596 22802 9608
rect 23201 9605 23213 9608
rect 23247 9605 23259 9639
rect 23201 9599 23259 9605
rect 23566 9596 23572 9648
rect 23624 9636 23630 9648
rect 24305 9639 24363 9645
rect 24305 9636 24317 9639
rect 23624 9608 24317 9636
rect 23624 9596 23630 9608
rect 24305 9605 24317 9608
rect 24351 9605 24363 9639
rect 24412 9636 24440 9676
rect 32858 9664 32864 9716
rect 32916 9704 32922 9716
rect 33318 9704 33324 9716
rect 32916 9676 33324 9704
rect 32916 9664 32922 9676
rect 33318 9664 33324 9676
rect 33376 9664 33382 9716
rect 38746 9664 38752 9716
rect 38804 9704 38810 9716
rect 40494 9704 40500 9716
rect 38804 9676 40500 9704
rect 38804 9664 38810 9676
rect 40494 9664 40500 9676
rect 40552 9664 40558 9716
rect 24486 9636 24492 9648
rect 24412 9608 24492 9636
rect 24305 9599 24363 9605
rect 24486 9596 24492 9608
rect 24544 9596 24550 9648
rect 24762 9596 24768 9648
rect 24820 9636 24826 9648
rect 25501 9639 25559 9645
rect 25501 9636 25513 9639
rect 24820 9608 25513 9636
rect 24820 9596 24826 9608
rect 25501 9605 25513 9608
rect 25547 9605 25559 9639
rect 25501 9599 25559 9605
rect 28537 9639 28595 9645
rect 28537 9605 28549 9639
rect 28583 9636 28595 9639
rect 29638 9636 29644 9648
rect 28583 9608 29644 9636
rect 28583 9605 28595 9608
rect 28537 9599 28595 9605
rect 20073 9571 20131 9577
rect 20073 9568 20085 9571
rect 20036 9540 20085 9568
rect 20036 9528 20042 9540
rect 20073 9537 20085 9540
rect 20119 9537 20131 9571
rect 20073 9531 20131 9537
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9537 20683 9571
rect 20625 9531 20683 9537
rect 21082 9528 21088 9580
rect 21140 9568 21146 9580
rect 21177 9571 21235 9577
rect 21177 9568 21189 9571
rect 21140 9540 21189 9568
rect 21140 9528 21146 9540
rect 21177 9537 21189 9540
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 19904 9472 20668 9500
rect 17236 9404 18368 9432
rect 18690 9392 18696 9444
rect 18748 9432 18754 9444
rect 20070 9432 20076 9444
rect 18748 9404 20076 9432
rect 18748 9392 18754 9404
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 20162 9392 20168 9444
rect 20220 9432 20226 9444
rect 20640 9432 20668 9472
rect 20714 9460 20720 9512
rect 20772 9460 20778 9512
rect 21192 9500 21220 9531
rect 21358 9528 21364 9580
rect 21416 9528 21422 9580
rect 21634 9528 21640 9580
rect 21692 9568 21698 9580
rect 21913 9571 21971 9577
rect 21913 9568 21925 9571
rect 21692 9540 21925 9568
rect 21692 9528 21698 9540
rect 21913 9537 21925 9540
rect 21959 9537 21971 9571
rect 22922 9568 22928 9580
rect 21913 9531 21971 9537
rect 22296 9540 22928 9568
rect 22097 9503 22155 9509
rect 22097 9500 22109 9503
rect 21192 9472 22109 9500
rect 22097 9469 22109 9472
rect 22143 9469 22155 9503
rect 22097 9463 22155 9469
rect 20806 9432 20812 9444
rect 20220 9404 20576 9432
rect 20640 9404 20812 9432
rect 20220 9392 20226 9404
rect 12710 9324 12716 9376
rect 12768 9364 12774 9376
rect 13630 9364 13636 9376
rect 12768 9336 13636 9364
rect 12768 9324 12774 9336
rect 13630 9324 13636 9336
rect 13688 9364 13694 9376
rect 13817 9367 13875 9373
rect 13817 9364 13829 9367
rect 13688 9336 13829 9364
rect 13688 9324 13694 9336
rect 13817 9333 13829 9336
rect 13863 9333 13875 9367
rect 13817 9327 13875 9333
rect 15197 9367 15255 9373
rect 15197 9333 15209 9367
rect 15243 9364 15255 9367
rect 15378 9364 15384 9376
rect 15243 9336 15384 9364
rect 15243 9333 15255 9336
rect 15197 9327 15255 9333
rect 15378 9324 15384 9336
rect 15436 9324 15442 9376
rect 15749 9367 15807 9373
rect 15749 9333 15761 9367
rect 15795 9364 15807 9367
rect 15838 9364 15844 9376
rect 15795 9336 15844 9364
rect 15795 9333 15807 9336
rect 15749 9327 15807 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 17405 9367 17463 9373
rect 17405 9333 17417 9367
rect 17451 9364 17463 9367
rect 17862 9364 17868 9376
rect 17451 9336 17868 9364
rect 17451 9333 17463 9336
rect 17405 9327 17463 9333
rect 17862 9324 17868 9336
rect 17920 9324 17926 9376
rect 18138 9324 18144 9376
rect 18196 9324 18202 9376
rect 18598 9324 18604 9376
rect 18656 9324 18662 9376
rect 19061 9367 19119 9373
rect 19061 9333 19073 9367
rect 19107 9364 19119 9367
rect 19334 9364 19340 9376
rect 19107 9336 19340 9364
rect 19107 9333 19119 9336
rect 19061 9327 19119 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 19429 9367 19487 9373
rect 19429 9333 19441 9367
rect 19475 9364 19487 9367
rect 19518 9364 19524 9376
rect 19475 9336 19524 9364
rect 19475 9333 19487 9336
rect 19429 9327 19487 9333
rect 19518 9324 19524 9336
rect 19576 9324 19582 9376
rect 19978 9324 19984 9376
rect 20036 9364 20042 9376
rect 20441 9367 20499 9373
rect 20441 9364 20453 9367
rect 20036 9336 20453 9364
rect 20036 9324 20042 9336
rect 20441 9333 20453 9336
rect 20487 9333 20499 9367
rect 20548 9364 20576 9404
rect 20806 9392 20812 9404
rect 20864 9392 20870 9444
rect 20898 9392 20904 9444
rect 20956 9432 20962 9444
rect 22296 9432 22324 9540
rect 22922 9528 22928 9540
rect 22980 9528 22986 9580
rect 23014 9528 23020 9580
rect 23072 9568 23078 9580
rect 23937 9571 23995 9577
rect 23937 9568 23949 9571
rect 23072 9540 23949 9568
rect 23072 9528 23078 9540
rect 23937 9537 23949 9540
rect 23983 9537 23995 9571
rect 23937 9531 23995 9537
rect 24026 9528 24032 9580
rect 24084 9568 24090 9580
rect 24581 9571 24639 9577
rect 24581 9568 24593 9571
rect 24084 9540 24593 9568
rect 24084 9528 24090 9540
rect 24581 9537 24593 9540
rect 24627 9537 24639 9571
rect 24581 9531 24639 9537
rect 23845 9503 23903 9509
rect 23845 9469 23857 9503
rect 23891 9500 23903 9503
rect 24118 9500 24124 9512
rect 23891 9472 24124 9500
rect 23891 9469 23903 9472
rect 23845 9463 23903 9469
rect 24118 9460 24124 9472
rect 24176 9460 24182 9512
rect 28074 9460 28080 9512
rect 28132 9500 28138 9512
rect 28169 9503 28227 9509
rect 28169 9500 28181 9503
rect 28132 9472 28181 9500
rect 28132 9460 28138 9472
rect 28169 9469 28181 9472
rect 28215 9469 28227 9503
rect 28169 9463 28227 9469
rect 28353 9503 28411 9509
rect 28353 9469 28365 9503
rect 28399 9500 28411 9503
rect 28552 9500 28580 9599
rect 29638 9596 29644 9608
rect 29696 9596 29702 9648
rect 28399 9472 28580 9500
rect 28399 9469 28411 9472
rect 28353 9463 28411 9469
rect 20956 9404 22324 9432
rect 20956 9392 20962 9404
rect 22554 9392 22560 9444
rect 22612 9392 22618 9444
rect 25406 9392 25412 9444
rect 25464 9392 25470 9444
rect 21453 9367 21511 9373
rect 21453 9364 21465 9367
rect 20548 9336 21465 9364
rect 20441 9327 20499 9333
rect 21453 9333 21465 9336
rect 21499 9333 21511 9367
rect 21453 9327 21511 9333
rect 21726 9324 21732 9376
rect 21784 9324 21790 9376
rect 23477 9367 23535 9373
rect 23477 9333 23489 9367
rect 23523 9364 23535 9367
rect 23750 9364 23756 9376
rect 23523 9336 23756 9364
rect 23523 9333 23535 9336
rect 23477 9327 23535 9333
rect 23750 9324 23756 9336
rect 23808 9324 23814 9376
rect 23842 9324 23848 9376
rect 23900 9364 23906 9376
rect 24121 9367 24179 9373
rect 24121 9364 24133 9367
rect 23900 9336 24133 9364
rect 23900 9324 23906 9336
rect 24121 9333 24133 9336
rect 24167 9333 24179 9367
rect 24121 9327 24179 9333
rect 24670 9324 24676 9376
rect 24728 9364 24734 9376
rect 24765 9367 24823 9373
rect 24765 9364 24777 9367
rect 24728 9336 24777 9364
rect 24728 9324 24734 9336
rect 24765 9333 24777 9336
rect 24811 9333 24823 9367
rect 24765 9327 24823 9333
rect 28350 9324 28356 9376
rect 28408 9324 28414 9376
rect 460 9274 43516 9296
rect 460 9222 1946 9274
rect 1998 9222 2010 9274
rect 2062 9222 2074 9274
rect 2126 9222 2138 9274
rect 2190 9222 2202 9274
rect 2254 9222 9946 9274
rect 9998 9222 10010 9274
rect 10062 9222 10074 9274
rect 10126 9222 10138 9274
rect 10190 9222 10202 9274
rect 10254 9222 33946 9274
rect 33998 9222 34010 9274
rect 34062 9222 34074 9274
rect 34126 9222 34138 9274
rect 34190 9222 34202 9274
rect 34254 9222 41946 9274
rect 41998 9222 42010 9274
rect 42062 9222 42074 9274
rect 42126 9222 42138 9274
rect 42190 9222 42202 9274
rect 42254 9222 43516 9274
rect 460 9200 43516 9222
rect 11609 9163 11667 9169
rect 11609 9160 11621 9163
rect 11440 9132 11621 9160
rect 10134 9052 10140 9104
rect 10192 9092 10198 9104
rect 11440 9101 11468 9132
rect 11609 9129 11621 9132
rect 11655 9160 11667 9163
rect 12250 9160 12256 9172
rect 11655 9132 12256 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 12250 9120 12256 9132
rect 12308 9120 12314 9172
rect 15654 9160 15660 9172
rect 12360 9132 12572 9160
rect 10505 9095 10563 9101
rect 10505 9092 10517 9095
rect 10192 9064 10517 9092
rect 10192 9052 10198 9064
rect 10505 9061 10517 9064
rect 10551 9092 10563 9095
rect 11425 9095 11483 9101
rect 10551 9064 11100 9092
rect 10551 9061 10563 9064
rect 10505 9055 10563 9061
rect 10870 8984 10876 9036
rect 10928 8984 10934 9036
rect 10965 9027 11023 9033
rect 10965 8993 10977 9027
rect 11011 8993 11023 9027
rect 11072 9024 11100 9064
rect 11425 9061 11437 9095
rect 11471 9061 11483 9095
rect 11425 9055 11483 9061
rect 12066 9052 12072 9104
rect 12124 9092 12130 9104
rect 12360 9092 12388 9132
rect 12124 9064 12388 9092
rect 12124 9052 12130 9064
rect 11974 9024 11980 9036
rect 11072 8996 11980 9024
rect 10965 8987 11023 8993
rect 10980 8956 11008 8987
rect 11974 8984 11980 8996
rect 12032 8984 12038 9036
rect 12434 8984 12440 9036
rect 12492 8984 12498 9036
rect 12544 9033 12572 9132
rect 13832 9132 15660 9160
rect 12986 9052 12992 9104
rect 13044 9052 13050 9104
rect 13832 9033 13860 9132
rect 15654 9120 15660 9132
rect 15712 9120 15718 9172
rect 16117 9163 16175 9169
rect 16117 9129 16129 9163
rect 16163 9160 16175 9163
rect 16390 9160 16396 9172
rect 16163 9132 16396 9160
rect 16163 9129 16175 9132
rect 16117 9123 16175 9129
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 16482 9120 16488 9172
rect 16540 9160 16546 9172
rect 18874 9160 18880 9172
rect 16540 9132 18880 9160
rect 16540 9120 16546 9132
rect 18874 9120 18880 9132
rect 18932 9120 18938 9172
rect 18966 9120 18972 9172
rect 19024 9120 19030 9172
rect 19058 9120 19064 9172
rect 19116 9160 19122 9172
rect 19116 9132 19196 9160
rect 19116 9120 19122 9132
rect 14366 9092 14372 9104
rect 13924 9064 14372 9092
rect 13924 9033 13952 9064
rect 14366 9052 14372 9064
rect 14424 9052 14430 9104
rect 14458 9052 14464 9104
rect 14516 9052 14522 9104
rect 15105 9095 15163 9101
rect 14568 9064 15056 9092
rect 12544 9027 12607 9033
rect 12544 8996 12561 9027
rect 12549 8993 12561 8996
rect 12595 8993 12607 9027
rect 13725 9027 13783 9033
rect 13725 9024 13737 9027
rect 12549 8987 12607 8993
rect 13096 8996 13737 9024
rect 10888 8928 11008 8956
rect 10888 8900 10916 8928
rect 11606 8916 11612 8968
rect 11664 8956 11670 8968
rect 11793 8959 11851 8965
rect 11793 8956 11805 8959
rect 11664 8928 11805 8956
rect 11664 8916 11670 8928
rect 11793 8925 11805 8928
rect 11839 8956 11851 8959
rect 12802 8956 12808 8968
rect 11839 8928 12808 8956
rect 11839 8925 11851 8928
rect 11793 8919 11851 8925
rect 12802 8916 12808 8928
rect 12860 8916 12866 8968
rect 10321 8891 10379 8897
rect 10321 8857 10333 8891
rect 10367 8888 10379 8891
rect 10870 8888 10876 8900
rect 10367 8860 10876 8888
rect 10367 8857 10379 8860
rect 10321 8851 10379 8857
rect 10870 8848 10876 8860
rect 10928 8848 10934 8900
rect 11974 8848 11980 8900
rect 12032 8888 12038 8900
rect 12032 8860 12204 8888
rect 12032 8848 12038 8860
rect 10502 8780 10508 8832
rect 10560 8820 10566 8832
rect 10597 8823 10655 8829
rect 10597 8820 10609 8823
rect 10560 8792 10609 8820
rect 10560 8780 10566 8792
rect 10597 8789 10609 8792
rect 10643 8789 10655 8823
rect 10597 8783 10655 8789
rect 11882 8780 11888 8832
rect 11940 8780 11946 8832
rect 12066 8780 12072 8832
rect 12124 8780 12130 8832
rect 12176 8820 12204 8860
rect 12253 8823 12311 8829
rect 12253 8820 12265 8823
rect 12176 8792 12265 8820
rect 12253 8789 12265 8792
rect 12299 8820 12311 8823
rect 13096 8820 13124 8996
rect 13725 8993 13737 8996
rect 13771 8993 13783 9027
rect 13725 8987 13783 8993
rect 13817 9027 13875 9033
rect 13817 8993 13829 9027
rect 13863 8993 13875 9027
rect 13817 8987 13875 8993
rect 13909 9027 13967 9033
rect 13909 8993 13921 9027
rect 13955 8993 13967 9027
rect 13909 8987 13967 8993
rect 14001 9027 14059 9033
rect 14001 8993 14013 9027
rect 14047 8993 14059 9027
rect 14001 8987 14059 8993
rect 13630 8848 13636 8900
rect 13688 8888 13694 8900
rect 14016 8888 14044 8987
rect 14274 8984 14280 9036
rect 14332 9024 14338 9036
rect 14568 9024 14596 9064
rect 14332 8996 14596 9024
rect 14332 8984 14338 8996
rect 14642 8984 14648 9036
rect 14700 8984 14706 9036
rect 14553 8959 14611 8965
rect 14553 8925 14565 8959
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 13688 8860 14044 8888
rect 13688 8848 13694 8860
rect 12299 8792 13124 8820
rect 13173 8823 13231 8829
rect 12299 8789 12311 8792
rect 12253 8783 12311 8789
rect 13173 8789 13185 8823
rect 13219 8820 13231 8823
rect 13541 8823 13599 8829
rect 13541 8820 13553 8823
rect 13219 8792 13553 8820
rect 13219 8789 13231 8792
rect 13173 8783 13231 8789
rect 13541 8789 13553 8792
rect 13587 8820 13599 8823
rect 14182 8820 14188 8832
rect 13587 8792 14188 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 14182 8780 14188 8792
rect 14240 8780 14246 8832
rect 14568 8820 14596 8919
rect 15028 8888 15056 9064
rect 15105 9061 15117 9095
rect 15151 9092 15163 9095
rect 15562 9092 15568 9104
rect 15151 9064 15568 9092
rect 15151 9061 15163 9064
rect 15105 9055 15163 9061
rect 15562 9052 15568 9064
rect 15620 9052 15626 9104
rect 17770 9052 17776 9104
rect 17828 9052 17834 9104
rect 18414 9052 18420 9104
rect 18472 9052 18478 9104
rect 18509 9095 18567 9101
rect 18509 9061 18521 9095
rect 18555 9092 18567 9095
rect 18984 9092 19012 9120
rect 18555 9064 19012 9092
rect 18555 9061 18567 9064
rect 18509 9055 18567 9061
rect 15194 8984 15200 9036
rect 15252 8984 15258 9036
rect 15470 8984 15476 9036
rect 15528 9024 15534 9036
rect 15657 9027 15715 9033
rect 15657 9024 15669 9027
rect 15528 8996 15669 9024
rect 15528 8984 15534 8996
rect 15657 8993 15669 8996
rect 15703 8993 15715 9027
rect 15657 8987 15715 8993
rect 16758 8984 16764 9036
rect 16816 9024 16822 9036
rect 17037 9027 17095 9033
rect 17037 9024 17049 9027
rect 16816 8996 17049 9024
rect 16816 8984 16822 8996
rect 17037 8993 17049 8996
rect 17083 8993 17095 9027
rect 17037 8987 17095 8993
rect 17218 8984 17224 9036
rect 17276 8984 17282 9036
rect 17310 8984 17316 9036
rect 17368 8984 17374 9036
rect 17494 8984 17500 9036
rect 17552 9024 17558 9036
rect 17957 9027 18015 9033
rect 17957 9024 17969 9027
rect 17552 8996 17969 9024
rect 17552 8984 17558 8996
rect 17957 8993 17969 8996
rect 18003 8993 18015 9027
rect 17957 8987 18015 8993
rect 18138 8984 18144 9036
rect 18196 9024 18202 9036
rect 19168 9033 19196 9132
rect 19978 9120 19984 9172
rect 20036 9160 20042 9172
rect 20036 9132 21220 9160
rect 20036 9120 20042 9132
rect 19705 9095 19763 9101
rect 19705 9061 19717 9095
rect 19751 9092 19763 9095
rect 19794 9092 19800 9104
rect 19751 9064 19800 9092
rect 19751 9061 19763 9064
rect 19705 9055 19763 9061
rect 19794 9052 19800 9064
rect 19852 9052 19858 9104
rect 20346 9052 20352 9104
rect 20404 9052 20410 9104
rect 20898 9092 20904 9104
rect 20456 9064 20904 9092
rect 18969 9027 19027 9033
rect 18969 9024 18981 9027
rect 18196 8996 18981 9024
rect 18196 8984 18202 8996
rect 18969 8993 18981 8996
rect 19015 8993 19027 9027
rect 18969 8987 19027 8993
rect 19153 9027 19211 9033
rect 19153 8993 19165 9027
rect 19199 8993 19211 9027
rect 19153 8987 19211 8993
rect 19242 8984 19248 9036
rect 19300 8984 19306 9036
rect 19426 8984 19432 9036
rect 19484 9024 19490 9036
rect 19886 9024 19892 9036
rect 19484 8996 19892 9024
rect 19484 8984 19490 8996
rect 19886 8984 19892 8996
rect 19944 8984 19950 9036
rect 20456 9033 20484 9064
rect 20898 9052 20904 9064
rect 20956 9052 20962 9104
rect 20990 9052 20996 9104
rect 21048 9052 21054 9104
rect 21192 9092 21220 9132
rect 22370 9120 22376 9172
rect 22428 9160 22434 9172
rect 25958 9160 25964 9172
rect 22428 9132 22508 9160
rect 22428 9120 22434 9132
rect 21192 9064 21404 9092
rect 20441 9027 20499 9033
rect 20441 8993 20453 9027
rect 20487 8993 20499 9027
rect 20441 8987 20499 8993
rect 20530 8984 20536 9036
rect 20588 8984 20594 9036
rect 21082 8984 21088 9036
rect 21140 9030 21146 9036
rect 21376 9033 21404 9064
rect 21634 9052 21640 9104
rect 21692 9092 21698 9104
rect 21821 9095 21879 9101
rect 21821 9092 21833 9095
rect 21692 9064 21833 9092
rect 21692 9052 21698 9064
rect 21821 9061 21833 9064
rect 21867 9061 21879 9095
rect 21821 9055 21879 9061
rect 21913 9095 21971 9101
rect 21913 9061 21925 9095
rect 21959 9092 21971 9095
rect 22186 9092 22192 9104
rect 21959 9064 22192 9092
rect 21959 9061 21971 9064
rect 21913 9055 21971 9061
rect 22186 9052 22192 9064
rect 22244 9052 22250 9104
rect 21269 9030 21327 9033
rect 21140 9027 21327 9030
rect 21140 9002 21281 9027
rect 21140 8984 21146 9002
rect 21269 8993 21281 9002
rect 21315 8993 21327 9027
rect 21269 8987 21327 8993
rect 21361 9027 21419 9033
rect 21361 8993 21373 9027
rect 21407 8993 21419 9027
rect 21361 8987 21419 8993
rect 21726 8984 21732 9036
rect 21784 9024 21790 9036
rect 22373 9027 22431 9033
rect 22373 9024 22385 9027
rect 21784 8996 22385 9024
rect 21784 8984 21790 8996
rect 22373 8993 22385 8996
rect 22419 8993 22431 9027
rect 22480 9024 22508 9132
rect 23860 9132 25964 9160
rect 22554 9052 22560 9104
rect 22612 9092 22618 9104
rect 22612 9064 22784 9092
rect 22612 9052 22618 9064
rect 22756 9033 22784 9064
rect 23014 9052 23020 9104
rect 23072 9092 23078 9104
rect 23201 9095 23259 9101
rect 23201 9092 23213 9095
rect 23072 9064 23213 9092
rect 23072 9052 23078 9064
rect 23201 9061 23213 9064
rect 23247 9061 23259 9095
rect 23201 9055 23259 9061
rect 22649 9027 22707 9033
rect 22649 9024 22661 9027
rect 22480 8996 22661 9024
rect 22373 8987 22431 8993
rect 22649 8993 22661 8996
rect 22695 8993 22707 9027
rect 22649 8987 22707 8993
rect 22741 9027 22799 9033
rect 22741 8993 22753 9027
rect 22787 8993 22799 9027
rect 22741 8987 22799 8993
rect 23750 8984 23756 9036
rect 23808 8984 23814 9036
rect 23860 9033 23888 9132
rect 25958 9120 25964 9132
rect 26016 9120 26022 9172
rect 27065 9163 27123 9169
rect 27065 9129 27077 9163
rect 27111 9160 27123 9163
rect 27798 9160 27804 9172
rect 27111 9132 27804 9160
rect 27111 9129 27123 9132
rect 27065 9123 27123 9129
rect 23937 9095 23995 9101
rect 23937 9061 23949 9095
rect 23983 9092 23995 9095
rect 24026 9092 24032 9104
rect 23983 9064 24032 9092
rect 23983 9061 23995 9064
rect 23937 9055 23995 9061
rect 24026 9052 24032 9064
rect 24084 9052 24090 9104
rect 24670 9052 24676 9104
rect 24728 9052 24734 9104
rect 24762 9052 24768 9104
rect 24820 9092 24826 9104
rect 24857 9095 24915 9101
rect 24857 9092 24869 9095
rect 24820 9064 24869 9092
rect 24820 9052 24826 9064
rect 24857 9061 24869 9064
rect 24903 9061 24915 9095
rect 26602 9092 26608 9104
rect 24857 9055 24915 9061
rect 25428 9064 26608 9092
rect 23845 9027 23903 9033
rect 23845 8993 23857 9027
rect 23891 8993 23903 9027
rect 23845 8987 23903 8993
rect 24397 9027 24455 9033
rect 24397 8993 24409 9027
rect 24443 8993 24455 9027
rect 24688 9024 24716 9052
rect 25428 9033 25456 9064
rect 26602 9052 26608 9064
rect 26660 9052 26666 9104
rect 25317 9027 25375 9033
rect 25317 9024 25329 9027
rect 24688 8996 25329 9024
rect 24397 8987 24455 8993
rect 25317 8993 25329 8996
rect 25363 8993 25375 9027
rect 25317 8987 25375 8993
rect 25409 9027 25467 9033
rect 25409 8993 25421 9027
rect 25455 8993 25467 9027
rect 25409 8987 25467 8993
rect 15749 8959 15807 8965
rect 15749 8925 15761 8959
rect 15795 8956 15807 8959
rect 15930 8956 15936 8968
rect 15795 8928 15936 8956
rect 15795 8925 15807 8928
rect 15749 8919 15807 8925
rect 15930 8916 15936 8928
rect 15988 8916 15994 8968
rect 17129 8959 17187 8965
rect 16224 8928 17080 8956
rect 16224 8888 16252 8928
rect 15028 8860 16252 8888
rect 16301 8891 16359 8897
rect 16301 8857 16313 8891
rect 16347 8888 16359 8891
rect 17052 8888 17080 8928
rect 17129 8925 17141 8959
rect 17175 8956 17187 8959
rect 17402 8956 17408 8968
rect 17175 8928 17408 8956
rect 17175 8925 17187 8928
rect 17129 8919 17187 8925
rect 17402 8916 17408 8928
rect 17460 8916 17466 8968
rect 17770 8916 17776 8968
rect 17828 8956 17834 8968
rect 17865 8959 17923 8965
rect 17865 8956 17877 8959
rect 17828 8928 17877 8956
rect 17828 8916 17834 8928
rect 17865 8925 17877 8928
rect 17911 8925 17923 8959
rect 17865 8919 17923 8925
rect 19061 8959 19119 8965
rect 19061 8925 19073 8959
rect 19107 8925 19119 8959
rect 19061 8919 19119 8925
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8925 19855 8959
rect 19797 8919 19855 8925
rect 17218 8888 17224 8900
rect 16347 8860 16896 8888
rect 17052 8860 17224 8888
rect 16347 8857 16359 8860
rect 16301 8851 16359 8857
rect 16022 8820 16028 8832
rect 14568 8792 16028 8820
rect 16022 8780 16028 8792
rect 16080 8780 16086 8832
rect 16206 8780 16212 8832
rect 16264 8820 16270 8832
rect 16868 8829 16896 8860
rect 17218 8848 17224 8860
rect 17276 8848 17282 8900
rect 16393 8823 16451 8829
rect 16393 8820 16405 8823
rect 16264 8792 16405 8820
rect 16264 8780 16270 8792
rect 16393 8789 16405 8792
rect 16439 8789 16451 8823
rect 16393 8783 16451 8789
rect 16853 8823 16911 8829
rect 16853 8789 16865 8823
rect 16899 8820 16911 8823
rect 17126 8820 17132 8832
rect 16899 8792 17132 8820
rect 16899 8789 16911 8792
rect 16853 8783 16911 8789
rect 17126 8780 17132 8792
rect 17184 8780 17190 8832
rect 19076 8820 19104 8919
rect 19812 8888 19840 8919
rect 20254 8916 20260 8968
rect 20312 8956 20318 8968
rect 22465 8959 22523 8965
rect 20312 8928 22416 8956
rect 20312 8916 20318 8928
rect 22002 8888 22008 8900
rect 19812 8860 22008 8888
rect 22002 8848 22008 8860
rect 22060 8848 22066 8900
rect 22388 8888 22416 8928
rect 22465 8925 22477 8959
rect 22511 8956 22523 8959
rect 23474 8956 23480 8968
rect 22511 8928 23480 8956
rect 22511 8925 22523 8928
rect 22465 8919 22523 8925
rect 23474 8916 23480 8928
rect 23532 8916 23538 8968
rect 23106 8888 23112 8900
rect 22388 8860 23112 8888
rect 23106 8848 23112 8860
rect 23164 8848 23170 8900
rect 23842 8848 23848 8900
rect 23900 8888 23906 8900
rect 24412 8888 24440 8987
rect 25866 8984 25872 9036
rect 25924 9033 25930 9036
rect 25924 9027 25978 9033
rect 25924 8993 25932 9027
rect 25966 8993 25978 9027
rect 25924 8987 25978 8993
rect 26053 9027 26111 9033
rect 26053 8993 26065 9027
rect 26099 9024 26111 9027
rect 26697 9027 26755 9033
rect 26099 8996 26648 9024
rect 26099 8993 26111 8996
rect 26053 8987 26111 8993
rect 25924 8984 25930 8987
rect 24489 8959 24547 8965
rect 24489 8925 24501 8959
rect 24535 8925 24547 8959
rect 24489 8919 24547 8925
rect 23900 8860 24440 8888
rect 24504 8888 24532 8919
rect 24670 8916 24676 8968
rect 24728 8916 24734 8968
rect 25038 8916 25044 8968
rect 25096 8956 25102 8968
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25096 8928 25513 8956
rect 25096 8916 25102 8928
rect 25501 8925 25513 8928
rect 25547 8956 25559 8959
rect 26513 8959 26571 8965
rect 26513 8956 26525 8959
rect 25547 8928 26525 8956
rect 25547 8925 25559 8928
rect 25501 8919 25559 8925
rect 26513 8925 26525 8928
rect 26559 8925 26571 8959
rect 26513 8919 26571 8925
rect 26620 8888 26648 8996
rect 26697 8993 26709 9027
rect 26743 8993 26755 9027
rect 26697 8987 26755 8993
rect 26881 9027 26939 9033
rect 26881 8993 26893 9027
rect 26927 9024 26939 9027
rect 27080 9024 27108 9123
rect 27798 9120 27804 9132
rect 27856 9120 27862 9172
rect 26927 8996 27108 9024
rect 26927 8993 26939 8996
rect 26881 8987 26939 8993
rect 26712 8956 26740 8987
rect 28074 8956 28080 8968
rect 26712 8928 28080 8956
rect 28074 8916 28080 8928
rect 28132 8916 28138 8968
rect 26878 8888 26884 8900
rect 24504 8860 26004 8888
rect 26620 8860 26884 8888
rect 23900 8848 23906 8860
rect 19794 8820 19800 8832
rect 19076 8792 19800 8820
rect 19794 8780 19800 8792
rect 19852 8780 19858 8832
rect 20346 8780 20352 8832
rect 20404 8820 20410 8832
rect 23382 8820 23388 8832
rect 20404 8792 23388 8820
rect 20404 8780 20410 8792
rect 23382 8780 23388 8792
rect 23440 8780 23446 8832
rect 23566 8780 23572 8832
rect 23624 8780 23630 8832
rect 25976 8820 26004 8860
rect 26878 8848 26884 8860
rect 26936 8848 26942 8900
rect 26234 8820 26240 8832
rect 25976 8792 26240 8820
rect 26234 8780 26240 8792
rect 26292 8780 26298 8832
rect 26326 8780 26332 8832
rect 26384 8780 26390 8832
rect 26786 8780 26792 8832
rect 26844 8780 26850 8832
rect 460 8730 43516 8752
rect 460 8678 1306 8730
rect 1358 8678 1370 8730
rect 1422 8678 1434 8730
rect 1486 8678 1498 8730
rect 1550 8678 1562 8730
rect 1614 8678 9306 8730
rect 9358 8678 9370 8730
rect 9422 8678 9434 8730
rect 9486 8678 9498 8730
rect 9550 8678 9562 8730
rect 9614 8678 41306 8730
rect 41358 8678 41370 8730
rect 41422 8678 41434 8730
rect 41486 8678 41498 8730
rect 41550 8678 41562 8730
rect 41614 8678 43516 8730
rect 460 8656 43516 8678
rect 6454 8576 6460 8628
rect 6512 8576 6518 8628
rect 7558 8576 7564 8628
rect 7616 8576 7622 8628
rect 8386 8576 8392 8628
rect 8444 8576 8450 8628
rect 9214 8576 9220 8628
rect 9272 8576 9278 8628
rect 9858 8576 9864 8628
rect 9916 8616 9922 8628
rect 10045 8619 10103 8625
rect 10045 8616 10057 8619
rect 9916 8588 10057 8616
rect 9916 8576 9922 8588
rect 10045 8585 10057 8588
rect 10091 8616 10103 8619
rect 10594 8616 10600 8628
rect 10091 8588 10600 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10594 8576 10600 8588
rect 10652 8576 10658 8628
rect 10965 8619 11023 8625
rect 10965 8585 10977 8619
rect 11011 8616 11023 8619
rect 11977 8619 12035 8625
rect 11011 8588 11284 8616
rect 11011 8585 11023 8588
rect 10965 8579 11023 8585
rect 9030 8508 9036 8560
rect 9088 8548 9094 8560
rect 9769 8551 9827 8557
rect 9769 8548 9781 8551
rect 9088 8520 9781 8548
rect 9088 8508 9094 8520
rect 9769 8517 9781 8520
rect 9815 8517 9827 8551
rect 9769 8511 9827 8517
rect 10502 8508 10508 8560
rect 10560 8548 10566 8560
rect 11256 8548 11284 8588
rect 11977 8585 11989 8619
rect 12023 8616 12035 8619
rect 12345 8619 12403 8625
rect 12345 8616 12357 8619
rect 12023 8588 12357 8616
rect 12023 8585 12035 8588
rect 11977 8579 12035 8585
rect 12345 8585 12357 8588
rect 12391 8616 12403 8619
rect 13906 8616 13912 8628
rect 12391 8588 13912 8616
rect 12391 8585 12403 8588
rect 12345 8579 12403 8585
rect 13906 8576 13912 8588
rect 13964 8576 13970 8628
rect 14277 8619 14335 8625
rect 14277 8585 14289 8619
rect 14323 8616 14335 8619
rect 15286 8616 15292 8628
rect 14323 8588 15292 8616
rect 14323 8585 14335 8588
rect 14277 8579 14335 8585
rect 11330 8548 11336 8560
rect 10560 8520 11192 8548
rect 11256 8520 11336 8548
rect 10560 8508 10566 8520
rect 10134 8440 10140 8492
rect 10192 8440 10198 8492
rect 10686 8440 10692 8492
rect 10744 8440 10750 8492
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 6822 8372 6828 8424
rect 6880 8412 6886 8424
rect 7653 8415 7711 8421
rect 7653 8412 7665 8415
rect 6880 8384 7665 8412
rect 6880 8372 6886 8384
rect 7653 8381 7665 8384
rect 7699 8381 7711 8415
rect 7653 8375 7711 8381
rect 8018 8372 8024 8424
rect 8076 8412 8082 8424
rect 9309 8415 9367 8421
rect 9309 8412 9321 8415
rect 8076 8384 9321 8412
rect 8076 8372 8082 8384
rect 9309 8381 9321 8384
rect 9355 8412 9367 8415
rect 9490 8412 9496 8424
rect 9355 8384 9496 8412
rect 9355 8381 9367 8384
rect 9309 8375 9367 8381
rect 9490 8372 9496 8384
rect 9548 8372 9554 8424
rect 9674 8372 9680 8424
rect 9732 8412 9738 8424
rect 11164 8421 11192 8520
rect 11330 8508 11336 8520
rect 11388 8548 11394 8560
rect 12526 8548 12532 8560
rect 11388 8520 12532 8548
rect 11388 8508 11394 8520
rect 12526 8508 12532 8520
rect 12584 8508 12590 8560
rect 13725 8551 13783 8557
rect 13725 8517 13737 8551
rect 13771 8548 13783 8551
rect 14292 8548 14320 8579
rect 15286 8576 15292 8588
rect 15344 8576 15350 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16390 8616 16396 8628
rect 16347 8588 16396 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16390 8576 16396 8588
rect 16448 8576 16454 8628
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8616 16911 8619
rect 17405 8619 17463 8625
rect 17405 8616 17417 8619
rect 16899 8588 17417 8616
rect 16899 8585 16911 8588
rect 16853 8579 16911 8585
rect 17405 8585 17417 8588
rect 17451 8616 17463 8619
rect 17586 8616 17592 8628
rect 17451 8588 17592 8616
rect 17451 8585 17463 8588
rect 17405 8579 17463 8585
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 18049 8619 18107 8625
rect 18049 8585 18061 8619
rect 18095 8616 18107 8619
rect 18506 8616 18512 8628
rect 18095 8588 18512 8616
rect 18095 8585 18107 8588
rect 18049 8579 18107 8585
rect 14918 8548 14924 8560
rect 13771 8520 14320 8548
rect 14476 8520 14924 8548
rect 13771 8517 13783 8520
rect 13725 8511 13783 8517
rect 11606 8440 11612 8492
rect 11664 8440 11670 8492
rect 11793 8483 11851 8489
rect 11793 8449 11805 8483
rect 11839 8480 11851 8483
rect 12158 8480 12164 8492
rect 11839 8452 12164 8480
rect 11839 8449 11851 8452
rect 11793 8443 11851 8449
rect 12158 8440 12164 8452
rect 12216 8480 12222 8492
rect 13265 8483 13323 8489
rect 12216 8452 12848 8480
rect 12216 8440 12222 8452
rect 10597 8415 10655 8421
rect 10597 8412 10609 8415
rect 9732 8384 10609 8412
rect 9732 8372 9738 8384
rect 10597 8381 10609 8384
rect 10643 8381 10655 8415
rect 10597 8375 10655 8381
rect 11149 8415 11207 8421
rect 11149 8381 11161 8415
rect 11195 8381 11207 8415
rect 11149 8375 11207 8381
rect 11422 8372 11428 8424
rect 11480 8412 11486 8424
rect 11882 8412 11888 8424
rect 11480 8384 11888 8412
rect 11480 8372 11486 8384
rect 11882 8372 11888 8384
rect 11940 8412 11946 8424
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 11940 8384 12541 8412
rect 11940 8372 11946 8384
rect 12529 8381 12541 8384
rect 12575 8381 12587 8415
rect 12529 8375 12587 8381
rect 12618 8372 12624 8424
rect 12676 8372 12682 8424
rect 12820 8421 12848 8452
rect 13265 8449 13277 8483
rect 13311 8480 13323 8483
rect 13814 8480 13820 8492
rect 13311 8452 13820 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13814 8440 13820 8452
rect 13872 8440 13878 8492
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8480 13967 8483
rect 14366 8480 14372 8492
rect 13955 8452 14372 8480
rect 13955 8449 13967 8452
rect 13909 8443 13967 8449
rect 14366 8440 14372 8452
rect 14424 8440 14430 8492
rect 14476 8480 14504 8520
rect 14918 8508 14924 8520
rect 14976 8508 14982 8560
rect 16942 8548 16948 8560
rect 15212 8520 16948 8548
rect 14543 8483 14601 8489
rect 14543 8480 14555 8483
rect 14476 8452 14555 8480
rect 14543 8449 14555 8452
rect 14589 8449 14601 8483
rect 14543 8443 14601 8449
rect 14645 8483 14703 8489
rect 14645 8449 14657 8483
rect 14691 8480 14703 8483
rect 15010 8480 15016 8492
rect 14691 8452 15016 8480
rect 14691 8449 14703 8452
rect 14645 8443 14703 8449
rect 15010 8440 15016 8452
rect 15068 8440 15074 8492
rect 15212 8489 15240 8520
rect 16942 8508 16948 8520
rect 17000 8508 17006 8560
rect 17037 8551 17095 8557
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 18064 8548 18092 8579
rect 18506 8576 18512 8588
rect 18564 8576 18570 8628
rect 18969 8619 19027 8625
rect 18969 8585 18981 8619
rect 19015 8616 19027 8619
rect 19150 8616 19156 8628
rect 19015 8588 19156 8616
rect 19015 8585 19027 8588
rect 18969 8579 19027 8585
rect 19150 8576 19156 8588
rect 19208 8576 19214 8628
rect 19613 8619 19671 8625
rect 19613 8585 19625 8619
rect 19659 8616 19671 8619
rect 19702 8616 19708 8628
rect 19659 8588 19708 8616
rect 19659 8585 19671 8588
rect 19613 8579 19671 8585
rect 19702 8576 19708 8588
rect 19760 8576 19766 8628
rect 20993 8619 21051 8625
rect 20993 8585 21005 8619
rect 21039 8616 21051 8619
rect 21545 8619 21603 8625
rect 21545 8616 21557 8619
rect 21039 8588 21557 8616
rect 21039 8585 21051 8588
rect 20993 8579 21051 8585
rect 21545 8585 21557 8588
rect 21591 8616 21603 8619
rect 21910 8616 21916 8628
rect 21591 8588 21916 8616
rect 21591 8585 21603 8588
rect 21545 8579 21603 8585
rect 21910 8576 21916 8588
rect 21968 8576 21974 8628
rect 22738 8576 22744 8628
rect 22796 8616 22802 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22796 8588 22845 8616
rect 22796 8576 22802 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 25406 8616 25412 8628
rect 22833 8579 22891 8585
rect 23676 8588 25412 8616
rect 20254 8548 20260 8560
rect 17083 8520 18092 8548
rect 18708 8520 20260 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 15197 8483 15255 8489
rect 15197 8449 15209 8483
rect 15243 8449 15255 8483
rect 15197 8443 15255 8449
rect 15289 8483 15347 8489
rect 15289 8449 15301 8483
rect 15335 8480 15347 8483
rect 15841 8483 15899 8489
rect 15335 8452 15792 8480
rect 15335 8449 15347 8452
rect 15289 8443 15347 8449
rect 12713 8415 12771 8421
rect 12713 8381 12725 8415
rect 12759 8381 12771 8415
rect 12713 8375 12771 8381
rect 12805 8415 12863 8421
rect 12805 8381 12817 8415
rect 12851 8381 12863 8415
rect 14461 8415 14519 8421
rect 14461 8412 14473 8415
rect 12805 8375 12863 8381
rect 13464 8384 14473 8412
rect 5258 8304 5264 8356
rect 5316 8344 5322 8356
rect 6638 8344 6644 8356
rect 5316 8316 6644 8344
rect 5316 8304 5322 8316
rect 6638 8304 6644 8316
rect 6696 8304 6702 8356
rect 6914 8304 6920 8356
rect 6972 8344 6978 8356
rect 8570 8344 8576 8356
rect 6972 8316 8576 8344
rect 6972 8304 6978 8316
rect 8570 8304 8576 8316
rect 8628 8304 8634 8356
rect 10686 8344 10692 8356
rect 9968 8316 10692 8344
rect 5442 8236 5448 8288
rect 5500 8276 5506 8288
rect 5537 8279 5595 8285
rect 5537 8276 5549 8279
rect 5500 8248 5549 8276
rect 5500 8236 5506 8248
rect 5537 8245 5549 8248
rect 5583 8245 5595 8279
rect 5537 8239 5595 8245
rect 5813 8279 5871 8285
rect 5813 8245 5825 8279
rect 5859 8276 5871 8279
rect 5994 8276 6000 8288
rect 5859 8248 6000 8276
rect 5859 8245 5871 8248
rect 5813 8239 5871 8245
rect 5994 8236 6000 8248
rect 6052 8236 6058 8288
rect 6362 8236 6368 8288
rect 6420 8276 6426 8288
rect 9968 8276 9996 8316
rect 10686 8304 10692 8316
rect 10744 8304 10750 8356
rect 12728 8344 12756 8375
rect 13464 8356 13492 8384
rect 14461 8381 14473 8384
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 14734 8372 14740 8424
rect 14792 8372 14798 8424
rect 15378 8372 15384 8424
rect 15436 8372 15442 8424
rect 15764 8412 15792 8452
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16114 8480 16120 8492
rect 15887 8452 16120 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 16264 8452 17632 8480
rect 16264 8440 16270 8452
rect 15764 8384 16436 8412
rect 13262 8344 13268 8356
rect 12728 8316 13268 8344
rect 13262 8304 13268 8316
rect 13320 8304 13326 8356
rect 13446 8304 13452 8356
rect 13504 8304 13510 8356
rect 13998 8304 14004 8356
rect 14056 8344 14062 8356
rect 14056 8316 15976 8344
rect 14056 8304 14062 8316
rect 6420 8248 9996 8276
rect 6420 8236 6426 8248
rect 10410 8236 10416 8288
rect 10468 8276 10474 8288
rect 15838 8276 15844 8288
rect 10468 8248 15844 8276
rect 10468 8236 10474 8248
rect 15838 8236 15844 8248
rect 15896 8236 15902 8288
rect 15948 8276 15976 8316
rect 16022 8304 16028 8356
rect 16080 8344 16086 8356
rect 16298 8344 16304 8356
rect 16080 8316 16304 8344
rect 16080 8304 16086 8316
rect 16298 8304 16304 8316
rect 16356 8304 16362 8356
rect 16408 8344 16436 8384
rect 16482 8372 16488 8424
rect 16540 8372 16546 8424
rect 16574 8372 16580 8424
rect 16632 8372 16638 8424
rect 17604 8421 17632 8452
rect 17678 8440 17684 8492
rect 17736 8440 17742 8492
rect 18708 8489 18736 8520
rect 20254 8508 20260 8520
rect 20312 8508 20318 8560
rect 22002 8548 22008 8560
rect 21928 8520 22008 8548
rect 18693 8483 18751 8489
rect 17788 8452 18460 8480
rect 17589 8415 17647 8421
rect 17589 8381 17601 8415
rect 17635 8381 17647 8415
rect 17589 8375 17647 8381
rect 16408 8316 17632 8344
rect 17310 8276 17316 8288
rect 15948 8248 17316 8276
rect 17310 8236 17316 8248
rect 17368 8236 17374 8288
rect 17604 8276 17632 8316
rect 17678 8304 17684 8356
rect 17736 8344 17742 8356
rect 17788 8344 17816 8452
rect 17862 8372 17868 8424
rect 17920 8412 17926 8424
rect 18233 8415 18291 8421
rect 18233 8412 18245 8415
rect 17920 8384 18245 8412
rect 17920 8372 17926 8384
rect 18233 8381 18245 8384
rect 18279 8381 18291 8415
rect 18233 8375 18291 8381
rect 18325 8415 18383 8421
rect 18325 8381 18337 8415
rect 18371 8381 18383 8415
rect 18432 8412 18460 8452
rect 18693 8449 18705 8483
rect 18739 8449 18751 8483
rect 18693 8443 18751 8449
rect 19337 8483 19395 8489
rect 19337 8449 19349 8483
rect 19383 8480 19395 8483
rect 20346 8480 20352 8492
rect 19383 8452 20352 8480
rect 19383 8449 19395 8452
rect 19337 8443 19395 8449
rect 20346 8440 20352 8452
rect 20404 8440 20410 8492
rect 20533 8483 20591 8489
rect 20533 8449 20545 8483
rect 20579 8480 20591 8483
rect 21450 8480 21456 8492
rect 20579 8452 21456 8480
rect 20579 8449 20591 8452
rect 20533 8443 20591 8449
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 21928 8489 21956 8520
rect 22002 8508 22008 8520
rect 22060 8508 22066 8560
rect 21913 8483 21971 8489
rect 21913 8449 21925 8483
rect 21959 8449 21971 8483
rect 21913 8443 21971 8449
rect 22462 8440 22468 8492
rect 22520 8480 22526 8492
rect 23201 8483 23259 8489
rect 23201 8480 23213 8483
rect 22520 8452 23213 8480
rect 22520 8440 22526 8452
rect 23201 8449 23213 8452
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 18598 8412 18604 8424
rect 18432 8384 18604 8412
rect 18325 8375 18383 8381
rect 17736 8316 17816 8344
rect 18340 8344 18368 8375
rect 18598 8372 18604 8384
rect 18656 8412 18662 8424
rect 18785 8415 18843 8421
rect 18785 8412 18797 8415
rect 18656 8384 18797 8412
rect 18656 8372 18662 8384
rect 18785 8381 18797 8384
rect 18831 8381 18843 8415
rect 18785 8375 18843 8381
rect 19426 8372 19432 8424
rect 19484 8372 19490 8424
rect 20438 8372 20444 8424
rect 20496 8372 20502 8424
rect 20714 8372 20720 8424
rect 20772 8412 20778 8424
rect 21174 8412 21180 8424
rect 20772 8384 21180 8412
rect 20772 8372 20778 8384
rect 21174 8372 21180 8384
rect 21232 8372 21238 8424
rect 21358 8372 21364 8424
rect 21416 8412 21422 8424
rect 21726 8412 21732 8424
rect 21416 8384 21732 8412
rect 21416 8372 21422 8384
rect 21726 8372 21732 8384
rect 21784 8372 21790 8424
rect 21818 8372 21824 8424
rect 21876 8372 21882 8424
rect 22005 8415 22063 8421
rect 22005 8381 22017 8415
rect 22051 8381 22063 8415
rect 22005 8375 22063 8381
rect 19886 8344 19892 8356
rect 18340 8316 19892 8344
rect 17736 8304 17742 8316
rect 19886 8304 19892 8316
rect 19944 8304 19950 8356
rect 19981 8347 20039 8353
rect 19981 8313 19993 8347
rect 20027 8344 20039 8347
rect 20162 8344 20168 8356
rect 20027 8316 20168 8344
rect 20027 8313 20039 8316
rect 19981 8307 20039 8313
rect 20162 8304 20168 8316
rect 20220 8304 20226 8356
rect 20990 8276 20996 8288
rect 17604 8248 20996 8276
rect 20990 8236 20996 8248
rect 21048 8236 21054 8288
rect 21174 8236 21180 8288
rect 21232 8276 21238 8288
rect 22020 8276 22048 8375
rect 23014 8372 23020 8424
rect 23072 8372 23078 8424
rect 23109 8415 23167 8421
rect 23109 8381 23121 8415
rect 23155 8412 23167 8415
rect 23676 8412 23704 8588
rect 25406 8576 25412 8588
rect 25464 8576 25470 8628
rect 25774 8576 25780 8628
rect 25832 8616 25838 8628
rect 26605 8619 26663 8625
rect 26605 8616 26617 8619
rect 25832 8588 26617 8616
rect 25832 8576 25838 8588
rect 26605 8585 26617 8588
rect 26651 8616 26663 8619
rect 27157 8619 27215 8625
rect 27157 8616 27169 8619
rect 26651 8588 27169 8616
rect 26651 8585 26663 8588
rect 26605 8579 26663 8585
rect 27157 8585 27169 8588
rect 27203 8585 27215 8619
rect 27157 8579 27215 8585
rect 26142 8548 26148 8560
rect 24320 8520 26148 8548
rect 23934 8480 23940 8492
rect 23155 8384 23704 8412
rect 23768 8452 23940 8480
rect 23155 8381 23167 8384
rect 23109 8375 23167 8381
rect 23032 8344 23060 8372
rect 23768 8353 23796 8452
rect 23934 8440 23940 8452
rect 23992 8440 23998 8492
rect 24320 8489 24348 8520
rect 26142 8508 26148 8520
rect 26200 8508 26206 8560
rect 24305 8483 24363 8489
rect 24305 8449 24317 8483
rect 24351 8449 24363 8483
rect 24305 8443 24363 8449
rect 25866 8440 25872 8492
rect 25924 8480 25930 8492
rect 26053 8483 26111 8489
rect 26053 8480 26065 8483
rect 25924 8452 26065 8480
rect 25924 8440 25930 8452
rect 26053 8449 26065 8452
rect 26099 8449 26111 8483
rect 26053 8443 26111 8449
rect 24118 8372 24124 8424
rect 24176 8412 24182 8424
rect 24213 8415 24271 8421
rect 24213 8412 24225 8415
rect 24176 8384 24225 8412
rect 24176 8372 24182 8384
rect 24213 8381 24225 8384
rect 24259 8381 24271 8415
rect 24213 8375 24271 8381
rect 24857 8415 24915 8421
rect 24857 8381 24869 8415
rect 24903 8381 24915 8415
rect 24857 8375 24915 8381
rect 23385 8347 23443 8353
rect 23385 8344 23397 8347
rect 23032 8316 23397 8344
rect 23385 8313 23397 8316
rect 23431 8313 23443 8347
rect 23385 8307 23443 8313
rect 23753 8347 23811 8353
rect 23753 8313 23765 8347
rect 23799 8313 23811 8347
rect 23753 8307 23811 8313
rect 24394 8304 24400 8356
rect 24452 8304 24458 8356
rect 24670 8304 24676 8356
rect 24728 8344 24734 8356
rect 24872 8344 24900 8375
rect 24946 8372 24952 8424
rect 25004 8372 25010 8424
rect 25038 8372 25044 8424
rect 25096 8372 25102 8424
rect 25498 8372 25504 8424
rect 25556 8372 25562 8424
rect 25593 8415 25651 8421
rect 25593 8381 25605 8415
rect 25639 8412 25651 8415
rect 26510 8412 26516 8424
rect 25639 8384 26516 8412
rect 25639 8381 25651 8384
rect 25593 8375 25651 8381
rect 26510 8372 26516 8384
rect 26568 8372 26574 8424
rect 26602 8372 26608 8424
rect 26660 8412 26666 8424
rect 26789 8415 26847 8421
rect 26789 8412 26801 8415
rect 26660 8384 26801 8412
rect 26660 8372 26666 8384
rect 26789 8381 26801 8384
rect 26835 8381 26847 8415
rect 26789 8375 26847 8381
rect 26881 8415 26939 8421
rect 26881 8381 26893 8415
rect 26927 8412 26939 8415
rect 27062 8412 27068 8424
rect 26927 8384 27068 8412
rect 26927 8381 26939 8384
rect 26881 8375 26939 8381
rect 24728 8316 24900 8344
rect 25516 8344 25544 8372
rect 25869 8347 25927 8353
rect 25869 8344 25881 8347
rect 25516 8316 25881 8344
rect 24728 8304 24734 8316
rect 25869 8313 25881 8316
rect 25915 8313 25927 8347
rect 26804 8344 26832 8375
rect 27062 8372 27068 8384
rect 27120 8372 27126 8424
rect 26973 8347 27031 8353
rect 26973 8344 26985 8347
rect 26804 8316 26985 8344
rect 25869 8307 25927 8313
rect 26973 8313 26985 8316
rect 27019 8313 27031 8347
rect 26973 8307 27031 8313
rect 27246 8304 27252 8356
rect 27304 8344 27310 8356
rect 31846 8344 31852 8356
rect 27304 8316 31852 8344
rect 27304 8304 27310 8316
rect 31846 8304 31852 8316
rect 31904 8304 31910 8356
rect 21232 8248 22048 8276
rect 21232 8236 21238 8248
rect 23934 8236 23940 8288
rect 23992 8276 23998 8288
rect 25685 8279 25743 8285
rect 25685 8276 25697 8279
rect 23992 8248 25697 8276
rect 23992 8236 23998 8248
rect 25685 8245 25697 8248
rect 25731 8245 25743 8279
rect 25685 8239 25743 8245
rect 460 8186 43516 8208
rect 460 8134 1946 8186
rect 1998 8134 2010 8186
rect 2062 8134 2074 8186
rect 2126 8134 2138 8186
rect 2190 8134 2202 8186
rect 2254 8134 9946 8186
rect 9998 8134 10010 8186
rect 10062 8134 10074 8186
rect 10126 8134 10138 8186
rect 10190 8134 10202 8186
rect 10254 8134 33946 8186
rect 33998 8134 34010 8186
rect 34062 8134 34074 8186
rect 34126 8134 34138 8186
rect 34190 8134 34202 8186
rect 34254 8134 41946 8186
rect 41998 8134 42010 8186
rect 42062 8134 42074 8186
rect 42126 8134 42138 8186
rect 42190 8134 42202 8186
rect 42254 8134 43516 8186
rect 460 8112 43516 8134
rect 4246 8032 4252 8084
rect 4304 8072 4310 8084
rect 4433 8075 4491 8081
rect 4433 8072 4445 8075
rect 4304 8044 4445 8072
rect 4304 8032 4310 8044
rect 4433 8041 4445 8044
rect 4479 8072 4491 8075
rect 5074 8072 5080 8084
rect 4479 8044 5080 8072
rect 4479 8041 4491 8044
rect 4433 8035 4491 8041
rect 5074 8032 5080 8044
rect 5132 8032 5138 8084
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 6178 8072 6184 8084
rect 5592 8044 6184 8072
rect 5592 8032 5598 8044
rect 6178 8032 6184 8044
rect 6236 8032 6242 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6604 8044 6745 8072
rect 6604 8032 6610 8044
rect 6733 8041 6745 8044
rect 6779 8072 6791 8075
rect 7282 8072 7288 8084
rect 6779 8044 7288 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 7282 8032 7288 8044
rect 7340 8032 7346 8084
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 8110 8072 8116 8084
rect 7524 8044 8116 8072
rect 7524 8032 7530 8044
rect 8110 8032 8116 8044
rect 8168 8032 8174 8084
rect 9125 8075 9183 8081
rect 9125 8041 9137 8075
rect 9171 8072 9183 8075
rect 10318 8072 10324 8084
rect 9171 8044 10324 8072
rect 9171 8041 9183 8044
rect 9125 8035 9183 8041
rect 4338 7964 4344 8016
rect 4396 8004 4402 8016
rect 5994 8004 6000 8016
rect 4396 7976 6000 8004
rect 4396 7964 4402 7976
rect 5828 7945 5856 7976
rect 5994 7964 6000 7976
rect 6052 7964 6058 8016
rect 6273 8007 6331 8013
rect 6273 7973 6285 8007
rect 6319 8004 6331 8007
rect 6454 8004 6460 8016
rect 6319 7976 6460 8004
rect 6319 7973 6331 7976
rect 6273 7967 6331 7973
rect 6454 7964 6460 7976
rect 6512 7964 6518 8016
rect 6822 8004 6828 8016
rect 6564 7976 6828 8004
rect 5169 7939 5227 7945
rect 5169 7936 5181 7939
rect 4172 7908 5181 7936
rect 2774 7692 2780 7744
rect 2832 7732 2838 7744
rect 4172 7741 4200 7908
rect 5169 7905 5181 7908
rect 5215 7905 5227 7939
rect 5169 7899 5227 7905
rect 5813 7939 5871 7945
rect 5813 7905 5825 7939
rect 5859 7905 5871 7939
rect 5813 7899 5871 7905
rect 6086 7896 6092 7948
rect 6144 7936 6150 7948
rect 6564 7936 6592 7976
rect 6822 7964 6828 7976
rect 6880 8004 6886 8016
rect 7377 8007 7435 8013
rect 6880 7976 7236 8004
rect 6880 7964 6886 7976
rect 6144 7908 6592 7936
rect 6144 7896 6150 7908
rect 6638 7896 6644 7948
rect 6696 7936 6702 7948
rect 6917 7939 6975 7945
rect 6917 7936 6929 7939
rect 6696 7908 6929 7936
rect 6696 7896 6702 7908
rect 6917 7905 6929 7908
rect 6963 7905 6975 7939
rect 7208 7936 7236 7976
rect 7377 7973 7389 8007
rect 7423 8004 7435 8007
rect 7558 8004 7564 8016
rect 7423 7976 7564 8004
rect 7423 7973 7435 7976
rect 7377 7967 7435 7973
rect 7558 7964 7564 7976
rect 7616 7964 7622 8016
rect 8205 8007 8263 8013
rect 8205 7973 8217 8007
rect 8251 8004 8263 8007
rect 8386 8004 8392 8016
rect 8251 7976 8392 8004
rect 8251 7973 8263 7976
rect 8205 7967 8263 7973
rect 8386 7964 8392 7976
rect 8444 7964 8450 8016
rect 9033 8007 9091 8013
rect 8496 7976 8984 8004
rect 7745 7939 7803 7945
rect 7745 7936 7757 7939
rect 7208 7908 7757 7936
rect 6917 7899 6975 7905
rect 7745 7905 7757 7908
rect 7791 7905 7803 7939
rect 8496 7936 8524 7976
rect 7745 7899 7803 7905
rect 8404 7908 8524 7936
rect 5261 7871 5319 7877
rect 5261 7868 5273 7871
rect 5184 7840 5273 7868
rect 5184 7812 5212 7840
rect 5261 7837 5273 7840
rect 5307 7837 5319 7871
rect 5261 7831 5319 7837
rect 5721 7871 5779 7877
rect 5721 7837 5733 7871
rect 5767 7837 5779 7871
rect 5721 7831 5779 7837
rect 5166 7760 5172 7812
rect 5224 7760 5230 7812
rect 5736 7800 5764 7831
rect 6822 7828 6828 7880
rect 6880 7828 6886 7880
rect 7653 7871 7711 7877
rect 7653 7837 7665 7871
rect 7699 7868 7711 7871
rect 8404 7868 8432 7908
rect 8570 7896 8576 7948
rect 8628 7896 8634 7948
rect 7699 7840 8432 7868
rect 8481 7871 8539 7877
rect 7699 7837 7711 7840
rect 7653 7831 7711 7837
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8956 7868 8984 7976
rect 9033 7973 9045 8007
rect 9079 8004 9091 8007
rect 9214 8004 9220 8016
rect 9079 7976 9220 8004
rect 9079 7973 9091 7976
rect 9033 7967 9091 7973
rect 9214 7964 9220 7976
rect 9272 7964 9278 8016
rect 9324 8013 9352 8044
rect 10318 8032 10324 8044
rect 10376 8032 10382 8084
rect 10612 8044 10916 8072
rect 9309 8007 9367 8013
rect 9309 7973 9321 8007
rect 9355 7973 9367 8007
rect 9309 7967 9367 7973
rect 9490 7964 9496 8016
rect 9548 8004 9554 8016
rect 10612 8004 10640 8044
rect 9548 7976 9812 8004
rect 9548 7964 9554 7976
rect 9784 7945 9812 7976
rect 9876 7976 10640 8004
rect 10888 8004 10916 8044
rect 10962 8032 10968 8084
rect 11020 8032 11026 8084
rect 11238 8032 11244 8084
rect 11296 8072 11302 8084
rect 13998 8072 14004 8084
rect 11296 8044 14004 8072
rect 11296 8032 11302 8044
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 14550 8032 14556 8084
rect 14608 8072 14614 8084
rect 18598 8072 18604 8084
rect 14608 8044 18604 8072
rect 14608 8032 14614 8044
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 18690 8032 18696 8084
rect 18748 8072 18754 8084
rect 19518 8072 19524 8084
rect 18748 8044 19524 8072
rect 18748 8032 18754 8044
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 19794 8032 19800 8084
rect 19852 8072 19858 8084
rect 23198 8072 23204 8084
rect 19852 8044 23204 8072
rect 19852 8032 19858 8044
rect 23198 8032 23204 8044
rect 23256 8032 23262 8084
rect 23474 8032 23480 8084
rect 23532 8072 23538 8084
rect 25038 8072 25044 8084
rect 23532 8044 25044 8072
rect 23532 8032 23538 8044
rect 25038 8032 25044 8044
rect 25096 8032 25102 8084
rect 29178 8032 29184 8084
rect 29236 8072 29242 8084
rect 34974 8072 34980 8084
rect 29236 8044 34980 8072
rect 29236 8032 29242 8044
rect 34974 8032 34980 8044
rect 35032 8032 35038 8084
rect 17126 8004 17132 8016
rect 10888 7976 17132 8004
rect 9876 7945 9904 7976
rect 17126 7964 17132 7976
rect 17184 7964 17190 8016
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 17954 8004 17960 8016
rect 17276 7976 17960 8004
rect 17276 7964 17282 7976
rect 17954 7964 17960 7976
rect 18012 7964 18018 8016
rect 18874 7964 18880 8016
rect 18932 8004 18938 8016
rect 20254 8004 20260 8016
rect 18932 7976 20260 8004
rect 18932 7964 18938 7976
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 21082 7964 21088 8016
rect 21140 8004 21146 8016
rect 24670 8004 24676 8016
rect 21140 7976 24676 8004
rect 21140 7964 21146 7976
rect 24670 7964 24676 7976
rect 24728 7964 24734 8016
rect 30098 7964 30104 8016
rect 30156 8004 30162 8016
rect 36078 8004 36084 8016
rect 30156 7976 36084 8004
rect 30156 7964 30162 7976
rect 36078 7964 36084 7976
rect 36136 7964 36142 8016
rect 9769 7939 9827 7945
rect 9769 7905 9781 7939
rect 9815 7905 9827 7939
rect 9769 7899 9827 7905
rect 9861 7939 9919 7945
rect 9861 7905 9873 7939
rect 9907 7905 9919 7939
rect 9861 7899 9919 7905
rect 10045 7939 10103 7945
rect 10045 7905 10057 7939
rect 10091 7936 10103 7939
rect 10229 7939 10287 7945
rect 10229 7936 10241 7939
rect 10091 7908 10241 7936
rect 10091 7905 10103 7908
rect 10045 7899 10103 7905
rect 10229 7905 10241 7908
rect 10275 7936 10287 7939
rect 16390 7936 16396 7948
rect 10275 7908 10364 7936
rect 10275 7905 10287 7908
rect 10229 7899 10287 7905
rect 10336 7880 10364 7908
rect 10612 7908 16396 7936
rect 9950 7868 9956 7880
rect 8956 7840 9956 7868
rect 8481 7831 8539 7837
rect 8496 7800 8524 7831
rect 9950 7828 9956 7840
rect 10008 7828 10014 7880
rect 10134 7828 10140 7880
rect 10192 7828 10198 7880
rect 10318 7828 10324 7880
rect 10376 7828 10382 7880
rect 10612 7800 10640 7908
rect 16390 7896 16396 7908
rect 16448 7896 16454 7948
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 20622 7936 20628 7948
rect 16540 7908 20628 7936
rect 16540 7896 16546 7908
rect 20622 7896 20628 7908
rect 20680 7896 20686 7948
rect 20806 7896 20812 7948
rect 20864 7936 20870 7948
rect 20864 7908 23612 7936
rect 20864 7896 20870 7908
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 11330 7868 11336 7880
rect 10735 7840 11336 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 11330 7828 11336 7840
rect 11388 7828 11394 7880
rect 11882 7828 11888 7880
rect 11940 7868 11946 7880
rect 14734 7868 14740 7880
rect 11940 7840 14740 7868
rect 11940 7828 11946 7840
rect 14734 7828 14740 7840
rect 14792 7828 14798 7880
rect 15102 7828 15108 7880
rect 15160 7868 15166 7880
rect 18690 7868 18696 7880
rect 15160 7840 18696 7868
rect 15160 7828 15166 7840
rect 18690 7828 18696 7840
rect 18748 7828 18754 7880
rect 19886 7828 19892 7880
rect 19944 7868 19950 7880
rect 22462 7868 22468 7880
rect 19944 7840 22468 7868
rect 19944 7828 19950 7840
rect 22462 7828 22468 7840
rect 22520 7828 22526 7880
rect 5736 7772 8432 7800
rect 8496 7772 10640 7800
rect 10980 7772 11744 7800
rect 4157 7735 4215 7741
rect 4157 7732 4169 7735
rect 2832 7704 4169 7732
rect 2832 7692 2838 7704
rect 4157 7701 4169 7704
rect 4203 7701 4215 7735
rect 4157 7695 4215 7701
rect 4617 7735 4675 7741
rect 4617 7701 4629 7735
rect 4663 7732 4675 7735
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 4663 7704 4997 7732
rect 4663 7701 4675 7704
rect 4617 7695 4675 7701
rect 4985 7701 4997 7704
rect 5031 7732 5043 7735
rect 5350 7732 5356 7744
rect 5031 7704 5356 7732
rect 5031 7701 5043 7704
rect 4985 7695 5043 7701
rect 5350 7692 5356 7704
rect 5408 7692 5414 7744
rect 5810 7692 5816 7744
rect 5868 7732 5874 7744
rect 6454 7732 6460 7744
rect 5868 7704 6460 7732
rect 5868 7692 5874 7704
rect 6454 7692 6460 7704
rect 6512 7692 6518 7744
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 8202 7732 8208 7744
rect 7248 7704 8208 7732
rect 7248 7692 7254 7704
rect 8202 7692 8208 7704
rect 8260 7732 8266 7744
rect 8297 7735 8355 7741
rect 8297 7732 8309 7735
rect 8260 7704 8309 7732
rect 8260 7692 8266 7704
rect 8297 7701 8309 7704
rect 8343 7701 8355 7735
rect 8404 7732 8432 7772
rect 10980 7732 11008 7772
rect 8404 7704 11008 7732
rect 8297 7695 8355 7701
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11149 7735 11207 7741
rect 11149 7732 11161 7735
rect 11112 7704 11161 7732
rect 11112 7692 11118 7704
rect 11149 7701 11161 7704
rect 11195 7701 11207 7735
rect 11149 7695 11207 7701
rect 460 7642 11592 7664
rect 460 7590 1306 7642
rect 1358 7590 1370 7642
rect 1422 7590 1434 7642
rect 1486 7590 1498 7642
rect 1550 7590 1562 7642
rect 1614 7590 9306 7642
rect 9358 7590 9370 7642
rect 9422 7590 9434 7642
rect 9486 7590 9498 7642
rect 9550 7590 9562 7642
rect 9614 7590 11592 7642
rect 460 7568 11592 7590
rect 11716 7596 11744 7772
rect 13538 7760 13544 7812
rect 13596 7800 13602 7812
rect 19150 7800 19156 7812
rect 13596 7772 19156 7800
rect 13596 7760 13602 7772
rect 19150 7760 19156 7772
rect 19208 7760 19214 7812
rect 23584 7744 23612 7908
rect 29362 7828 29368 7880
rect 29420 7868 29426 7880
rect 35250 7868 35256 7880
rect 29420 7840 35256 7868
rect 29420 7828 29426 7840
rect 35250 7828 35256 7840
rect 35308 7828 35314 7880
rect 29914 7760 29920 7812
rect 29972 7800 29978 7812
rect 36446 7800 36452 7812
rect 29972 7772 36452 7800
rect 29972 7760 29978 7772
rect 36446 7760 36452 7772
rect 36504 7760 36510 7812
rect 11790 7692 11796 7744
rect 11848 7732 11854 7744
rect 17494 7732 17500 7744
rect 11848 7704 17500 7732
rect 11848 7692 11854 7704
rect 17494 7692 17500 7704
rect 17552 7692 17558 7744
rect 21450 7692 21456 7744
rect 21508 7732 21514 7744
rect 21508 7704 23520 7732
rect 21508 7692 21514 7704
rect 12894 7624 12900 7676
rect 12952 7664 12958 7676
rect 13354 7664 13360 7676
rect 12952 7636 13360 7664
rect 12952 7624 12958 7636
rect 13354 7624 13360 7636
rect 13412 7624 13418 7676
rect 13446 7624 13452 7676
rect 13504 7664 13510 7676
rect 15930 7664 15936 7676
rect 13504 7636 15936 7664
rect 13504 7624 13510 7636
rect 15930 7624 15936 7636
rect 15988 7624 15994 7676
rect 16298 7624 16304 7676
rect 16356 7664 16362 7676
rect 16356 7636 21634 7664
rect 16356 7624 16362 7636
rect 21606 7608 21634 7636
rect 14596 7596 14602 7608
rect 11716 7568 14602 7596
rect 14596 7556 14602 7568
rect 14654 7556 14660 7608
rect 16620 7596 16626 7608
rect 15304 7568 16626 7596
rect 4522 7488 4528 7540
rect 4580 7528 4586 7540
rect 4617 7531 4675 7537
rect 4617 7528 4629 7531
rect 4580 7500 4629 7528
rect 4580 7488 4586 7500
rect 4617 7497 4629 7500
rect 4663 7528 4675 7531
rect 5718 7528 5724 7540
rect 4663 7500 5724 7528
rect 4663 7497 4675 7500
rect 4617 7491 4675 7497
rect 5718 7488 5724 7500
rect 5776 7488 5782 7540
rect 5905 7531 5963 7537
rect 5905 7497 5917 7531
rect 5951 7528 5963 7531
rect 5994 7528 6000 7540
rect 5951 7500 6000 7528
rect 5951 7497 5963 7500
rect 5905 7491 5963 7497
rect 5994 7488 6000 7500
rect 6052 7528 6058 7540
rect 6730 7528 6736 7540
rect 6052 7500 6736 7528
rect 6052 7488 6058 7500
rect 6730 7488 6736 7500
rect 6788 7488 6794 7540
rect 7374 7528 7380 7540
rect 6932 7500 7380 7528
rect 6362 7460 6368 7472
rect 3712 7432 6368 7460
rect 3712 7401 3740 7432
rect 6362 7420 6368 7432
rect 6420 7420 6426 7472
rect 3697 7395 3755 7401
rect 3697 7361 3709 7395
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 4246 7352 4252 7404
rect 4304 7352 4310 7404
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5534 7352 5540 7404
rect 5592 7352 5598 7404
rect 5718 7352 5724 7404
rect 5776 7392 5782 7404
rect 5776 7364 6408 7392
rect 5776 7352 5782 7364
rect 3789 7327 3847 7333
rect 3789 7293 3801 7327
rect 3835 7293 3847 7327
rect 3789 7287 3847 7293
rect 3804 7256 3832 7287
rect 4154 7284 4160 7336
rect 4212 7324 4218 7336
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 4212 7296 4813 7324
rect 4212 7284 4218 7296
rect 4801 7293 4813 7296
rect 4847 7293 4859 7327
rect 4801 7287 4859 7293
rect 5077 7327 5135 7333
rect 5077 7293 5089 7327
rect 5123 7293 5135 7327
rect 5442 7324 5448 7336
rect 5077 7287 5135 7293
rect 5368 7296 5448 7324
rect 3528 7228 3832 7256
rect 3050 7148 3056 7200
rect 3108 7188 3114 7200
rect 3528 7197 3556 7228
rect 4614 7216 4620 7268
rect 4672 7256 4678 7268
rect 5092 7256 5120 7287
rect 4672 7228 5120 7256
rect 4672 7216 4678 7228
rect 3513 7191 3571 7197
rect 3513 7188 3525 7191
rect 3108 7160 3525 7188
rect 3108 7148 3114 7160
rect 3513 7157 3525 7160
rect 3559 7157 3571 7191
rect 3513 7151 3571 7157
rect 4430 7148 4436 7200
rect 4488 7188 4494 7200
rect 5368 7188 5396 7296
rect 5442 7284 5448 7296
rect 5500 7324 5506 7336
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5500 7296 6101 7324
rect 5500 7284 5506 7296
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 6089 7287 6147 7293
rect 6181 7327 6239 7333
rect 6181 7293 6193 7327
rect 6227 7293 6239 7327
rect 6181 7287 6239 7293
rect 4488 7160 5396 7188
rect 6196 7188 6224 7287
rect 6270 7284 6276 7336
rect 6328 7284 6334 7336
rect 6380 7333 6408 7364
rect 6546 7352 6552 7404
rect 6604 7392 6610 7404
rect 6825 7395 6883 7401
rect 6825 7392 6837 7395
rect 6604 7364 6837 7392
rect 6604 7352 6610 7364
rect 6825 7361 6837 7364
rect 6871 7361 6883 7395
rect 6825 7355 6883 7361
rect 6932 7333 6960 7500
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 8573 7531 8631 7537
rect 8573 7497 8585 7531
rect 8619 7528 8631 7531
rect 8941 7531 8999 7537
rect 8941 7528 8953 7531
rect 8619 7500 8953 7528
rect 8619 7497 8631 7500
rect 8573 7491 8631 7497
rect 8941 7497 8953 7500
rect 8987 7528 8999 7531
rect 9122 7528 9128 7540
rect 8987 7500 9128 7528
rect 8987 7497 8999 7500
rect 8941 7491 8999 7497
rect 9122 7488 9128 7500
rect 9180 7488 9186 7540
rect 10965 7531 11023 7537
rect 9784 7500 10180 7528
rect 9784 7460 9812 7500
rect 10042 7460 10048 7472
rect 7576 7432 9812 7460
rect 9876 7432 10048 7460
rect 7466 7352 7472 7404
rect 7524 7352 7530 7404
rect 7576 7401 7604 7432
rect 7561 7395 7619 7401
rect 7561 7361 7573 7395
rect 7607 7361 7619 7395
rect 7561 7355 7619 7361
rect 8113 7395 8171 7401
rect 8113 7361 8125 7395
rect 8159 7392 8171 7395
rect 8662 7392 8668 7404
rect 8159 7364 8668 7392
rect 8159 7361 8171 7364
rect 8113 7355 8171 7361
rect 8662 7352 8668 7364
rect 8720 7352 8726 7404
rect 9876 7401 9904 7432
rect 10042 7420 10048 7432
rect 10100 7420 10106 7472
rect 10152 7460 10180 7500
rect 10965 7497 10977 7531
rect 11011 7528 11023 7531
rect 11146 7528 11152 7540
rect 11011 7500 11152 7528
rect 11011 7497 11023 7500
rect 10965 7491 11023 7497
rect 11146 7488 11152 7500
rect 11204 7488 11210 7540
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 15148 7528 15154 7540
rect 12400 7500 15154 7528
rect 12400 7488 12406 7500
rect 15148 7488 15154 7500
rect 15206 7488 15212 7540
rect 13446 7460 13452 7472
rect 10152 7432 13452 7460
rect 13446 7420 13452 7432
rect 13504 7420 13510 7472
rect 9217 7395 9275 7401
rect 9217 7361 9229 7395
rect 9263 7392 9275 7395
rect 9861 7395 9919 7401
rect 9263 7364 9812 7392
rect 9263 7361 9275 7364
rect 9217 7355 9275 7361
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7293 6423 7327
rect 6365 7287 6423 7293
rect 6917 7327 6975 7333
rect 6917 7293 6929 7327
rect 6963 7293 6975 7327
rect 6917 7287 6975 7293
rect 7009 7327 7067 7333
rect 7009 7293 7021 7327
rect 7055 7293 7067 7327
rect 7009 7287 7067 7293
rect 6454 7216 6460 7268
rect 6512 7256 6518 7268
rect 7024 7256 7052 7287
rect 7374 7284 7380 7336
rect 7432 7324 7438 7336
rect 7653 7327 7711 7333
rect 7653 7324 7665 7327
rect 7432 7296 7665 7324
rect 7432 7284 7438 7296
rect 7653 7293 7665 7296
rect 7699 7293 7711 7327
rect 7653 7287 7711 7293
rect 8202 7284 8208 7336
rect 8260 7324 8266 7336
rect 9125 7327 9183 7333
rect 9125 7324 9137 7327
rect 8260 7296 9137 7324
rect 8260 7284 8266 7296
rect 9125 7293 9137 7296
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9306 7284 9312 7336
rect 9364 7284 9370 7336
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7293 9459 7327
rect 9401 7287 9459 7293
rect 9416 7256 9444 7287
rect 6512 7228 7052 7256
rect 8312 7228 9444 7256
rect 9784 7256 9812 7364
rect 9861 7361 9873 7395
rect 9907 7361 9919 7395
rect 9861 7355 9919 7361
rect 9953 7395 10011 7401
rect 9953 7361 9965 7395
rect 9999 7392 10011 7395
rect 10686 7392 10692 7404
rect 9999 7364 10692 7392
rect 9999 7361 10011 7364
rect 9953 7355 10011 7361
rect 10686 7352 10692 7364
rect 10744 7352 10750 7404
rect 11241 7395 11299 7401
rect 11241 7361 11253 7395
rect 11287 7392 11299 7395
rect 13538 7392 13544 7404
rect 11287 7364 13544 7392
rect 11287 7361 11299 7364
rect 11241 7355 11299 7361
rect 13538 7352 13544 7364
rect 13596 7352 13602 7404
rect 10045 7327 10103 7333
rect 10045 7293 10057 7327
rect 10091 7324 10103 7327
rect 10134 7324 10140 7336
rect 10091 7296 10140 7324
rect 10091 7293 10103 7296
rect 10045 7287 10103 7293
rect 10134 7284 10140 7296
rect 10192 7284 10198 7336
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 10962 7324 10968 7336
rect 10551 7296 10968 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 10962 7284 10968 7296
rect 11020 7284 11026 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 11149 7327 11207 7333
rect 11149 7324 11161 7327
rect 11112 7296 11161 7324
rect 11112 7284 11118 7296
rect 11149 7293 11161 7296
rect 11195 7293 11207 7327
rect 11149 7287 11207 7293
rect 15304 7256 15332 7568
rect 16620 7556 16626 7568
rect 16678 7556 16684 7608
rect 19748 7596 19754 7608
rect 16776 7568 19754 7596
rect 15562 7488 15568 7540
rect 15620 7528 15626 7540
rect 16776 7528 16804 7568
rect 19748 7556 19754 7568
rect 19806 7556 19812 7608
rect 21588 7556 21594 7608
rect 21646 7556 21652 7608
rect 23492 7596 23520 7704
rect 23566 7692 23572 7744
rect 23624 7692 23630 7744
rect 29546 7692 29552 7744
rect 29604 7732 29610 7744
rect 36170 7732 36176 7744
rect 29604 7704 36176 7732
rect 29604 7692 29610 7704
rect 36170 7692 36176 7704
rect 36228 7692 36234 7744
rect 32476 7642 43516 7664
rect 23796 7596 23802 7608
rect 23492 7568 23802 7596
rect 23796 7556 23802 7568
rect 23854 7556 23860 7608
rect 24946 7556 24952 7608
rect 25004 7596 25010 7608
rect 25820 7596 25826 7608
rect 25004 7568 25826 7596
rect 25004 7556 25010 7568
rect 25820 7556 25826 7568
rect 25878 7556 25884 7608
rect 28396 7556 28402 7608
rect 28454 7596 28460 7608
rect 30834 7596 30840 7608
rect 28454 7568 30840 7596
rect 28454 7556 28460 7568
rect 30834 7556 30840 7568
rect 30892 7556 30898 7608
rect 32476 7590 41306 7642
rect 41358 7590 41370 7642
rect 41422 7590 41434 7642
rect 41486 7590 41498 7642
rect 41550 7590 41562 7642
rect 41614 7590 43516 7642
rect 32476 7568 43516 7590
rect 15620 7500 16804 7528
rect 15620 7488 15626 7500
rect 17724 7488 17730 7540
rect 17782 7488 17788 7540
rect 17954 7488 17960 7540
rect 18012 7528 18018 7540
rect 18012 7500 19334 7528
rect 18012 7488 18018 7500
rect 17742 7460 17770 7488
rect 9784 7228 15332 7256
rect 15396 7432 17770 7460
rect 19306 7460 19334 7500
rect 20116 7488 20122 7540
rect 20174 7488 20180 7540
rect 22002 7488 22008 7540
rect 22060 7528 22066 7540
rect 25268 7528 25274 7540
rect 22060 7500 25274 7528
rect 22060 7488 22066 7500
rect 25268 7488 25274 7500
rect 25326 7488 25332 7540
rect 27292 7488 27298 7540
rect 27350 7488 27356 7540
rect 28948 7488 28954 7540
rect 29006 7528 29012 7540
rect 36354 7528 36360 7540
rect 29006 7500 36360 7528
rect 29006 7488 29012 7500
rect 36354 7488 36360 7500
rect 36412 7488 36418 7540
rect 20134 7460 20162 7488
rect 19306 7432 20162 7460
rect 6512 7216 6518 7228
rect 8312 7200 8340 7228
rect 8110 7188 8116 7200
rect 6196 7160 8116 7188
rect 4488 7148 4494 7160
rect 8110 7148 8116 7160
rect 8168 7148 8174 7200
rect 8294 7148 8300 7200
rect 8352 7148 8358 7200
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 10134 7188 10140 7200
rect 9088 7160 10140 7188
rect 9088 7148 9094 7160
rect 10134 7148 10140 7160
rect 10192 7148 10198 7200
rect 10686 7148 10692 7200
rect 10744 7188 10750 7200
rect 15396 7188 15424 7432
rect 27310 7392 27338 7488
rect 32769 7395 32827 7401
rect 32769 7392 32781 7395
rect 27310 7364 32781 7392
rect 32769 7361 32781 7364
rect 32815 7361 32827 7395
rect 32769 7355 32827 7361
rect 33318 7352 33324 7404
rect 33376 7352 33382 7404
rect 32306 7284 32312 7336
rect 32364 7324 32370 7336
rect 32861 7327 32919 7333
rect 32861 7324 32873 7327
rect 32364 7296 32873 7324
rect 32364 7284 32370 7296
rect 32861 7293 32873 7296
rect 32907 7324 32919 7327
rect 33413 7327 33471 7333
rect 33413 7324 33425 7327
rect 32907 7296 33425 7324
rect 32907 7293 32919 7296
rect 32861 7287 32919 7293
rect 33413 7293 33425 7296
rect 33459 7293 33471 7327
rect 33413 7287 33471 7293
rect 10744 7160 15424 7188
rect 10744 7148 10750 7160
rect 37642 7148 37648 7200
rect 37700 7188 37706 7200
rect 38378 7188 38384 7200
rect 37700 7160 38384 7188
rect 37700 7148 37706 7160
rect 38378 7148 38384 7160
rect 38436 7148 38442 7200
rect 460 7098 11592 7120
rect 460 7046 1946 7098
rect 1998 7046 2010 7098
rect 2062 7046 2074 7098
rect 2126 7046 2138 7098
rect 2190 7046 2202 7098
rect 2254 7046 9946 7098
rect 9998 7046 10010 7098
rect 10062 7046 10074 7098
rect 10126 7046 10138 7098
rect 10190 7046 10202 7098
rect 10254 7046 11592 7098
rect 460 7024 11592 7046
rect 32476 7098 43516 7120
rect 32476 7046 33946 7098
rect 33998 7046 34010 7098
rect 34062 7046 34074 7098
rect 34126 7046 34138 7098
rect 34190 7046 34202 7098
rect 34254 7046 41946 7098
rect 41998 7046 42010 7098
rect 42062 7046 42074 7098
rect 42126 7046 42138 7098
rect 42190 7046 42202 7098
rect 42254 7046 43516 7098
rect 32476 7024 43516 7046
rect 4522 6944 4528 6996
rect 4580 6944 4586 6996
rect 5994 6944 6000 6996
rect 6052 6944 6058 6996
rect 6270 6944 6276 6996
rect 6328 6984 6334 6996
rect 12342 6984 12348 6996
rect 6328 6956 12348 6984
rect 6328 6944 6334 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 9306 6876 9312 6928
rect 9364 6916 9370 6928
rect 11238 6916 11244 6928
rect 9364 6888 11244 6916
rect 9364 6876 9370 6888
rect 11238 6876 11244 6888
rect 11296 6876 11302 6928
rect 12894 6916 12900 6928
rect 12406 6888 12900 6916
rect 4985 6851 5043 6857
rect 4985 6817 4997 6851
rect 5031 6817 5043 6851
rect 4985 6811 5043 6817
rect 5445 6851 5503 6857
rect 5445 6817 5457 6851
rect 5491 6848 5503 6851
rect 5626 6848 5632 6860
rect 5491 6820 5632 6848
rect 5491 6817 5503 6820
rect 5445 6811 5503 6817
rect 3878 6740 3884 6792
rect 3936 6780 3942 6792
rect 4341 6783 4399 6789
rect 4341 6780 4353 6783
rect 3936 6752 4353 6780
rect 3936 6740 3942 6752
rect 4341 6749 4353 6752
rect 4387 6780 4399 6783
rect 4614 6780 4620 6792
rect 4387 6752 4620 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4614 6740 4620 6752
rect 4672 6740 4678 6792
rect 4890 6740 4896 6792
rect 4948 6740 4954 6792
rect 3326 6672 3332 6724
rect 3384 6712 3390 6724
rect 4709 6715 4767 6721
rect 4709 6712 4721 6715
rect 3384 6684 4721 6712
rect 3384 6672 3390 6684
rect 4709 6681 4721 6684
rect 4755 6712 4767 6715
rect 5000 6712 5028 6811
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 6365 6851 6423 6857
rect 6365 6817 6377 6851
rect 6411 6817 6423 6851
rect 6365 6811 6423 6817
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 7006 6848 7012 6860
rect 6871 6820 7012 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5718 6780 5724 6792
rect 5132 6752 5724 6780
rect 5132 6740 5138 6752
rect 5718 6740 5724 6752
rect 5776 6740 5782 6792
rect 6270 6740 6276 6792
rect 6328 6740 6334 6792
rect 6089 6715 6147 6721
rect 6089 6712 6101 6715
rect 4755 6684 5028 6712
rect 5644 6684 6101 6712
rect 4755 6681 4767 6684
rect 4709 6675 4767 6681
rect 3602 6604 3608 6656
rect 3660 6644 3666 6656
rect 4154 6644 4160 6656
rect 3660 6616 4160 6644
rect 3660 6604 3666 6616
rect 4154 6604 4160 6616
rect 4212 6604 4218 6656
rect 4798 6604 4804 6656
rect 4856 6644 4862 6656
rect 5644 6644 5672 6684
rect 6089 6681 6101 6684
rect 6135 6712 6147 6715
rect 6380 6712 6408 6811
rect 7006 6808 7012 6820
rect 7064 6808 7070 6860
rect 7193 6851 7251 6857
rect 7193 6817 7205 6851
rect 7239 6817 7251 6851
rect 7193 6811 7251 6817
rect 7653 6851 7711 6857
rect 7653 6817 7665 6851
rect 7699 6848 7711 6851
rect 7834 6848 7840 6860
rect 7699 6820 7840 6848
rect 7699 6817 7711 6820
rect 7653 6811 7711 6817
rect 7098 6740 7104 6792
rect 7156 6740 7162 6792
rect 6135 6684 6408 6712
rect 6135 6681 6147 6684
rect 6089 6675 6147 6681
rect 6822 6672 6828 6724
rect 6880 6712 6886 6724
rect 7208 6712 7236 6811
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 8665 6851 8723 6857
rect 8665 6817 8677 6851
rect 8711 6817 8723 6851
rect 8665 6811 8723 6817
rect 8680 6780 8708 6811
rect 8754 6808 8760 6860
rect 8812 6808 8818 6860
rect 8941 6851 8999 6857
rect 8941 6817 8953 6851
rect 8987 6817 8999 6851
rect 8941 6811 8999 6817
rect 6880 6684 7236 6712
rect 7668 6752 8708 6780
rect 6880 6672 6886 6684
rect 4856 6616 5672 6644
rect 4856 6604 4862 6616
rect 6638 6604 6644 6656
rect 6696 6644 6702 6656
rect 7668 6644 7696 6752
rect 8846 6740 8852 6792
rect 8904 6740 8910 6792
rect 7742 6672 7748 6724
rect 7800 6712 7806 6724
rect 8956 6712 8984 6811
rect 9490 6808 9496 6860
rect 9548 6808 9554 6860
rect 9585 6851 9643 6857
rect 9585 6817 9597 6851
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9600 6780 9628 6811
rect 9950 6808 9956 6860
rect 10008 6848 10014 6860
rect 10249 6851 10307 6857
rect 10249 6848 10261 6851
rect 10008 6820 10261 6848
rect 10008 6808 10014 6820
rect 10249 6817 10261 6820
rect 10295 6817 10307 6851
rect 10249 6811 10307 6817
rect 11146 6808 11152 6860
rect 11204 6848 11210 6860
rect 12406 6848 12434 6888
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 36078 6876 36084 6928
rect 36136 6916 36142 6928
rect 36446 6916 36452 6928
rect 36136 6888 36452 6916
rect 36136 6876 36142 6888
rect 36446 6876 36452 6888
rect 36504 6876 36510 6928
rect 11204 6820 12434 6848
rect 11204 6808 11210 6820
rect 32858 6808 32864 6860
rect 32916 6808 32922 6860
rect 32953 6851 33011 6857
rect 32953 6817 32965 6851
rect 32999 6817 33011 6851
rect 32953 6811 33011 6817
rect 33413 6851 33471 6857
rect 33413 6817 33425 6851
rect 33459 6848 33471 6851
rect 33965 6851 34023 6857
rect 33965 6848 33977 6851
rect 33459 6820 33977 6848
rect 33459 6817 33471 6820
rect 33413 6811 33471 6817
rect 33965 6817 33977 6820
rect 34011 6817 34023 6851
rect 33965 6811 34023 6817
rect 9180 6752 9628 6780
rect 10045 6783 10103 6789
rect 9180 6740 9186 6752
rect 10045 6749 10057 6783
rect 10091 6749 10103 6783
rect 10045 6743 10103 6749
rect 7800 6684 8984 6712
rect 10060 6712 10088 6743
rect 10134 6740 10140 6792
rect 10192 6740 10198 6792
rect 10689 6783 10747 6789
rect 10689 6749 10701 6783
rect 10735 6780 10747 6783
rect 10965 6783 11023 6789
rect 10965 6780 10977 6783
rect 10735 6752 10977 6780
rect 10735 6749 10747 6752
rect 10689 6743 10747 6749
rect 10965 6749 10977 6752
rect 11011 6780 11023 6783
rect 11698 6780 11704 6792
rect 11011 6752 11704 6780
rect 11011 6749 11023 6752
rect 10965 6743 11023 6749
rect 11698 6740 11704 6752
rect 11756 6740 11762 6792
rect 32490 6740 32496 6792
rect 32548 6780 32554 6792
rect 32968 6780 32996 6811
rect 34606 6808 34612 6860
rect 34664 6848 34670 6860
rect 34793 6851 34851 6857
rect 34793 6848 34805 6851
rect 34664 6820 34805 6848
rect 34664 6808 34670 6820
rect 34793 6817 34805 6820
rect 34839 6817 34851 6851
rect 34793 6811 34851 6817
rect 33505 6783 33563 6789
rect 33505 6780 33517 6783
rect 32548 6752 33517 6780
rect 32548 6740 32554 6752
rect 33505 6749 33517 6752
rect 33551 6749 33563 6783
rect 33505 6743 33563 6749
rect 34333 6783 34391 6789
rect 34333 6749 34345 6783
rect 34379 6780 34391 6783
rect 35618 6780 35624 6792
rect 34379 6752 35624 6780
rect 34379 6749 34391 6752
rect 34333 6743 34391 6749
rect 35618 6740 35624 6752
rect 35676 6740 35682 6792
rect 10410 6712 10416 6724
rect 10060 6684 10416 6712
rect 7800 6672 7806 6684
rect 10410 6672 10416 6684
rect 10468 6672 10474 6724
rect 7837 6647 7895 6653
rect 7837 6644 7849 6647
rect 6696 6616 7849 6644
rect 6696 6604 6702 6616
rect 7837 6613 7849 6616
rect 7883 6613 7895 6647
rect 7837 6607 7895 6613
rect 8113 6647 8171 6653
rect 8113 6613 8125 6647
rect 8159 6644 8171 6647
rect 8481 6647 8539 6653
rect 8481 6644 8493 6647
rect 8159 6616 8493 6644
rect 8159 6613 8171 6616
rect 8113 6607 8171 6613
rect 8481 6613 8493 6616
rect 8527 6644 8539 6647
rect 8938 6644 8944 6656
rect 8527 6616 8944 6644
rect 8527 6613 8539 6616
rect 8481 6607 8539 6613
rect 8938 6604 8944 6616
rect 8996 6604 9002 6656
rect 9125 6647 9183 6653
rect 9125 6613 9137 6647
rect 9171 6644 9183 6647
rect 9858 6644 9864 6656
rect 9171 6616 9864 6644
rect 9171 6613 9183 6616
rect 9125 6607 9183 6613
rect 9858 6604 9864 6616
rect 9916 6644 9922 6656
rect 10502 6644 10508 6656
rect 9916 6616 10508 6644
rect 9916 6604 9922 6616
rect 10502 6604 10508 6616
rect 10560 6604 10566 6656
rect 13078 6644 13084 6656
rect 11624 6616 13084 6644
rect 460 6554 11592 6576
rect 460 6502 1306 6554
rect 1358 6502 1370 6554
rect 1422 6502 1434 6554
rect 1486 6502 1498 6554
rect 1550 6502 1562 6554
rect 1614 6502 9306 6554
rect 9358 6502 9370 6554
rect 9422 6502 9434 6554
rect 9486 6502 9498 6554
rect 9550 6502 9562 6554
rect 9614 6502 11592 6554
rect 460 6480 11592 6502
rect 5626 6400 5632 6452
rect 5684 6400 5690 6452
rect 7834 6400 7840 6452
rect 7892 6400 7898 6452
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 8662 6440 8668 6452
rect 8435 6412 8668 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8662 6400 8668 6412
rect 8720 6400 8726 6452
rect 8846 6400 8852 6452
rect 8904 6440 8910 6452
rect 11330 6440 11336 6452
rect 8904 6412 11336 6440
rect 8904 6400 8910 6412
rect 11330 6400 11336 6412
rect 11388 6400 11394 6452
rect 9766 6372 9772 6384
rect 9508 6344 9772 6372
rect 9508 6313 9536 6344
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 10502 6372 10508 6384
rect 10336 6344 10508 6372
rect 10336 6313 10364 6344
rect 10502 6332 10508 6344
rect 10560 6372 10566 6384
rect 10778 6372 10784 6384
rect 10560 6344 10784 6372
rect 10560 6332 10566 6344
rect 10778 6332 10784 6344
rect 10836 6332 10842 6384
rect 11514 6372 11520 6384
rect 11164 6344 11520 6372
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 10321 6307 10379 6313
rect 9493 6267 9551 6273
rect 9784 6276 10272 6304
rect 8938 6196 8944 6248
rect 8996 6196 9002 6248
rect 9784 6245 9812 6276
rect 9033 6239 9091 6245
rect 9033 6205 9045 6239
rect 9079 6205 9091 6239
rect 9033 6199 9091 6205
rect 9769 6239 9827 6245
rect 9769 6205 9781 6239
rect 9815 6205 9827 6239
rect 9769 6199 9827 6205
rect 9861 6239 9919 6245
rect 9861 6205 9873 6239
rect 9907 6205 9919 6239
rect 9861 6199 9919 6205
rect 6362 6128 6368 6180
rect 6420 6168 6426 6180
rect 7374 6168 7380 6180
rect 6420 6140 7380 6168
rect 6420 6128 6426 6140
rect 7374 6128 7380 6140
rect 7432 6128 7438 6180
rect 7466 6128 7472 6180
rect 7524 6168 7530 6180
rect 8481 6171 8539 6177
rect 8481 6168 8493 6171
rect 7524 6140 8493 6168
rect 7524 6128 7530 6140
rect 8481 6137 8493 6140
rect 8527 6168 8539 6171
rect 9048 6168 9076 6199
rect 8527 6140 9076 6168
rect 8527 6137 8539 6140
rect 8481 6131 8539 6137
rect 9582 6128 9588 6180
rect 9640 6168 9646 6180
rect 9876 6168 9904 6199
rect 9640 6140 9904 6168
rect 9640 6128 9646 6140
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6822 6100 6828 6112
rect 5592 6072 6828 6100
rect 5592 6060 5598 6072
rect 6822 6060 6828 6072
rect 6880 6100 6886 6112
rect 6917 6103 6975 6109
rect 6917 6100 6929 6103
rect 6880 6072 6929 6100
rect 6880 6060 6886 6072
rect 6917 6069 6929 6072
rect 6963 6069 6975 6103
rect 6917 6063 6975 6069
rect 7742 6060 7748 6112
rect 7800 6100 7806 6112
rect 8665 6103 8723 6109
rect 8665 6100 8677 6103
rect 7800 6072 8677 6100
rect 7800 6060 7806 6072
rect 8665 6069 8677 6072
rect 8711 6069 8723 6103
rect 8665 6063 8723 6069
rect 9214 6060 9220 6112
rect 9272 6100 9278 6112
rect 9677 6103 9735 6109
rect 9677 6100 9689 6103
rect 9272 6072 9689 6100
rect 9272 6060 9278 6072
rect 9677 6069 9689 6072
rect 9723 6100 9735 6103
rect 9950 6100 9956 6112
rect 9723 6072 9956 6100
rect 9723 6069 9735 6072
rect 9677 6063 9735 6069
rect 9950 6060 9956 6072
rect 10008 6060 10014 6112
rect 10244 6100 10272 6276
rect 10321 6273 10333 6307
rect 10367 6273 10379 6307
rect 10321 6267 10379 6273
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6304 10747 6307
rect 11164 6304 11192 6344
rect 11514 6332 11520 6344
rect 11572 6332 11578 6384
rect 10735 6276 11192 6304
rect 11241 6307 11299 6313
rect 10735 6273 10747 6276
rect 10689 6267 10747 6273
rect 11241 6273 11253 6307
rect 11287 6304 11299 6307
rect 11624 6304 11652 6616
rect 13078 6604 13084 6616
rect 13136 6604 13142 6656
rect 31478 6604 31484 6656
rect 31536 6644 31542 6656
rect 31536 6616 32444 6644
rect 31536 6604 31542 6616
rect 32416 6440 32444 6616
rect 32476 6554 43516 6576
rect 32476 6502 41306 6554
rect 41358 6502 41370 6554
rect 41422 6502 41434 6554
rect 41486 6502 41498 6554
rect 41550 6502 41562 6554
rect 41614 6502 43516 6554
rect 32476 6480 43516 6502
rect 32416 6412 33088 6440
rect 33060 6313 33088 6412
rect 37918 6400 37924 6452
rect 37976 6440 37982 6452
rect 39850 6440 39856 6452
rect 37976 6412 39856 6440
rect 37976 6400 37982 6412
rect 39850 6400 39856 6412
rect 39908 6400 39914 6452
rect 11287 6276 11652 6304
rect 11287 6273 11299 6276
rect 11241 6267 11299 6273
rect 10778 6196 10784 6248
rect 10836 6196 10842 6248
rect 10597 6171 10655 6177
rect 10597 6137 10609 6171
rect 10643 6168 10655 6171
rect 10796 6168 10824 6196
rect 10643 6140 10824 6168
rect 10643 6137 10655 6140
rect 10597 6131 10655 6137
rect 11514 6100 11520 6112
rect 10244 6072 11520 6100
rect 11514 6060 11520 6072
rect 11572 6060 11578 6112
rect 460 6010 11592 6032
rect 460 5958 1946 6010
rect 1998 5958 2010 6010
rect 2062 5958 2074 6010
rect 2126 5958 2138 6010
rect 2190 5958 2202 6010
rect 2254 5958 9946 6010
rect 9998 5958 10010 6010
rect 10062 5958 10074 6010
rect 10126 5958 10138 6010
rect 10190 5958 10202 6010
rect 10254 5958 11592 6010
rect 460 5936 11592 5958
rect 9766 5856 9772 5908
rect 9824 5856 9830 5908
rect 10229 5899 10287 5905
rect 10229 5865 10241 5899
rect 10275 5896 10287 5899
rect 10410 5896 10416 5908
rect 10275 5868 10416 5896
rect 10275 5865 10287 5868
rect 10229 5859 10287 5865
rect 10410 5856 10416 5868
rect 10468 5856 10474 5908
rect 10502 5856 10508 5908
rect 10560 5856 10566 5908
rect 11241 5899 11299 5905
rect 11241 5865 11253 5899
rect 11287 5896 11299 5899
rect 11624 5896 11652 6276
rect 33045 6307 33103 6313
rect 33045 6273 33057 6307
rect 33091 6273 33103 6307
rect 33045 6267 33103 6273
rect 34609 6307 34667 6313
rect 34609 6273 34621 6307
rect 34655 6304 34667 6307
rect 35986 6304 35992 6316
rect 34655 6276 35992 6304
rect 34655 6273 34667 6276
rect 34609 6267 34667 6273
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 33137 6239 33195 6245
rect 33137 6236 33149 6239
rect 32876 6208 33149 6236
rect 32876 6112 32904 6208
rect 33137 6205 33149 6208
rect 33183 6205 33195 6239
rect 33137 6199 33195 6205
rect 33597 6239 33655 6245
rect 33597 6205 33609 6239
rect 33643 6236 33655 6239
rect 34241 6239 34299 6245
rect 34241 6236 34253 6239
rect 33643 6208 34253 6236
rect 33643 6205 33655 6208
rect 33597 6199 33655 6205
rect 34241 6205 34253 6208
rect 34287 6205 34299 6239
rect 34241 6199 34299 6205
rect 34882 6196 34888 6248
rect 34940 6236 34946 6248
rect 35161 6239 35219 6245
rect 35161 6236 35173 6239
rect 34940 6208 35173 6236
rect 34940 6196 34946 6208
rect 35161 6205 35173 6208
rect 35207 6205 35219 6239
rect 35161 6199 35219 6205
rect 35618 6196 35624 6248
rect 35676 6196 35682 6248
rect 32858 6060 32864 6112
rect 32916 6060 32922 6112
rect 35713 6103 35771 6109
rect 35713 6069 35725 6103
rect 35759 6100 35771 6103
rect 35989 6103 36047 6109
rect 35989 6100 36001 6103
rect 35759 6072 36001 6100
rect 35759 6069 35771 6072
rect 35713 6063 35771 6069
rect 35989 6069 36001 6072
rect 36035 6100 36047 6103
rect 36998 6100 37004 6112
rect 36035 6072 37004 6100
rect 36035 6069 36047 6072
rect 35989 6063 36047 6069
rect 36998 6060 37004 6072
rect 37056 6060 37062 6112
rect 32476 6010 43516 6032
rect 32476 5958 33946 6010
rect 33998 5958 34010 6010
rect 34062 5958 34074 6010
rect 34126 5958 34138 6010
rect 34190 5958 34202 6010
rect 34254 5958 41946 6010
rect 41998 5958 42010 6010
rect 42062 5958 42074 6010
rect 42126 5958 42138 6010
rect 42190 5958 42202 6010
rect 42254 5958 43516 6010
rect 32476 5936 43516 5958
rect 11287 5868 11652 5896
rect 11287 5865 11299 5868
rect 11241 5859 11299 5865
rect 9585 5831 9643 5837
rect 9585 5797 9597 5831
rect 9631 5828 9643 5831
rect 9858 5828 9864 5840
rect 9631 5800 9864 5828
rect 9631 5797 9643 5800
rect 9585 5791 9643 5797
rect 9858 5788 9864 5800
rect 9916 5788 9922 5840
rect 11330 5788 11336 5840
rect 11388 5828 11394 5840
rect 12066 5828 12072 5840
rect 11388 5800 12072 5828
rect 11388 5788 11394 5800
rect 12066 5788 12072 5800
rect 12124 5788 12130 5840
rect 8938 5720 8944 5772
rect 8996 5760 9002 5772
rect 11882 5760 11888 5772
rect 8996 5732 11888 5760
rect 8996 5720 9002 5732
rect 11882 5720 11888 5732
rect 11940 5720 11946 5772
rect 8570 5584 8576 5636
rect 8628 5624 8634 5636
rect 9582 5624 9588 5636
rect 8628 5596 9588 5624
rect 8628 5584 8634 5596
rect 9582 5584 9588 5596
rect 9640 5624 9646 5636
rect 9861 5627 9919 5633
rect 9861 5624 9873 5627
rect 9640 5596 9873 5624
rect 9640 5584 9646 5596
rect 9861 5593 9873 5596
rect 9907 5593 9919 5627
rect 9861 5587 9919 5593
rect 9122 5516 9128 5568
rect 9180 5556 9186 5568
rect 9309 5559 9367 5565
rect 9309 5556 9321 5559
rect 9180 5528 9321 5556
rect 9180 5516 9186 5528
rect 9309 5525 9321 5528
rect 9355 5525 9367 5559
rect 9309 5519 9367 5525
rect 460 5466 11592 5488
rect 460 5414 1306 5466
rect 1358 5414 1370 5466
rect 1422 5414 1434 5466
rect 1486 5414 1498 5466
rect 1550 5414 1562 5466
rect 1614 5414 9306 5466
rect 9358 5414 9370 5466
rect 9422 5414 9434 5466
rect 9486 5414 9498 5466
rect 9550 5414 9562 5466
rect 9614 5414 11592 5466
rect 460 5392 11592 5414
rect 32476 5466 43516 5488
rect 32476 5414 41306 5466
rect 41358 5414 41370 5466
rect 41422 5414 41434 5466
rect 41486 5414 41498 5466
rect 41550 5414 41562 5466
rect 41614 5414 43516 5466
rect 32476 5392 43516 5414
rect 32122 5176 32128 5228
rect 32180 5216 32186 5228
rect 33137 5219 33195 5225
rect 33137 5216 33149 5219
rect 32180 5188 33149 5216
rect 32180 5176 32186 5188
rect 33137 5185 33149 5188
rect 33183 5185 33195 5219
rect 33137 5179 33195 5185
rect 32582 5108 32588 5160
rect 32640 5148 32646 5160
rect 33321 5151 33379 5157
rect 33321 5148 33333 5151
rect 32640 5120 33333 5148
rect 32640 5108 32646 5120
rect 33321 5117 33333 5120
rect 33367 5117 33379 5151
rect 33321 5111 33379 5117
rect 35986 5108 35992 5160
rect 36044 5108 36050 5160
rect 31938 5040 31944 5092
rect 31996 5080 32002 5092
rect 32953 5083 33011 5089
rect 32953 5080 32965 5083
rect 31996 5052 32965 5080
rect 31996 5040 32002 5052
rect 32953 5049 32965 5052
rect 32999 5049 33011 5083
rect 32953 5043 33011 5049
rect 32769 5015 32827 5021
rect 32769 5012 32781 5015
rect 32232 4984 32781 5012
rect 460 4922 11592 4944
rect 460 4870 1946 4922
rect 1998 4870 2010 4922
rect 2062 4870 2074 4922
rect 2126 4870 2138 4922
rect 2190 4870 2202 4922
rect 2254 4870 11592 4922
rect 460 4848 11592 4870
rect 460 4378 11592 4400
rect 460 4326 1306 4378
rect 1358 4326 1370 4378
rect 1422 4326 1434 4378
rect 1486 4326 1498 4378
rect 1550 4326 1562 4378
rect 1614 4326 9306 4378
rect 9358 4326 9370 4378
rect 9422 4326 9434 4378
rect 9486 4326 9498 4378
rect 9550 4326 9562 4378
rect 9614 4326 11592 4378
rect 29914 4360 29920 4412
rect 29972 4400 29978 4412
rect 32232 4400 32260 4984
rect 32769 4981 32781 4984
rect 32815 4981 32827 5015
rect 32769 4975 32827 4981
rect 33686 4972 33692 5024
rect 33744 5012 33750 5024
rect 33965 5015 34023 5021
rect 33965 5012 33977 5015
rect 33744 4984 33977 5012
rect 33744 4972 33750 4984
rect 33965 4981 33977 4984
rect 34011 4981 34023 5015
rect 33965 4975 34023 4981
rect 36081 5015 36139 5021
rect 36081 4981 36093 5015
rect 36127 5012 36139 5015
rect 36357 5015 36415 5021
rect 36357 5012 36369 5015
rect 36127 4984 36369 5012
rect 36127 4981 36139 4984
rect 36081 4975 36139 4981
rect 36357 4981 36369 4984
rect 36403 5012 36415 5015
rect 37274 5012 37280 5024
rect 36403 4984 37280 5012
rect 36403 4981 36415 4984
rect 36357 4975 36415 4981
rect 37274 4972 37280 4984
rect 37332 4972 37338 5024
rect 32476 4922 43516 4944
rect 32476 4870 33946 4922
rect 33998 4870 34010 4922
rect 34062 4870 34074 4922
rect 34126 4870 34138 4922
rect 34190 4870 34202 4922
rect 34254 4870 41946 4922
rect 41998 4870 42010 4922
rect 42062 4870 42074 4922
rect 42126 4870 42138 4922
rect 42190 4870 42202 4922
rect 42254 4870 43516 4922
rect 32476 4848 43516 4870
rect 32766 4632 32772 4684
rect 32824 4632 32830 4684
rect 32950 4632 32956 4684
rect 33008 4672 33014 4684
rect 33137 4675 33195 4681
rect 33137 4672 33149 4675
rect 33008 4644 33149 4672
rect 33008 4632 33014 4644
rect 33137 4641 33149 4644
rect 33183 4641 33195 4675
rect 33137 4635 33195 4641
rect 33226 4632 33232 4684
rect 33284 4632 33290 4684
rect 33689 4675 33747 4681
rect 33689 4641 33701 4675
rect 33735 4672 33747 4675
rect 34517 4675 34575 4681
rect 34517 4672 34529 4675
rect 33735 4644 34529 4672
rect 33735 4641 33747 4644
rect 33689 4635 33747 4641
rect 34517 4641 34529 4644
rect 34563 4641 34575 4675
rect 34517 4635 34575 4641
rect 35158 4632 35164 4684
rect 35216 4672 35222 4684
rect 35345 4675 35403 4681
rect 35345 4672 35357 4675
rect 35216 4644 35357 4672
rect 35216 4632 35222 4644
rect 35345 4641 35357 4644
rect 35391 4641 35403 4675
rect 35345 4635 35403 4641
rect 33244 4604 33272 4632
rect 33781 4607 33839 4613
rect 33781 4604 33793 4607
rect 33244 4576 33793 4604
rect 33781 4573 33793 4576
rect 33827 4573 33839 4607
rect 33781 4567 33839 4573
rect 34885 4607 34943 4613
rect 34885 4573 34897 4607
rect 34931 4604 34943 4607
rect 35894 4604 35900 4616
rect 34931 4576 35900 4604
rect 34931 4573 34943 4576
rect 34885 4567 34943 4573
rect 35894 4564 35900 4576
rect 35952 4564 35958 4616
rect 32861 4539 32919 4545
rect 32861 4505 32873 4539
rect 32907 4536 32919 4539
rect 32907 4508 34928 4536
rect 32907 4505 32919 4508
rect 32861 4499 32919 4505
rect 34900 4480 34928 4508
rect 32950 4428 32956 4480
rect 33008 4468 33014 4480
rect 33965 4471 34023 4477
rect 33965 4468 33977 4471
rect 33008 4440 33977 4468
rect 33008 4428 33014 4440
rect 33965 4437 33977 4440
rect 34011 4437 34023 4471
rect 33965 4431 34023 4437
rect 34330 4428 34336 4480
rect 34388 4428 34394 4480
rect 34882 4428 34888 4480
rect 34940 4428 34946 4480
rect 35618 4428 35624 4480
rect 35676 4428 35682 4480
rect 29972 4372 32260 4400
rect 32476 4378 43516 4400
rect 29972 4360 29978 4372
rect 460 4304 11592 4326
rect 32476 4326 41306 4378
rect 41358 4326 41370 4378
rect 41422 4326 41434 4378
rect 41486 4326 41498 4378
rect 41550 4326 41562 4378
rect 41614 4326 43516 4378
rect 32476 4304 43516 4326
rect 34333 4267 34391 4273
rect 34333 4264 34345 4267
rect 32968 4236 34345 4264
rect 9858 4156 9864 4208
rect 9916 4196 9922 4208
rect 10870 4196 10876 4208
rect 9916 4168 10876 4196
rect 9916 4156 9922 4168
rect 10870 4156 10876 4168
rect 10928 4156 10934 4208
rect 32858 4088 32864 4140
rect 32916 4128 32922 4140
rect 32968 4128 32996 4236
rect 34333 4233 34345 4236
rect 34379 4233 34391 4267
rect 34333 4227 34391 4233
rect 36078 4224 36084 4276
rect 36136 4264 36142 4276
rect 36906 4264 36912 4276
rect 36136 4236 36912 4264
rect 36136 4224 36142 4236
rect 36906 4224 36912 4236
rect 36964 4264 36970 4276
rect 37093 4267 37151 4273
rect 37093 4264 37105 4267
rect 36964 4236 37105 4264
rect 36964 4224 36970 4236
rect 37093 4233 37105 4236
rect 37139 4233 37151 4267
rect 37093 4227 37151 4233
rect 33042 4156 33048 4208
rect 33100 4156 33106 4208
rect 34514 4156 34520 4208
rect 34572 4156 34578 4208
rect 35989 4199 36047 4205
rect 35989 4165 36001 4199
rect 36035 4196 36047 4199
rect 36035 4168 36308 4196
rect 36035 4165 36047 4168
rect 35989 4159 36047 4165
rect 32916 4100 32996 4128
rect 32916 4088 32922 4100
rect 32674 4020 32680 4072
rect 32732 4060 32738 4072
rect 33060 4069 33088 4156
rect 34885 4131 34943 4137
rect 34885 4128 34897 4131
rect 33704 4100 34897 4128
rect 32769 4063 32827 4069
rect 32769 4060 32781 4063
rect 32732 4032 32781 4060
rect 32732 4020 32738 4032
rect 32769 4029 32781 4032
rect 32815 4029 32827 4063
rect 32769 4023 32827 4029
rect 33045 4063 33103 4069
rect 33045 4029 33057 4063
rect 33091 4029 33103 4063
rect 33045 4023 33103 4029
rect 33410 4020 33416 4072
rect 33468 4020 33474 4072
rect 33502 4020 33508 4072
rect 33560 4060 33566 4072
rect 33704 4060 33732 4100
rect 34885 4097 34897 4100
rect 34931 4097 34943 4131
rect 34885 4091 34943 4097
rect 35342 4088 35348 4140
rect 35400 4128 35406 4140
rect 36173 4131 36231 4137
rect 36173 4128 36185 4131
rect 35400 4100 36185 4128
rect 35400 4088 35406 4100
rect 36173 4097 36185 4100
rect 36219 4097 36231 4131
rect 36280 4128 36308 4168
rect 36449 4131 36507 4137
rect 36449 4128 36461 4131
rect 36280 4100 36461 4128
rect 36173 4091 36231 4097
rect 36449 4097 36461 4100
rect 36495 4128 36507 4131
rect 37918 4128 37924 4140
rect 36495 4100 37924 4128
rect 36495 4097 36507 4100
rect 36449 4091 36507 4097
rect 37918 4088 37924 4100
rect 37976 4088 37982 4140
rect 33560 4032 33732 4060
rect 33560 4020 33566 4032
rect 33778 4020 33784 4072
rect 33836 4060 33842 4072
rect 34057 4063 34115 4069
rect 34057 4060 34069 4063
rect 33836 4032 34069 4060
rect 33836 4020 33842 4032
rect 34057 4029 34069 4032
rect 34103 4029 34115 4063
rect 34057 4023 34115 4029
rect 34422 4020 34428 4072
rect 34480 4060 34486 4072
rect 35621 4063 35679 4069
rect 35621 4060 35633 4063
rect 34480 4032 35633 4060
rect 34480 4020 34486 4032
rect 35621 4029 35633 4032
rect 35667 4029 35679 4063
rect 35621 4023 35679 4029
rect 35894 4020 35900 4072
rect 35952 4020 35958 4072
rect 32861 3995 32919 4001
rect 32861 3961 32873 3995
rect 32907 3992 32919 3995
rect 33870 3992 33876 4004
rect 32907 3964 33876 3992
rect 32907 3961 32919 3964
rect 32861 3955 32919 3961
rect 33870 3952 33876 3964
rect 33928 3952 33934 4004
rect 33965 3995 34023 4001
rect 33965 3961 33977 3995
rect 34011 3992 34023 3995
rect 34790 3992 34796 4004
rect 34011 3964 34796 3992
rect 34011 3961 34023 3964
rect 33965 3955 34023 3961
rect 34790 3952 34796 3964
rect 34848 3952 34854 4004
rect 35802 3952 35808 4004
rect 35860 3992 35866 4004
rect 36541 3995 36599 4001
rect 36541 3992 36553 3995
rect 35860 3964 36553 3992
rect 35860 3952 35866 3964
rect 36541 3961 36553 3964
rect 36587 3961 36599 3995
rect 36541 3955 36599 3961
rect 37001 3995 37059 4001
rect 37001 3961 37013 3995
rect 37047 3992 37059 3995
rect 37734 3992 37740 4004
rect 37047 3964 37740 3992
rect 37047 3961 37059 3964
rect 37001 3955 37059 3961
rect 37734 3952 37740 3964
rect 37792 3952 37798 4004
rect 32030 3884 32036 3936
rect 32088 3924 32094 3936
rect 32674 3924 32680 3936
rect 32088 3896 32680 3924
rect 32088 3884 32094 3896
rect 32674 3884 32680 3896
rect 32732 3884 32738 3936
rect 32950 3884 32956 3936
rect 33008 3924 33014 3936
rect 33137 3927 33195 3933
rect 33137 3924 33149 3927
rect 33008 3896 33149 3924
rect 33008 3884 33014 3896
rect 33137 3893 33149 3896
rect 33183 3893 33195 3927
rect 33137 3887 33195 3893
rect 34149 3927 34207 3933
rect 34149 3893 34161 3927
rect 34195 3924 34207 3927
rect 34606 3924 34612 3936
rect 34195 3896 34612 3924
rect 34195 3893 34207 3896
rect 34149 3887 34207 3893
rect 34606 3884 34612 3896
rect 34664 3884 34670 3936
rect 34698 3884 34704 3936
rect 34756 3884 34762 3936
rect 35158 3884 35164 3936
rect 35216 3884 35222 3936
rect 35434 3884 35440 3936
rect 35492 3884 35498 3936
rect 35894 3884 35900 3936
rect 35952 3924 35958 3936
rect 36354 3924 36360 3936
rect 35952 3896 36360 3924
rect 35952 3884 35958 3896
rect 36354 3884 36360 3896
rect 36412 3884 36418 3936
rect 36722 3884 36728 3936
rect 36780 3884 36786 3936
rect 460 3834 11592 3856
rect 460 3782 1946 3834
rect 1998 3782 2010 3834
rect 2062 3782 2074 3834
rect 2126 3782 2138 3834
rect 2190 3782 2202 3834
rect 2254 3782 9946 3834
rect 9998 3782 10010 3834
rect 10062 3782 10074 3834
rect 10126 3782 10138 3834
rect 10190 3782 10202 3834
rect 10254 3782 11592 3834
rect 28350 3816 28356 3868
rect 28408 3856 28414 3868
rect 31846 3856 31852 3868
rect 28408 3828 31852 3856
rect 28408 3816 28414 3828
rect 31846 3816 31852 3828
rect 31904 3816 31910 3868
rect 32476 3834 43516 3856
rect 460 3760 11592 3782
rect 32476 3782 33946 3834
rect 33998 3782 34010 3834
rect 34062 3782 34074 3834
rect 34126 3782 34138 3834
rect 34190 3782 34202 3834
rect 34254 3782 41946 3834
rect 41998 3782 42010 3834
rect 42062 3782 42074 3834
rect 42126 3782 42138 3834
rect 42190 3782 42202 3834
rect 42254 3782 43516 3834
rect 32476 3760 43516 3782
rect 30466 3680 30472 3732
rect 30524 3720 30530 3732
rect 32858 3720 32864 3732
rect 30524 3692 32864 3720
rect 30524 3680 30530 3692
rect 32858 3680 32864 3692
rect 32916 3680 32922 3732
rect 34333 3723 34391 3729
rect 34072 3692 34284 3720
rect 31294 3612 31300 3664
rect 31352 3652 31358 3664
rect 34072 3652 34100 3692
rect 31352 3624 34100 3652
rect 34256 3652 34284 3692
rect 34333 3689 34345 3723
rect 34379 3720 34391 3723
rect 34379 3692 36492 3720
rect 34379 3689 34391 3692
rect 34333 3683 34391 3689
rect 36464 3664 36492 3692
rect 37090 3680 37096 3732
rect 37148 3720 37154 3732
rect 37921 3723 37979 3729
rect 37921 3720 37933 3723
rect 37148 3692 37933 3720
rect 37148 3680 37154 3692
rect 37921 3689 37933 3692
rect 37967 3689 37979 3723
rect 37921 3683 37979 3689
rect 34698 3652 34704 3664
rect 34256 3624 34704 3652
rect 31352 3612 31358 3624
rect 34698 3612 34704 3624
rect 34756 3612 34762 3664
rect 36446 3612 36452 3664
rect 36504 3612 36510 3664
rect 36817 3655 36875 3661
rect 36817 3621 36829 3655
rect 36863 3652 36875 3655
rect 37826 3652 37832 3664
rect 36863 3624 37832 3652
rect 36863 3621 36875 3624
rect 36817 3615 36875 3621
rect 37826 3612 37832 3624
rect 37884 3612 37890 3664
rect 32950 3544 32956 3596
rect 33008 3544 33014 3596
rect 33594 3544 33600 3596
rect 33652 3584 33658 3596
rect 34054 3584 34060 3596
rect 33652 3556 34060 3584
rect 33652 3544 33658 3556
rect 34054 3544 34060 3556
rect 34112 3544 34118 3596
rect 34146 3544 34152 3596
rect 34204 3584 34210 3596
rect 34241 3587 34299 3593
rect 34241 3584 34253 3587
rect 34204 3556 34253 3584
rect 34204 3544 34210 3556
rect 34241 3553 34253 3556
rect 34287 3553 34299 3587
rect 34241 3547 34299 3553
rect 34517 3587 34575 3593
rect 34517 3553 34529 3587
rect 34563 3553 34575 3587
rect 34517 3547 34575 3553
rect 31110 3476 31116 3528
rect 31168 3516 31174 3528
rect 33965 3519 34023 3525
rect 33965 3516 33977 3519
rect 31168 3488 33977 3516
rect 31168 3476 31174 3488
rect 33965 3485 33977 3488
rect 34011 3516 34023 3519
rect 34330 3516 34336 3528
rect 34011 3488 34336 3516
rect 34011 3485 34023 3488
rect 33965 3479 34023 3485
rect 34330 3476 34336 3488
rect 34388 3476 34394 3528
rect 29822 3408 29828 3460
rect 29880 3448 29886 3460
rect 33778 3448 33784 3460
rect 29880 3420 33784 3448
rect 29880 3408 29886 3420
rect 33778 3408 33784 3420
rect 33836 3408 33842 3460
rect 30374 3340 30380 3392
rect 30432 3380 30438 3392
rect 33318 3380 33324 3392
rect 30432 3352 33324 3380
rect 30432 3340 30438 3352
rect 33318 3340 33324 3352
rect 33376 3340 33382 3392
rect 34054 3340 34060 3392
rect 34112 3380 34118 3392
rect 34532 3380 34560 3547
rect 34790 3544 34796 3596
rect 34848 3544 34854 3596
rect 35342 3544 35348 3596
rect 35400 3544 35406 3596
rect 35434 3544 35440 3596
rect 35492 3584 35498 3596
rect 35713 3587 35771 3593
rect 35713 3584 35725 3587
rect 35492 3556 35725 3584
rect 35492 3544 35498 3556
rect 35713 3553 35725 3556
rect 35759 3553 35771 3587
rect 35713 3547 35771 3553
rect 35802 3544 35808 3596
rect 35860 3584 35866 3596
rect 36357 3587 36415 3593
rect 36357 3584 36369 3587
rect 35860 3556 36369 3584
rect 35860 3544 35866 3556
rect 36357 3553 36369 3556
rect 36403 3553 36415 3587
rect 36357 3547 36415 3553
rect 36538 3544 36544 3596
rect 36596 3584 36602 3596
rect 36909 3587 36967 3593
rect 36909 3584 36921 3587
rect 36596 3556 36921 3584
rect 36596 3544 36602 3556
rect 36909 3553 36921 3556
rect 36955 3553 36967 3587
rect 36909 3547 36967 3553
rect 37001 3587 37059 3593
rect 37001 3553 37013 3587
rect 37047 3553 37059 3587
rect 37001 3547 37059 3553
rect 34606 3476 34612 3528
rect 34664 3516 34670 3528
rect 35526 3516 35532 3528
rect 34664 3488 35532 3516
rect 34664 3476 34670 3488
rect 35526 3476 35532 3488
rect 35584 3476 35590 3528
rect 35621 3519 35679 3525
rect 35621 3485 35633 3519
rect 35667 3485 35679 3519
rect 35621 3479 35679 3485
rect 35250 3408 35256 3460
rect 35308 3448 35314 3460
rect 35636 3448 35664 3479
rect 36078 3476 36084 3528
rect 36136 3516 36142 3528
rect 36265 3519 36323 3525
rect 36265 3516 36277 3519
rect 36136 3488 36277 3516
rect 36136 3476 36142 3488
rect 36265 3485 36277 3488
rect 36311 3485 36323 3519
rect 36265 3479 36323 3485
rect 35308 3420 35664 3448
rect 35308 3408 35314 3420
rect 36170 3408 36176 3460
rect 36228 3448 36234 3460
rect 36722 3448 36728 3460
rect 36228 3420 36728 3448
rect 36228 3408 36234 3420
rect 36722 3408 36728 3420
rect 36780 3448 36786 3460
rect 37016 3448 37044 3547
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 38105 3587 38163 3593
rect 38105 3584 38117 3587
rect 37424 3556 38117 3584
rect 37424 3544 37430 3556
rect 38105 3553 38117 3556
rect 38151 3584 38163 3587
rect 38562 3584 38568 3596
rect 38151 3556 38568 3584
rect 38151 3553 38163 3556
rect 38105 3547 38163 3553
rect 38562 3544 38568 3556
rect 38620 3544 38626 3596
rect 37461 3519 37519 3525
rect 37461 3485 37473 3519
rect 37507 3516 37519 3519
rect 37642 3516 37648 3528
rect 37507 3488 37648 3516
rect 37507 3485 37519 3488
rect 37461 3479 37519 3485
rect 37642 3476 37648 3488
rect 37700 3476 37706 3528
rect 36780 3420 37044 3448
rect 36780 3408 36786 3420
rect 37182 3408 37188 3460
rect 37240 3448 37246 3460
rect 37737 3451 37795 3457
rect 37737 3448 37749 3451
rect 37240 3420 37749 3448
rect 37240 3408 37246 3420
rect 37737 3417 37749 3420
rect 37783 3417 37795 3451
rect 37737 3411 37795 3417
rect 34112 3352 34560 3380
rect 34112 3340 34118 3352
rect 34606 3340 34612 3392
rect 34664 3340 34670 3392
rect 34885 3383 34943 3389
rect 34885 3349 34897 3383
rect 34931 3380 34943 3383
rect 35802 3380 35808 3392
rect 34931 3352 35808 3380
rect 34931 3349 34943 3352
rect 34885 3343 34943 3349
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 35897 3383 35955 3389
rect 35897 3349 35909 3383
rect 35943 3380 35955 3383
rect 37458 3380 37464 3392
rect 35943 3352 37464 3380
rect 35943 3349 35955 3352
rect 35897 3343 35955 3349
rect 37458 3340 37464 3352
rect 37516 3340 37522 3392
rect 460 3290 43516 3312
rect 460 3238 1306 3290
rect 1358 3238 1370 3290
rect 1422 3238 1434 3290
rect 1486 3238 1498 3290
rect 1550 3238 1562 3290
rect 1614 3238 9306 3290
rect 9358 3238 9370 3290
rect 9422 3238 9434 3290
rect 9486 3238 9498 3290
rect 9550 3238 9562 3290
rect 9614 3238 41306 3290
rect 41358 3238 41370 3290
rect 41422 3238 41434 3290
rect 41486 3238 41498 3290
rect 41550 3238 41562 3290
rect 41614 3238 43516 3290
rect 460 3216 43516 3238
rect 31021 3179 31079 3185
rect 31021 3145 31033 3179
rect 31067 3176 31079 3179
rect 31067 3148 33640 3176
rect 31067 3145 31079 3148
rect 31021 3139 31079 3145
rect 32214 3108 32220 3120
rect 30392 3080 32220 3108
rect 28074 3000 28080 3052
rect 28132 3040 28138 3052
rect 29822 3040 29828 3052
rect 28132 3012 29828 3040
rect 28132 3000 28138 3012
rect 29822 3000 29828 3012
rect 29880 3000 29886 3052
rect 30392 3040 30420 3080
rect 32214 3068 32220 3080
rect 32272 3068 32278 3120
rect 33612 3108 33640 3148
rect 33778 3136 33784 3188
rect 33836 3136 33842 3188
rect 36354 3136 36360 3188
rect 36412 3176 36418 3188
rect 36538 3176 36544 3188
rect 36412 3148 36544 3176
rect 36412 3136 36418 3148
rect 36538 3136 36544 3148
rect 36596 3136 36602 3188
rect 36725 3179 36783 3185
rect 36725 3145 36737 3179
rect 36771 3176 36783 3179
rect 39022 3176 39028 3188
rect 36771 3148 39028 3176
rect 36771 3145 36783 3148
rect 36725 3139 36783 3145
rect 39022 3136 39028 3148
rect 39080 3136 39086 3188
rect 33962 3108 33968 3120
rect 32324 3080 33548 3108
rect 33612 3080 33968 3108
rect 30300 3012 30420 3040
rect 30745 3043 30803 3049
rect 27709 2975 27767 2981
rect 27709 2941 27721 2975
rect 27755 2972 27767 2975
rect 28166 2972 28172 2984
rect 27755 2944 28172 2972
rect 27755 2941 27767 2944
rect 27709 2935 27767 2941
rect 28166 2932 28172 2944
rect 28224 2932 28230 2984
rect 28442 2932 28448 2984
rect 28500 2932 28506 2984
rect 28718 2932 28724 2984
rect 28776 2932 28782 2984
rect 30300 2981 30328 3012
rect 30745 3009 30757 3043
rect 30791 3040 30803 3043
rect 32030 3040 32036 3052
rect 30791 3012 32036 3040
rect 30791 3009 30803 3012
rect 30745 3003 30803 3009
rect 32030 3000 32036 3012
rect 32088 3000 32094 3052
rect 30285 2975 30343 2981
rect 30285 2941 30297 2975
rect 30331 2941 30343 2975
rect 30285 2935 30343 2941
rect 30374 2932 30380 2984
rect 30432 2932 30438 2984
rect 30650 2932 30656 2984
rect 30708 2932 30714 2984
rect 30929 2975 30987 2981
rect 30929 2941 30941 2975
rect 30975 2972 30987 2975
rect 31662 2972 31668 2984
rect 30975 2944 31668 2972
rect 30975 2941 30987 2944
rect 30929 2935 30987 2941
rect 31662 2932 31668 2944
rect 31720 2932 31726 2984
rect 31846 2932 31852 2984
rect 31904 2972 31910 2984
rect 32324 2972 32352 3080
rect 32398 3000 32404 3052
rect 32456 3040 32462 3052
rect 32456 3012 32812 3040
rect 32456 3000 32462 3012
rect 31904 2944 32352 2972
rect 32677 2975 32735 2981
rect 31904 2932 31910 2944
rect 32677 2941 32689 2975
rect 32723 2941 32735 2975
rect 32784 2972 32812 3012
rect 33318 3000 33324 3052
rect 33376 3000 33382 3052
rect 33520 3040 33548 3080
rect 33962 3068 33968 3080
rect 34020 3068 34026 3120
rect 36078 3068 36084 3120
rect 36136 3108 36142 3120
rect 37182 3108 37188 3120
rect 36136 3080 37188 3108
rect 36136 3068 36142 3080
rect 37182 3068 37188 3080
rect 37240 3108 37246 3120
rect 37240 3080 37688 3108
rect 37240 3068 37246 3080
rect 34517 3043 34575 3049
rect 34517 3040 34529 3043
rect 33520 3012 34529 3040
rect 34517 3009 34529 3012
rect 34563 3040 34575 3043
rect 34882 3040 34888 3052
rect 34563 3012 34888 3040
rect 34563 3009 34575 3012
rect 34517 3003 34575 3009
rect 34882 3000 34888 3012
rect 34940 3000 34946 3052
rect 36354 3000 36360 3052
rect 36412 3040 36418 3052
rect 36412 3012 37136 3040
rect 36412 3000 36418 3012
rect 32953 2975 33011 2981
rect 32953 2972 32965 2975
rect 32784 2944 32965 2972
rect 32677 2935 32735 2941
rect 32953 2941 32965 2944
rect 32999 2941 33011 2975
rect 32953 2935 33011 2941
rect 24762 2864 24768 2916
rect 24820 2904 24826 2916
rect 26053 2907 26111 2913
rect 26053 2904 26065 2907
rect 24820 2876 26065 2904
rect 24820 2864 24826 2876
rect 26053 2873 26065 2876
rect 26099 2873 26111 2907
rect 26053 2867 26111 2873
rect 26326 2864 26332 2916
rect 26384 2904 26390 2916
rect 26513 2907 26571 2913
rect 26513 2904 26525 2907
rect 26384 2876 26525 2904
rect 26384 2864 26390 2876
rect 26513 2873 26525 2876
rect 26559 2904 26571 2907
rect 27801 2907 27859 2913
rect 27801 2904 27813 2907
rect 26559 2876 27813 2904
rect 26559 2873 26571 2876
rect 26513 2867 26571 2873
rect 27801 2873 27813 2876
rect 27847 2873 27859 2907
rect 27801 2867 27859 2873
rect 28353 2907 28411 2913
rect 28353 2873 28365 2907
rect 28399 2904 28411 2907
rect 29086 2904 29092 2916
rect 28399 2876 29092 2904
rect 28399 2873 28411 2876
rect 28353 2867 28411 2873
rect 29086 2864 29092 2876
rect 29144 2864 29150 2916
rect 30469 2907 30527 2913
rect 30469 2873 30481 2907
rect 30515 2904 30527 2907
rect 31478 2904 31484 2916
rect 30515 2876 31484 2904
rect 30515 2873 30527 2876
rect 30469 2867 30527 2873
rect 31478 2864 31484 2876
rect 31536 2864 31542 2916
rect 31757 2907 31815 2913
rect 31757 2873 31769 2907
rect 31803 2873 31815 2907
rect 32692 2904 32720 2935
rect 33226 2932 33232 2984
rect 33284 2932 33290 2984
rect 33336 2972 33364 3000
rect 33505 2975 33563 2981
rect 33505 2972 33517 2975
rect 33336 2944 33517 2972
rect 33505 2941 33517 2944
rect 33551 2941 33563 2975
rect 33505 2935 33563 2941
rect 34241 2975 34299 2981
rect 34241 2941 34253 2975
rect 34287 2972 34299 2975
rect 34606 2972 34612 2984
rect 34287 2944 34612 2972
rect 34287 2941 34299 2944
rect 34241 2935 34299 2941
rect 34606 2932 34612 2944
rect 34664 2932 34670 2984
rect 34974 2932 34980 2984
rect 35032 2972 35038 2984
rect 35529 2975 35587 2981
rect 35529 2972 35541 2975
rect 35032 2944 35541 2972
rect 35032 2932 35038 2944
rect 35529 2941 35541 2944
rect 35575 2941 35587 2975
rect 35529 2935 35587 2941
rect 35618 2932 35624 2984
rect 35676 2932 35682 2984
rect 35802 2932 35808 2984
rect 35860 2972 35866 2984
rect 36464 2981 36676 2982
rect 36173 2975 36231 2981
rect 36173 2972 36185 2975
rect 35860 2944 36185 2972
rect 35860 2932 35866 2944
rect 36173 2941 36185 2944
rect 36219 2941 36231 2975
rect 36173 2935 36231 2941
rect 36464 2975 36691 2981
rect 36464 2954 36645 2975
rect 33045 2907 33103 2913
rect 33045 2904 33057 2907
rect 32692 2876 33057 2904
rect 31757 2867 31815 2873
rect 33045 2873 33057 2876
rect 33091 2873 33103 2907
rect 33597 2907 33655 2913
rect 33597 2904 33609 2907
rect 33045 2867 33103 2873
rect 33152 2876 33609 2904
rect 25958 2796 25964 2848
rect 26016 2796 26022 2848
rect 27982 2796 27988 2848
rect 28040 2796 28046 2848
rect 28629 2839 28687 2845
rect 28629 2805 28641 2839
rect 28675 2836 28687 2839
rect 30374 2836 30380 2848
rect 28675 2808 30380 2836
rect 28675 2805 28687 2808
rect 28629 2799 28687 2805
rect 30374 2796 30380 2808
rect 30432 2796 30438 2848
rect 30558 2796 30564 2848
rect 30616 2836 30622 2848
rect 31205 2839 31263 2845
rect 31205 2836 31217 2839
rect 30616 2808 31217 2836
rect 30616 2796 30622 2808
rect 31205 2805 31217 2808
rect 31251 2805 31263 2839
rect 31205 2799 31263 2805
rect 31294 2796 31300 2848
rect 31352 2836 31358 2848
rect 31772 2836 31800 2867
rect 31352 2808 31800 2836
rect 31352 2796 31358 2808
rect 32950 2796 32956 2848
rect 33008 2836 33014 2848
rect 33152 2836 33180 2876
rect 33597 2873 33609 2876
rect 33643 2873 33655 2907
rect 33597 2867 33655 2873
rect 35066 2864 35072 2916
rect 35124 2904 35130 2916
rect 35636 2904 35664 2932
rect 35124 2876 35664 2904
rect 36081 2907 36139 2913
rect 35124 2864 35130 2876
rect 36081 2873 36093 2907
rect 36127 2904 36139 2907
rect 36464 2904 36492 2954
rect 36633 2941 36645 2954
rect 36679 2941 36691 2975
rect 36633 2935 36691 2941
rect 36127 2876 36492 2904
rect 37108 2904 37136 3012
rect 37458 3000 37464 3052
rect 37516 3000 37522 3052
rect 37182 2932 37188 2984
rect 37240 2932 37246 2984
rect 37553 2975 37611 2981
rect 37553 2941 37565 2975
rect 37599 2974 37611 2975
rect 37660 2974 37688 3080
rect 38010 3068 38016 3120
rect 38068 3108 38074 3120
rect 38657 3111 38715 3117
rect 38657 3108 38669 3111
rect 38068 3080 38669 3108
rect 38068 3068 38074 3080
rect 38657 3077 38669 3080
rect 38703 3077 38715 3111
rect 38657 3071 38715 3077
rect 38473 3043 38531 3049
rect 38473 3040 38485 3043
rect 37599 2946 37688 2974
rect 37844 3012 38485 3040
rect 37599 2941 37611 2946
rect 37553 2935 37611 2941
rect 37844 2904 37872 3012
rect 38473 3009 38485 3012
rect 38519 3009 38531 3043
rect 38473 3003 38531 3009
rect 38013 2975 38071 2981
rect 38013 2941 38025 2975
rect 38059 2941 38071 2975
rect 38013 2935 38071 2941
rect 37108 2876 37872 2904
rect 38028 2904 38056 2935
rect 38102 2932 38108 2984
rect 38160 2972 38166 2984
rect 38289 2975 38347 2981
rect 38289 2972 38301 2975
rect 38160 2944 38301 2972
rect 38160 2932 38166 2944
rect 38289 2941 38301 2944
rect 38335 2941 38347 2975
rect 38289 2935 38347 2941
rect 38194 2904 38200 2916
rect 38028 2876 38200 2904
rect 36127 2873 36139 2876
rect 36081 2867 36139 2873
rect 38194 2864 38200 2876
rect 38252 2864 38258 2916
rect 33008 2808 33180 2836
rect 33321 2839 33379 2845
rect 33008 2796 33014 2808
rect 33321 2805 33333 2839
rect 33367 2836 33379 2839
rect 34330 2836 34336 2848
rect 33367 2808 34336 2836
rect 33367 2805 33379 2808
rect 33321 2799 33379 2805
rect 34330 2796 34336 2808
rect 34388 2796 34394 2848
rect 36265 2839 36323 2845
rect 36265 2805 36277 2839
rect 36311 2836 36323 2839
rect 37734 2836 37740 2848
rect 36311 2808 37740 2836
rect 36311 2805 36323 2808
rect 36265 2799 36323 2805
rect 37734 2796 37740 2808
rect 37792 2796 37798 2848
rect 38010 2796 38016 2848
rect 38068 2836 38074 2848
rect 38105 2839 38163 2845
rect 38105 2836 38117 2839
rect 38068 2808 38117 2836
rect 38068 2796 38074 2808
rect 38105 2805 38117 2808
rect 38151 2805 38163 2839
rect 38105 2799 38163 2805
rect 38838 2796 38844 2848
rect 38896 2796 38902 2848
rect 460 2746 43516 2768
rect 460 2694 1946 2746
rect 1998 2694 2010 2746
rect 2062 2694 2074 2746
rect 2126 2694 2138 2746
rect 2190 2694 2202 2746
rect 2254 2694 9946 2746
rect 9998 2694 10010 2746
rect 10062 2694 10074 2746
rect 10126 2694 10138 2746
rect 10190 2694 10202 2746
rect 10254 2694 33946 2746
rect 33998 2694 34010 2746
rect 34062 2694 34074 2746
rect 34126 2694 34138 2746
rect 34190 2694 34202 2746
rect 34254 2694 41946 2746
rect 41998 2694 42010 2746
rect 42062 2694 42074 2746
rect 42126 2694 42138 2746
rect 42190 2694 42202 2746
rect 42254 2694 43516 2746
rect 460 2672 43516 2694
rect 27614 2592 27620 2644
rect 27672 2632 27678 2644
rect 27672 2604 29776 2632
rect 27672 2592 27678 2604
rect 24854 2524 24860 2576
rect 24912 2564 24918 2576
rect 26513 2567 26571 2573
rect 26513 2564 26525 2567
rect 24912 2536 26525 2564
rect 24912 2524 24918 2536
rect 26513 2533 26525 2536
rect 26559 2564 26571 2567
rect 27982 2564 27988 2576
rect 26559 2536 27988 2564
rect 26559 2533 26571 2536
rect 26513 2527 26571 2533
rect 27982 2524 27988 2536
rect 28040 2524 28046 2576
rect 29748 2564 29776 2604
rect 29822 2592 29828 2644
rect 29880 2632 29886 2644
rect 31294 2632 31300 2644
rect 29880 2604 31300 2632
rect 29880 2592 29886 2604
rect 31294 2592 31300 2604
rect 31352 2592 31358 2644
rect 31386 2592 31392 2644
rect 31444 2632 31450 2644
rect 34514 2632 34520 2644
rect 31444 2604 34520 2632
rect 31444 2592 31450 2604
rect 34514 2592 34520 2604
rect 34572 2592 34578 2644
rect 38933 2635 38991 2641
rect 38933 2632 38945 2635
rect 35636 2604 38945 2632
rect 30193 2567 30251 2573
rect 30193 2564 30205 2567
rect 29748 2536 30205 2564
rect 30193 2533 30205 2536
rect 30239 2564 30251 2567
rect 30466 2564 30472 2576
rect 30239 2536 30472 2564
rect 30239 2533 30251 2536
rect 30193 2527 30251 2533
rect 30466 2524 30472 2536
rect 30524 2524 30530 2576
rect 31570 2564 31576 2576
rect 30760 2536 31576 2564
rect 25130 2456 25136 2508
rect 25188 2496 25194 2508
rect 25593 2499 25651 2505
rect 25593 2496 25605 2499
rect 25188 2468 25605 2496
rect 25188 2456 25194 2468
rect 25593 2465 25605 2468
rect 25639 2465 25651 2499
rect 25593 2459 25651 2465
rect 27706 2456 27712 2508
rect 27764 2456 27770 2508
rect 28994 2456 29000 2508
rect 29052 2456 29058 2508
rect 29086 2456 29092 2508
rect 29144 2496 29150 2508
rect 29273 2499 29331 2505
rect 29273 2496 29285 2499
rect 29144 2468 29285 2496
rect 29144 2456 29150 2468
rect 29273 2465 29285 2468
rect 29319 2465 29331 2499
rect 30558 2496 30564 2508
rect 29273 2459 29331 2465
rect 30392 2468 30564 2496
rect 24302 2388 24308 2440
rect 24360 2428 24366 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24360 2400 24593 2428
rect 24360 2388 24366 2400
rect 24581 2397 24593 2400
rect 24627 2428 24639 2431
rect 25869 2431 25927 2437
rect 25869 2428 25881 2431
rect 24627 2400 25881 2428
rect 24627 2397 24639 2400
rect 24581 2391 24639 2397
rect 25869 2397 25881 2400
rect 25915 2397 25927 2431
rect 25869 2391 25927 2397
rect 26878 2388 26884 2440
rect 26936 2428 26942 2440
rect 27985 2431 28043 2437
rect 27985 2428 27997 2431
rect 26936 2400 27997 2428
rect 26936 2388 26942 2400
rect 27985 2397 27997 2400
rect 28031 2428 28043 2431
rect 30392 2428 30420 2468
rect 30558 2456 30564 2468
rect 30616 2456 30622 2508
rect 30760 2505 30788 2536
rect 31570 2524 31576 2536
rect 31628 2524 31634 2576
rect 32950 2524 32956 2576
rect 33008 2564 33014 2576
rect 35636 2573 35664 2604
rect 38933 2601 38945 2604
rect 38979 2601 38991 2635
rect 38933 2595 38991 2601
rect 39114 2592 39120 2644
rect 39172 2632 39178 2644
rect 39853 2635 39911 2641
rect 39853 2632 39865 2635
rect 39172 2604 39865 2632
rect 39172 2592 39178 2604
rect 39853 2601 39865 2604
rect 39899 2601 39911 2635
rect 39853 2595 39911 2601
rect 35621 2567 35679 2573
rect 35621 2564 35633 2567
rect 33008 2536 33088 2564
rect 33008 2524 33014 2536
rect 30745 2499 30803 2505
rect 30745 2465 30757 2499
rect 30791 2465 30803 2499
rect 30745 2459 30803 2465
rect 31018 2456 31024 2508
rect 31076 2456 31082 2508
rect 31478 2456 31484 2508
rect 31536 2456 31542 2508
rect 33060 2505 33088 2536
rect 34532 2536 35633 2564
rect 33045 2499 33103 2505
rect 31588 2468 32996 2496
rect 28031 2400 30420 2428
rect 28031 2397 28043 2400
rect 27985 2391 28043 2397
rect 30466 2388 30472 2440
rect 30524 2428 30530 2440
rect 31588 2428 31616 2468
rect 30524 2400 31616 2428
rect 30524 2388 30530 2400
rect 31662 2388 31668 2440
rect 31720 2428 31726 2440
rect 31941 2431 31999 2437
rect 31941 2428 31953 2431
rect 31720 2400 31953 2428
rect 31720 2388 31726 2400
rect 31941 2397 31953 2400
rect 31987 2428 31999 2431
rect 32122 2428 32128 2440
rect 31987 2400 32128 2428
rect 31987 2397 31999 2400
rect 31941 2391 31999 2397
rect 32122 2388 32128 2400
rect 32180 2388 32186 2440
rect 32968 2428 32996 2468
rect 33045 2465 33057 2499
rect 33091 2465 33103 2499
rect 33045 2459 33103 2465
rect 33413 2431 33471 2437
rect 33413 2428 33425 2431
rect 32968 2400 33425 2428
rect 33413 2397 33425 2400
rect 33459 2428 33471 2431
rect 33594 2428 33600 2440
rect 33459 2400 33600 2428
rect 33459 2397 33471 2400
rect 33413 2391 33471 2397
rect 33594 2388 33600 2400
rect 33652 2388 33658 2440
rect 31478 2320 31484 2372
rect 31536 2360 31542 2372
rect 34532 2360 34560 2536
rect 35621 2533 35633 2536
rect 35667 2533 35679 2567
rect 35621 2527 35679 2533
rect 36538 2524 36544 2576
rect 36596 2564 36602 2576
rect 38838 2564 38844 2576
rect 36596 2536 38332 2564
rect 36596 2524 36602 2536
rect 34609 2499 34667 2505
rect 34609 2465 34621 2499
rect 34655 2496 34667 2499
rect 34698 2496 34704 2508
rect 34655 2468 34704 2496
rect 34655 2465 34667 2468
rect 34609 2459 34667 2465
rect 34698 2456 34704 2468
rect 34756 2456 34762 2508
rect 35894 2456 35900 2508
rect 35952 2456 35958 2508
rect 35989 2499 36047 2505
rect 35989 2465 36001 2499
rect 36035 2465 36047 2499
rect 35989 2459 36047 2465
rect 36449 2499 36507 2505
rect 36449 2465 36461 2499
rect 36495 2496 36507 2499
rect 36633 2499 36691 2505
rect 36633 2496 36645 2499
rect 36495 2468 36645 2496
rect 36495 2465 36507 2468
rect 36449 2459 36507 2465
rect 36633 2465 36645 2468
rect 36679 2465 36691 2499
rect 36633 2459 36691 2465
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 36004 2428 36032 2459
rect 37274 2456 37280 2508
rect 37332 2456 37338 2508
rect 37458 2456 37464 2508
rect 37516 2456 37522 2508
rect 37550 2456 37556 2508
rect 37608 2496 37614 2508
rect 37608 2468 37872 2496
rect 37608 2456 37614 2468
rect 37844 2437 37872 2468
rect 38102 2456 38108 2508
rect 38160 2456 38166 2508
rect 38304 2505 38332 2536
rect 38396 2536 38844 2564
rect 38396 2505 38424 2536
rect 38838 2524 38844 2536
rect 38896 2524 38902 2576
rect 38289 2499 38347 2505
rect 38289 2465 38301 2499
rect 38335 2465 38347 2499
rect 38289 2459 38347 2465
rect 38381 2499 38439 2505
rect 38381 2465 38393 2499
rect 38427 2465 38439 2499
rect 38381 2459 38439 2465
rect 38470 2456 38476 2508
rect 38528 2496 38534 2508
rect 40678 2496 40684 2508
rect 38528 2468 40684 2496
rect 38528 2456 38534 2468
rect 40678 2456 40684 2468
rect 40736 2456 40742 2508
rect 34848 2400 36032 2428
rect 34848 2388 34854 2400
rect 31536 2332 34560 2360
rect 31536 2320 31542 2332
rect 34606 2320 34612 2372
rect 34664 2360 34670 2372
rect 36004 2360 36032 2400
rect 37001 2431 37059 2437
rect 37001 2397 37013 2431
rect 37047 2397 37059 2431
rect 37001 2391 37059 2397
rect 37829 2431 37887 2437
rect 37829 2397 37841 2431
rect 37875 2397 37887 2431
rect 37829 2391 37887 2397
rect 36814 2360 36820 2372
rect 34664 2332 35296 2360
rect 36004 2332 36820 2360
rect 34664 2320 34670 2332
rect 26050 2252 26056 2304
rect 26108 2252 26114 2304
rect 30837 2295 30895 2301
rect 30837 2261 30849 2295
rect 30883 2292 30895 2295
rect 31018 2292 31024 2304
rect 30883 2264 31024 2292
rect 30883 2261 30895 2264
rect 30837 2255 30895 2261
rect 31018 2252 31024 2264
rect 31076 2252 31082 2304
rect 31113 2295 31171 2301
rect 31113 2261 31125 2295
rect 31159 2292 31171 2295
rect 31846 2292 31852 2304
rect 31159 2264 31852 2292
rect 31159 2261 31171 2264
rect 31113 2255 31171 2261
rect 31846 2252 31852 2264
rect 31904 2252 31910 2304
rect 32122 2252 32128 2304
rect 32180 2292 32186 2304
rect 35158 2292 35164 2304
rect 32180 2264 35164 2292
rect 32180 2252 32186 2264
rect 35158 2252 35164 2264
rect 35216 2252 35222 2304
rect 35268 2292 35296 2332
rect 36814 2320 36820 2332
rect 36872 2320 36878 2372
rect 37016 2360 37044 2391
rect 38562 2388 38568 2440
rect 38620 2428 38626 2440
rect 38841 2431 38899 2437
rect 38620 2400 38792 2428
rect 38620 2388 38626 2400
rect 38654 2360 38660 2372
rect 37016 2332 38660 2360
rect 38654 2320 38660 2332
rect 38712 2320 38718 2372
rect 38764 2360 38792 2400
rect 38841 2397 38853 2431
rect 38887 2428 38899 2431
rect 39114 2428 39120 2440
rect 38887 2400 39120 2428
rect 38887 2397 38899 2400
rect 38841 2391 38899 2397
rect 39114 2388 39120 2400
rect 39172 2388 39178 2440
rect 39485 2363 39543 2369
rect 39485 2360 39497 2363
rect 38764 2332 39497 2360
rect 39485 2329 39497 2332
rect 39531 2329 39543 2363
rect 39485 2323 39543 2329
rect 39574 2320 39580 2372
rect 39632 2360 39638 2372
rect 40221 2363 40279 2369
rect 40221 2360 40233 2363
rect 39632 2332 40233 2360
rect 39632 2320 39638 2332
rect 40221 2329 40233 2332
rect 40267 2329 40279 2363
rect 40221 2323 40279 2329
rect 39117 2295 39175 2301
rect 39117 2292 39129 2295
rect 35268 2264 39129 2292
rect 39117 2261 39129 2264
rect 39163 2261 39175 2295
rect 39117 2255 39175 2261
rect 39206 2252 39212 2304
rect 39264 2292 39270 2304
rect 39301 2295 39359 2301
rect 39301 2292 39313 2295
rect 39264 2264 39313 2292
rect 39264 2252 39270 2264
rect 39301 2261 39313 2264
rect 39347 2261 39359 2295
rect 39301 2255 39359 2261
rect 39666 2252 39672 2304
rect 39724 2252 39730 2304
rect 39758 2252 39764 2304
rect 39816 2292 39822 2304
rect 40037 2295 40095 2301
rect 40037 2292 40049 2295
rect 39816 2264 40049 2292
rect 39816 2252 39822 2264
rect 40037 2261 40049 2264
rect 40083 2261 40095 2295
rect 40037 2255 40095 2261
rect 40494 2252 40500 2304
rect 40552 2252 40558 2304
rect 460 2202 43516 2224
rect 460 2150 1306 2202
rect 1358 2150 1370 2202
rect 1422 2150 1434 2202
rect 1486 2150 1498 2202
rect 1550 2150 1562 2202
rect 1614 2150 9306 2202
rect 9358 2150 9370 2202
rect 9422 2150 9434 2202
rect 9486 2150 9498 2202
rect 9550 2150 9562 2202
rect 9614 2150 17306 2202
rect 17358 2150 17370 2202
rect 17422 2150 17434 2202
rect 17486 2150 17498 2202
rect 17550 2150 17562 2202
rect 17614 2150 25306 2202
rect 25358 2150 25370 2202
rect 25422 2150 25434 2202
rect 25486 2150 25498 2202
rect 25550 2150 25562 2202
rect 25614 2150 33306 2202
rect 33358 2150 33370 2202
rect 33422 2150 33434 2202
rect 33486 2150 33498 2202
rect 33550 2150 33562 2202
rect 33614 2150 41306 2202
rect 41358 2150 41370 2202
rect 41422 2150 41434 2202
rect 41486 2150 41498 2202
rect 41550 2150 41562 2202
rect 41614 2150 43516 2202
rect 460 2128 43516 2150
rect 28166 2048 28172 2100
rect 28224 2088 28230 2100
rect 28353 2091 28411 2097
rect 28353 2088 28365 2091
rect 28224 2060 28365 2088
rect 28224 2048 28230 2060
rect 28353 2057 28365 2060
rect 28399 2057 28411 2091
rect 28353 2051 28411 2057
rect 28442 2048 28448 2100
rect 28500 2088 28506 2100
rect 32766 2088 32772 2100
rect 28500 2060 32772 2088
rect 28500 2048 28506 2060
rect 32766 2048 32772 2060
rect 32824 2048 32830 2100
rect 34514 2088 34520 2100
rect 32876 2060 34520 2088
rect 25958 1980 25964 2032
rect 26016 2020 26022 2032
rect 26418 2020 26424 2032
rect 26016 1992 26424 2020
rect 26016 1980 26022 1992
rect 26418 1980 26424 1992
rect 26476 1980 26482 2032
rect 29086 1980 29092 2032
rect 29144 2020 29150 2032
rect 31662 2020 31668 2032
rect 29144 1992 31668 2020
rect 29144 1980 29150 1992
rect 31662 1980 31668 1992
rect 31720 1980 31726 2032
rect 24578 1912 24584 1964
rect 24636 1952 24642 1964
rect 25777 1955 25835 1961
rect 25777 1952 25789 1955
rect 24636 1924 25789 1952
rect 24636 1912 24642 1924
rect 25777 1921 25789 1924
rect 25823 1952 25835 1955
rect 26050 1952 26056 1964
rect 25823 1924 26056 1952
rect 25823 1921 25835 1924
rect 25777 1915 25835 1921
rect 26050 1912 26056 1924
rect 26108 1912 26114 1964
rect 28718 1912 28724 1964
rect 28776 1952 28782 1964
rect 28776 1924 30512 1952
rect 28776 1912 28782 1924
rect 25038 1844 25044 1896
rect 25096 1844 25102 1896
rect 25501 1887 25559 1893
rect 25501 1853 25513 1887
rect 25547 1884 25559 1887
rect 25590 1884 25596 1896
rect 25547 1856 25596 1884
rect 25547 1853 25559 1856
rect 25501 1847 25559 1853
rect 25590 1844 25596 1856
rect 25648 1844 25654 1896
rect 26786 1844 26792 1896
rect 26844 1844 26850 1896
rect 28258 1844 28264 1896
rect 28316 1844 28322 1896
rect 28534 1844 28540 1896
rect 28592 1844 28598 1896
rect 28626 1844 28632 1896
rect 28684 1884 28690 1896
rect 28684 1856 30236 1884
rect 28684 1844 28690 1856
rect 23750 1776 23756 1828
rect 23808 1816 23814 1828
rect 24029 1819 24087 1825
rect 24029 1816 24041 1819
rect 23808 1788 24041 1816
rect 23808 1776 23814 1788
rect 24029 1785 24041 1788
rect 24075 1785 24087 1819
rect 24029 1779 24087 1785
rect 27890 1776 27896 1828
rect 27948 1776 27954 1828
rect 29089 1819 29147 1825
rect 29089 1816 29101 1819
rect 28552 1788 29101 1816
rect 27062 1708 27068 1760
rect 27120 1748 27126 1760
rect 28552 1748 28580 1788
rect 29089 1785 29101 1788
rect 29135 1816 29147 1819
rect 29914 1816 29920 1828
rect 29135 1788 29920 1816
rect 29135 1785 29147 1788
rect 29089 1779 29147 1785
rect 29914 1776 29920 1788
rect 29972 1776 29978 1828
rect 30208 1816 30236 1856
rect 30282 1844 30288 1896
rect 30340 1844 30346 1896
rect 30374 1844 30380 1896
rect 30432 1844 30438 1896
rect 30484 1884 30512 1924
rect 30834 1912 30840 1964
rect 30892 1952 30898 1964
rect 31938 1952 31944 1964
rect 30892 1924 31944 1952
rect 30892 1912 30898 1924
rect 31938 1912 31944 1924
rect 31996 1952 32002 1964
rect 32876 1952 32904 2060
rect 34514 2048 34520 2060
rect 34572 2048 34578 2100
rect 36722 2048 36728 2100
rect 36780 2088 36786 2100
rect 36780 2060 38654 2088
rect 36780 2048 36786 2060
rect 35158 1980 35164 2032
rect 35216 2020 35222 2032
rect 38470 2020 38476 2032
rect 35216 1992 35756 2020
rect 35216 1980 35222 1992
rect 31996 1924 32904 1952
rect 31996 1912 32002 1924
rect 33042 1912 33048 1964
rect 33100 1912 33106 1964
rect 33318 1912 33324 1964
rect 33376 1912 33382 1964
rect 34422 1952 34428 1964
rect 33428 1924 34428 1952
rect 30484 1856 31754 1884
rect 31386 1816 31392 1828
rect 30208 1788 31392 1816
rect 31386 1776 31392 1788
rect 31444 1776 31450 1828
rect 31726 1816 31754 1856
rect 31846 1844 31852 1896
rect 31904 1844 31910 1896
rect 33060 1816 33088 1912
rect 33428 1893 33456 1924
rect 34422 1912 34428 1924
rect 34480 1912 34486 1964
rect 34606 1912 34612 1964
rect 34664 1912 34670 1964
rect 35728 1952 35756 1992
rect 37292 1992 38476 2020
rect 35989 1955 36047 1961
rect 35989 1952 36001 1955
rect 35636 1924 36001 1952
rect 33413 1887 33471 1893
rect 33413 1853 33425 1887
rect 33459 1853 33471 1887
rect 33413 1847 33471 1853
rect 33873 1887 33931 1893
rect 33873 1853 33885 1887
rect 33919 1884 33931 1887
rect 33962 1884 33968 1896
rect 33919 1856 33968 1884
rect 33919 1853 33931 1856
rect 33873 1847 33931 1853
rect 33962 1844 33968 1856
rect 34020 1844 34026 1896
rect 34057 1887 34115 1893
rect 34057 1853 34069 1887
rect 34103 1853 34115 1887
rect 34057 1847 34115 1853
rect 31726 1788 33088 1816
rect 33778 1776 33784 1828
rect 33836 1816 33842 1828
rect 34072 1816 34100 1847
rect 35526 1844 35532 1896
rect 35584 1844 35590 1896
rect 33836 1788 34100 1816
rect 35636 1816 35664 1924
rect 35989 1921 36001 1924
rect 36035 1921 36047 1955
rect 35989 1915 36047 1921
rect 36630 1912 36636 1964
rect 36688 1952 36694 1964
rect 37292 1952 37320 1992
rect 38470 1980 38476 1992
rect 38528 1980 38534 2032
rect 38626 2020 38654 2060
rect 39574 2048 39580 2100
rect 39632 2048 39638 2100
rect 39853 2091 39911 2097
rect 39853 2057 39865 2091
rect 39899 2088 39911 2091
rect 40218 2088 40224 2100
rect 39899 2060 40224 2088
rect 39899 2057 39911 2060
rect 39853 2051 39911 2057
rect 40218 2048 40224 2060
rect 40276 2088 40282 2100
rect 40865 2091 40923 2097
rect 40865 2088 40877 2091
rect 40276 2060 40877 2088
rect 40276 2048 40282 2060
rect 40865 2057 40877 2060
rect 40911 2057 40923 2091
rect 40865 2051 40923 2057
rect 38746 2020 38752 2032
rect 38626 1992 38752 2020
rect 38746 1980 38752 1992
rect 38804 1980 38810 2032
rect 39301 2023 39359 2029
rect 39301 1989 39313 2023
rect 39347 2020 39359 2023
rect 39482 2020 39488 2032
rect 39347 1992 39488 2020
rect 39347 1989 39359 1992
rect 39301 1983 39359 1989
rect 39482 1980 39488 1992
rect 39540 2020 39546 2032
rect 39758 2020 39764 2032
rect 39540 1992 39764 2020
rect 39540 1980 39546 1992
rect 39758 1980 39764 1992
rect 39816 1980 39822 2032
rect 40129 2023 40187 2029
rect 40129 1989 40141 2023
rect 40175 2020 40187 2023
rect 40175 1992 40908 2020
rect 40175 1989 40187 1992
rect 40129 1983 40187 1989
rect 37369 1955 37427 1961
rect 37369 1952 37381 1955
rect 36688 1924 37136 1952
rect 37292 1924 37381 1952
rect 36688 1912 36694 1924
rect 35710 1844 35716 1896
rect 35768 1884 35774 1896
rect 37001 1887 37059 1893
rect 37001 1884 37013 1887
rect 35768 1856 37013 1884
rect 35768 1844 35774 1856
rect 37001 1853 37013 1856
rect 37047 1853 37059 1887
rect 37108 1884 37136 1924
rect 37369 1921 37381 1924
rect 37415 1921 37427 1955
rect 37369 1915 37427 1921
rect 38197 1955 38255 1961
rect 38197 1921 38209 1955
rect 38243 1952 38255 1955
rect 38243 1924 39712 1952
rect 38243 1921 38255 1924
rect 38197 1915 38255 1921
rect 37737 1887 37795 1893
rect 37737 1884 37749 1887
rect 37108 1856 37749 1884
rect 37001 1847 37059 1853
rect 37737 1853 37749 1856
rect 37783 1853 37795 1887
rect 37737 1847 37795 1853
rect 37550 1816 37556 1828
rect 35636 1788 37556 1816
rect 33836 1776 33842 1788
rect 37550 1776 37556 1788
rect 37608 1776 37614 1828
rect 27120 1720 28580 1748
rect 28629 1751 28687 1757
rect 27120 1708 27126 1720
rect 28629 1717 28641 1751
rect 28675 1748 28687 1751
rect 29270 1748 29276 1760
rect 28675 1720 29276 1748
rect 28675 1717 28687 1720
rect 28629 1711 28687 1717
rect 29270 1708 29276 1720
rect 29328 1708 29334 1760
rect 37752 1748 37780 1847
rect 37826 1844 37832 1896
rect 37884 1844 37890 1896
rect 38378 1844 38384 1896
rect 38436 1884 38442 1896
rect 38565 1887 38623 1893
rect 38565 1884 38577 1887
rect 38436 1856 38577 1884
rect 38436 1844 38442 1856
rect 38565 1853 38577 1856
rect 38611 1853 38623 1887
rect 38565 1847 38623 1853
rect 38580 1816 38608 1847
rect 38654 1844 38660 1896
rect 38712 1844 38718 1896
rect 39209 1887 39267 1893
rect 39209 1853 39221 1887
rect 39255 1884 39267 1887
rect 39298 1884 39304 1896
rect 39255 1856 39304 1884
rect 39255 1853 39267 1856
rect 39209 1847 39267 1853
rect 39298 1844 39304 1856
rect 39356 1844 39362 1896
rect 39390 1844 39396 1896
rect 39448 1884 39454 1896
rect 39485 1887 39543 1893
rect 39485 1884 39497 1887
rect 39448 1856 39497 1884
rect 39448 1844 39454 1856
rect 39485 1853 39497 1856
rect 39531 1853 39543 1887
rect 39485 1847 39543 1853
rect 39684 1878 39712 1924
rect 40880 1896 40908 1992
rect 39761 1887 39819 1893
rect 39761 1878 39773 1887
rect 39684 1853 39773 1878
rect 39807 1853 39819 1887
rect 39684 1850 39819 1853
rect 39761 1847 39819 1850
rect 40037 1887 40095 1893
rect 40037 1853 40049 1887
rect 40083 1884 40095 1887
rect 40126 1884 40132 1896
rect 40083 1856 40132 1884
rect 40083 1853 40095 1856
rect 40037 1847 40095 1853
rect 40126 1844 40132 1856
rect 40184 1844 40190 1896
rect 40862 1844 40868 1896
rect 40920 1884 40926 1896
rect 41049 1887 41107 1893
rect 41049 1884 41061 1887
rect 40920 1856 41061 1884
rect 40920 1844 40926 1856
rect 41049 1853 41061 1856
rect 41095 1853 41107 1887
rect 41049 1847 41107 1853
rect 38580 1788 39528 1816
rect 38562 1748 38568 1760
rect 37752 1720 38568 1748
rect 38562 1708 38568 1720
rect 38620 1708 38626 1760
rect 38746 1708 38752 1760
rect 38804 1708 38810 1760
rect 38933 1751 38991 1757
rect 38933 1717 38945 1751
rect 38979 1748 38991 1751
rect 39206 1748 39212 1760
rect 38979 1720 39212 1748
rect 38979 1717 38991 1720
rect 38933 1711 38991 1717
rect 39206 1708 39212 1720
rect 39264 1708 39270 1760
rect 39500 1748 39528 1788
rect 39850 1776 39856 1828
rect 39908 1816 39914 1828
rect 40497 1819 40555 1825
rect 40497 1816 40509 1819
rect 39908 1788 40509 1816
rect 39908 1776 39914 1788
rect 40497 1785 40509 1788
rect 40543 1785 40555 1819
rect 40497 1779 40555 1785
rect 40313 1751 40371 1757
rect 40313 1748 40325 1751
rect 39500 1720 40325 1748
rect 40313 1717 40325 1720
rect 40359 1717 40371 1751
rect 40313 1711 40371 1717
rect 40402 1708 40408 1760
rect 40460 1748 40466 1760
rect 40681 1751 40739 1757
rect 40681 1748 40693 1751
rect 40460 1720 40693 1748
rect 40460 1708 40466 1720
rect 40681 1717 40693 1720
rect 40727 1717 40739 1751
rect 40681 1711 40739 1717
rect 40770 1708 40776 1760
rect 40828 1748 40834 1760
rect 41233 1751 41291 1757
rect 41233 1748 41245 1751
rect 40828 1720 41245 1748
rect 40828 1708 40834 1720
rect 41233 1717 41245 1720
rect 41279 1717 41291 1751
rect 41233 1711 41291 1717
rect 460 1658 43516 1680
rect 460 1606 1946 1658
rect 1998 1606 2010 1658
rect 2062 1606 2074 1658
rect 2126 1606 2138 1658
rect 2190 1606 2202 1658
rect 2254 1606 9946 1658
rect 9998 1606 10010 1658
rect 10062 1606 10074 1658
rect 10126 1606 10138 1658
rect 10190 1606 10202 1658
rect 10254 1606 17946 1658
rect 17998 1606 18010 1658
rect 18062 1606 18074 1658
rect 18126 1606 18138 1658
rect 18190 1606 18202 1658
rect 18254 1606 25946 1658
rect 25998 1606 26010 1658
rect 26062 1606 26074 1658
rect 26126 1606 26138 1658
rect 26190 1606 26202 1658
rect 26254 1606 33946 1658
rect 33998 1606 34010 1658
rect 34062 1606 34074 1658
rect 34126 1606 34138 1658
rect 34190 1606 34202 1658
rect 34254 1606 41946 1658
rect 41998 1606 42010 1658
rect 42062 1606 42074 1658
rect 42126 1606 42138 1658
rect 42190 1606 42202 1658
rect 42254 1606 43516 1658
rect 460 1584 43516 1606
rect 25130 1504 25136 1556
rect 25188 1504 25194 1556
rect 25961 1547 26019 1553
rect 25961 1513 25973 1547
rect 26007 1544 26019 1547
rect 26786 1544 26792 1556
rect 26007 1516 26792 1544
rect 26007 1513 26019 1516
rect 25961 1507 26019 1513
rect 26786 1504 26792 1516
rect 26844 1504 26850 1556
rect 30098 1504 30104 1556
rect 30156 1544 30162 1556
rect 30156 1516 34008 1544
rect 30156 1504 30162 1516
rect 25593 1479 25651 1485
rect 25593 1445 25605 1479
rect 25639 1476 25651 1479
rect 25639 1448 26372 1476
rect 25639 1445 25651 1448
rect 25593 1439 25651 1445
rect 23566 1368 23572 1420
rect 23624 1368 23630 1420
rect 25222 1368 25228 1420
rect 25280 1368 25286 1420
rect 25682 1368 25688 1420
rect 25740 1368 25746 1420
rect 25774 1368 25780 1420
rect 25832 1408 25838 1420
rect 26344 1417 26372 1448
rect 26418 1436 26424 1488
rect 26476 1476 26482 1488
rect 28721 1479 28779 1485
rect 28721 1476 28733 1479
rect 26476 1448 28733 1476
rect 26476 1436 26482 1448
rect 28721 1445 28733 1448
rect 28767 1445 28779 1479
rect 28721 1439 28779 1445
rect 29362 1436 29368 1488
rect 29420 1476 29426 1488
rect 33980 1476 34008 1516
rect 34054 1504 34060 1556
rect 34112 1544 34118 1556
rect 39206 1544 39212 1556
rect 34112 1516 39212 1544
rect 34112 1504 34118 1516
rect 39206 1504 39212 1516
rect 39264 1504 39270 1556
rect 40034 1544 40040 1556
rect 39868 1516 40040 1544
rect 35345 1479 35403 1485
rect 35345 1476 35357 1479
rect 29420 1448 33456 1476
rect 33980 1448 35357 1476
rect 29420 1436 29426 1448
rect 26053 1411 26111 1417
rect 26053 1408 26065 1411
rect 25832 1380 26065 1408
rect 25832 1368 25838 1380
rect 26053 1377 26065 1380
rect 26099 1377 26111 1411
rect 26053 1371 26111 1377
rect 26329 1411 26387 1417
rect 26329 1377 26341 1411
rect 26375 1377 26387 1411
rect 26329 1371 26387 1377
rect 21542 1300 21548 1352
rect 21600 1340 21606 1352
rect 22554 1340 22560 1352
rect 21600 1312 22560 1340
rect 21600 1300 21606 1312
rect 22554 1300 22560 1312
rect 22612 1300 22618 1352
rect 23474 1300 23480 1352
rect 23532 1340 23538 1352
rect 24029 1343 24087 1349
rect 24029 1340 24041 1343
rect 23532 1312 24041 1340
rect 23532 1300 23538 1312
rect 24029 1309 24041 1312
rect 24075 1309 24087 1343
rect 24029 1303 24087 1309
rect 25958 1300 25964 1352
rect 26016 1340 26022 1352
rect 26436 1340 26464 1436
rect 27430 1368 27436 1420
rect 27488 1408 27494 1420
rect 27540 1408 27660 1414
rect 27488 1386 27660 1408
rect 27488 1380 27568 1386
rect 27488 1368 27494 1380
rect 26016 1312 26464 1340
rect 27632 1340 27660 1386
rect 27982 1368 27988 1420
rect 28040 1368 28046 1420
rect 29270 1368 29276 1420
rect 29328 1368 29334 1420
rect 29656 1380 29868 1408
rect 29656 1340 29684 1380
rect 27632 1312 29684 1340
rect 29733 1343 29791 1349
rect 26016 1300 26022 1312
rect 29733 1309 29745 1343
rect 29779 1309 29791 1343
rect 29733 1303 29791 1309
rect 23385 1275 23443 1281
rect 23385 1241 23397 1275
rect 23431 1272 23443 1275
rect 25774 1272 25780 1284
rect 23431 1244 25780 1272
rect 23431 1241 23443 1244
rect 23385 1235 23443 1241
rect 25774 1232 25780 1244
rect 25832 1232 25838 1284
rect 26510 1232 26516 1284
rect 26568 1272 26574 1284
rect 29748 1272 29776 1303
rect 26568 1244 29776 1272
rect 29840 1272 29868 1380
rect 30834 1368 30840 1420
rect 30892 1368 30898 1420
rect 31018 1368 31024 1420
rect 31076 1408 31082 1420
rect 31481 1411 31539 1417
rect 31481 1408 31493 1411
rect 31076 1380 31493 1408
rect 31076 1368 31082 1380
rect 31481 1377 31493 1380
rect 31527 1377 31539 1411
rect 31481 1371 31539 1377
rect 32030 1368 32036 1420
rect 32088 1408 32094 1420
rect 32953 1411 33011 1417
rect 32953 1408 32965 1411
rect 32088 1380 32965 1408
rect 32088 1368 32094 1380
rect 32953 1377 32965 1380
rect 32999 1377 33011 1411
rect 32953 1371 33011 1377
rect 30742 1300 30748 1352
rect 30800 1300 30806 1352
rect 31297 1343 31355 1349
rect 31297 1309 31309 1343
rect 31343 1309 31355 1343
rect 31297 1303 31355 1309
rect 32677 1343 32735 1349
rect 32677 1309 32689 1343
rect 32723 1340 32735 1343
rect 32766 1340 32772 1352
rect 32723 1312 32772 1340
rect 32723 1309 32735 1312
rect 32677 1303 32735 1309
rect 31202 1272 31208 1284
rect 29840 1244 31208 1272
rect 26568 1232 26574 1244
rect 23750 1164 23756 1216
rect 23808 1204 23814 1216
rect 25317 1207 25375 1213
rect 25317 1204 25329 1207
rect 23808 1176 25329 1204
rect 23808 1164 23814 1176
rect 25317 1173 25329 1176
rect 25363 1173 25375 1207
rect 29748 1204 29776 1244
rect 31202 1232 31208 1244
rect 31260 1232 31266 1284
rect 31312 1272 31340 1303
rect 32766 1300 32772 1312
rect 32824 1300 32830 1352
rect 33428 1349 33456 1448
rect 35345 1445 35357 1448
rect 35391 1476 35403 1479
rect 36354 1476 36360 1488
rect 35391 1448 36360 1476
rect 35391 1445 35403 1448
rect 35345 1439 35403 1445
rect 36354 1436 36360 1448
rect 36412 1436 36418 1488
rect 36722 1476 36728 1488
rect 36556 1448 36728 1476
rect 34238 1368 34244 1420
rect 34296 1408 34302 1420
rect 34425 1411 34483 1417
rect 34425 1408 34437 1411
rect 34296 1380 34437 1408
rect 34296 1368 34302 1380
rect 34425 1377 34437 1380
rect 34471 1377 34483 1411
rect 35989 1411 36047 1417
rect 35989 1408 36001 1411
rect 34425 1371 34483 1377
rect 35820 1380 36001 1408
rect 33413 1343 33471 1349
rect 33413 1309 33425 1343
rect 33459 1340 33471 1343
rect 34054 1340 34060 1352
rect 33459 1312 34060 1340
rect 33459 1309 33471 1312
rect 33413 1303 33471 1309
rect 34054 1300 34060 1312
rect 34112 1300 34118 1352
rect 34330 1300 34336 1352
rect 34388 1340 34394 1352
rect 35820 1340 35848 1380
rect 35989 1377 36001 1380
rect 36035 1408 36047 1411
rect 36556 1408 36584 1448
rect 36722 1436 36728 1448
rect 36780 1436 36786 1488
rect 36906 1436 36912 1488
rect 36964 1476 36970 1488
rect 39758 1476 39764 1488
rect 36964 1448 38056 1476
rect 36964 1436 36970 1448
rect 36035 1380 36584 1408
rect 36035 1377 36047 1380
rect 35989 1371 36047 1377
rect 36630 1368 36636 1420
rect 36688 1368 36694 1420
rect 36814 1368 36820 1420
rect 36872 1408 36878 1420
rect 37185 1411 37243 1417
rect 37185 1408 37197 1411
rect 36872 1380 37197 1408
rect 36872 1368 36878 1380
rect 37185 1377 37197 1380
rect 37231 1377 37243 1411
rect 37185 1371 37243 1377
rect 37461 1411 37519 1417
rect 37461 1377 37473 1411
rect 37507 1377 37519 1411
rect 37461 1371 37519 1377
rect 34388 1312 35848 1340
rect 35897 1343 35955 1349
rect 34388 1300 34394 1312
rect 35897 1309 35909 1343
rect 35943 1340 35955 1343
rect 36262 1340 36268 1352
rect 35943 1312 36268 1340
rect 35943 1309 35955 1312
rect 35897 1303 35955 1309
rect 36262 1300 36268 1312
rect 36320 1300 36326 1352
rect 36449 1343 36507 1349
rect 36449 1309 36461 1343
rect 36495 1340 36507 1343
rect 37476 1340 37504 1371
rect 37550 1368 37556 1420
rect 37608 1408 37614 1420
rect 37918 1408 37924 1420
rect 37608 1380 37924 1408
rect 37608 1368 37614 1380
rect 37918 1368 37924 1380
rect 37976 1368 37982 1420
rect 38028 1417 38056 1448
rect 39040 1448 39764 1476
rect 38013 1411 38071 1417
rect 38013 1377 38025 1411
rect 38059 1377 38071 1411
rect 38013 1371 38071 1377
rect 38194 1368 38200 1420
rect 38252 1408 38258 1420
rect 39040 1417 39068 1448
rect 39758 1436 39764 1448
rect 39816 1436 39822 1488
rect 38289 1411 38347 1417
rect 38289 1408 38301 1411
rect 38252 1380 38301 1408
rect 38252 1368 38258 1380
rect 38289 1377 38301 1380
rect 38335 1377 38347 1411
rect 38289 1371 38347 1377
rect 39025 1411 39083 1417
rect 39025 1377 39037 1411
rect 39071 1377 39083 1411
rect 39025 1371 39083 1377
rect 39114 1368 39120 1420
rect 39172 1368 39178 1420
rect 39868 1417 39896 1516
rect 40034 1504 40040 1516
rect 40092 1544 40098 1556
rect 41233 1547 41291 1553
rect 41233 1544 41245 1547
rect 40092 1516 41245 1544
rect 40092 1504 40098 1516
rect 41233 1513 41245 1516
rect 41279 1513 41291 1547
rect 41233 1507 41291 1513
rect 40865 1479 40923 1485
rect 40865 1445 40877 1479
rect 40911 1476 40923 1479
rect 41138 1476 41144 1488
rect 40911 1448 41144 1476
rect 40911 1445 40923 1448
rect 40865 1439 40923 1445
rect 41138 1436 41144 1448
rect 41196 1476 41202 1488
rect 41196 1448 41414 1476
rect 41196 1436 41202 1448
rect 39853 1411 39911 1417
rect 39853 1377 39865 1411
rect 39899 1377 39911 1411
rect 39853 1371 39911 1377
rect 40034 1368 40040 1420
rect 40092 1368 40098 1420
rect 40494 1368 40500 1420
rect 40552 1368 40558 1420
rect 40773 1411 40831 1417
rect 40773 1377 40785 1411
rect 40819 1377 40831 1411
rect 40773 1371 40831 1377
rect 36495 1312 37504 1340
rect 37829 1343 37887 1349
rect 36495 1309 36507 1312
rect 36449 1303 36507 1309
rect 37829 1309 37841 1343
rect 37875 1309 37887 1343
rect 37829 1303 37887 1309
rect 35710 1272 35716 1284
rect 31312 1244 35716 1272
rect 35710 1232 35716 1244
rect 35768 1232 35774 1284
rect 37844 1272 37872 1303
rect 38654 1300 38660 1352
rect 38712 1300 38718 1352
rect 39485 1343 39543 1349
rect 39485 1309 39497 1343
rect 39531 1340 39543 1343
rect 40126 1340 40132 1352
rect 39531 1312 40132 1340
rect 39531 1309 39543 1312
rect 39485 1303 39543 1309
rect 40126 1300 40132 1312
rect 40184 1300 40190 1352
rect 40313 1343 40371 1349
rect 40313 1309 40325 1343
rect 40359 1340 40371 1343
rect 40788 1340 40816 1371
rect 40359 1312 40816 1340
rect 41386 1340 41414 1448
rect 41785 1343 41843 1349
rect 41785 1340 41797 1343
rect 41386 1312 41797 1340
rect 40359 1309 40371 1312
rect 40313 1303 40371 1309
rect 41785 1309 41797 1312
rect 41831 1309 41843 1343
rect 41785 1303 41843 1309
rect 40402 1272 40408 1284
rect 37844 1244 40408 1272
rect 40402 1232 40408 1244
rect 40460 1232 40466 1284
rect 40954 1232 40960 1284
rect 41012 1272 41018 1284
rect 41012 1244 41184 1272
rect 41012 1232 41018 1244
rect 36354 1204 36360 1216
rect 29748 1176 36360 1204
rect 25317 1167 25375 1173
rect 36354 1164 36360 1176
rect 36412 1164 36418 1216
rect 36722 1164 36728 1216
rect 36780 1164 36786 1216
rect 36814 1164 36820 1216
rect 36872 1204 36878 1216
rect 39298 1204 39304 1216
rect 36872 1176 39304 1204
rect 36872 1164 36878 1176
rect 39298 1164 39304 1176
rect 39356 1164 39362 1216
rect 39942 1164 39948 1216
rect 40000 1204 40006 1216
rect 41049 1207 41107 1213
rect 41049 1204 41061 1207
rect 40000 1176 41061 1204
rect 40000 1164 40006 1176
rect 41049 1173 41061 1176
rect 41095 1173 41107 1207
rect 41156 1204 41184 1244
rect 41322 1232 41328 1284
rect 41380 1272 41386 1284
rect 42153 1275 42211 1281
rect 42153 1272 42165 1275
rect 41380 1244 42165 1272
rect 41380 1232 41386 1244
rect 42153 1241 42165 1244
rect 42199 1241 42211 1275
rect 42153 1235 42211 1241
rect 41417 1207 41475 1213
rect 41417 1204 41429 1207
rect 41156 1176 41429 1204
rect 41049 1167 41107 1173
rect 41417 1173 41429 1176
rect 41463 1173 41475 1207
rect 41417 1167 41475 1173
rect 41966 1164 41972 1216
rect 42024 1164 42030 1216
rect 460 1114 43516 1136
rect 460 1062 1306 1114
rect 1358 1062 1370 1114
rect 1422 1062 1434 1114
rect 1486 1062 1498 1114
rect 1550 1062 1562 1114
rect 1614 1062 9306 1114
rect 9358 1062 9370 1114
rect 9422 1062 9434 1114
rect 9486 1062 9498 1114
rect 9550 1062 9562 1114
rect 9614 1062 17306 1114
rect 17358 1062 17370 1114
rect 17422 1062 17434 1114
rect 17486 1062 17498 1114
rect 17550 1062 17562 1114
rect 17614 1062 25306 1114
rect 25358 1062 25370 1114
rect 25422 1062 25434 1114
rect 25486 1062 25498 1114
rect 25550 1062 25562 1114
rect 25614 1062 33306 1114
rect 33358 1062 33370 1114
rect 33422 1062 33434 1114
rect 33486 1062 33498 1114
rect 33550 1062 33562 1114
rect 33614 1062 41306 1114
rect 41358 1062 41370 1114
rect 41422 1062 41434 1114
rect 41486 1062 41498 1114
rect 41550 1062 41562 1114
rect 41614 1062 43516 1114
rect 460 1040 43516 1062
rect 23201 1003 23259 1009
rect 23201 969 23213 1003
rect 23247 1000 23259 1003
rect 23566 1000 23572 1012
rect 23247 972 23572 1000
rect 23247 969 23259 972
rect 23201 963 23259 969
rect 23566 960 23572 972
rect 23624 960 23630 1012
rect 25038 960 25044 1012
rect 25096 1000 25102 1012
rect 25317 1003 25375 1009
rect 25317 1000 25329 1003
rect 25096 972 25329 1000
rect 25096 960 25102 972
rect 25317 969 25329 972
rect 25363 969 25375 1003
rect 25317 963 25375 969
rect 25682 960 25688 1012
rect 25740 1000 25746 1012
rect 25869 1003 25927 1009
rect 25869 1000 25881 1003
rect 25740 972 25881 1000
rect 25740 960 25746 972
rect 25869 969 25881 972
rect 25915 969 25927 1003
rect 25869 963 25927 969
rect 27706 960 27712 1012
rect 27764 1000 27770 1012
rect 27893 1003 27951 1009
rect 27893 1000 27905 1003
rect 27764 972 27905 1000
rect 27764 960 27770 972
rect 27893 969 27905 972
rect 27939 969 27951 1003
rect 27893 963 27951 969
rect 27982 960 27988 1012
rect 28040 1000 28046 1012
rect 28169 1003 28227 1009
rect 28169 1000 28181 1003
rect 28040 972 28181 1000
rect 28040 960 28046 972
rect 28169 969 28181 972
rect 28215 969 28227 1003
rect 28169 963 28227 969
rect 30282 960 30288 1012
rect 30340 1000 30346 1012
rect 30745 1003 30803 1009
rect 30745 1000 30757 1003
rect 30340 972 30757 1000
rect 30340 960 30346 972
rect 30745 969 30757 972
rect 30791 969 30803 1003
rect 30745 963 30803 969
rect 31202 960 31208 1012
rect 31260 960 31266 1012
rect 32214 960 32220 1012
rect 32272 1000 32278 1012
rect 33045 1003 33103 1009
rect 33045 1000 33057 1003
rect 32272 972 33057 1000
rect 32272 960 32278 972
rect 33045 969 33057 972
rect 33091 969 33103 1003
rect 33045 963 33103 969
rect 36354 960 36360 1012
rect 36412 960 36418 1012
rect 38654 960 38660 1012
rect 38712 1000 38718 1012
rect 38712 972 40908 1000
rect 38712 960 38718 972
rect 23474 892 23480 944
rect 23532 932 23538 944
rect 26053 935 26111 941
rect 26053 932 26065 935
rect 23532 904 26065 932
rect 23532 892 23538 904
rect 26053 901 26065 904
rect 26099 901 26111 935
rect 26053 895 26111 901
rect 28994 892 29000 944
rect 29052 932 29058 944
rect 30469 935 30527 941
rect 30469 932 30481 935
rect 29052 904 30481 932
rect 29052 892 29058 904
rect 30469 901 30481 904
rect 30515 901 30527 935
rect 30469 895 30527 901
rect 30834 892 30840 944
rect 30892 932 30898 944
rect 34606 932 34612 944
rect 30892 904 34612 932
rect 30892 892 30898 904
rect 34606 892 34612 904
rect 34664 892 34670 944
rect 36722 892 36728 944
rect 36780 932 36786 944
rect 40221 935 40279 941
rect 36780 904 40172 932
rect 36780 892 36786 904
rect 23017 867 23075 873
rect 23017 833 23029 867
rect 23063 864 23075 867
rect 23198 864 23204 876
rect 23063 836 23204 864
rect 23063 833 23075 836
rect 23017 827 23075 833
rect 23198 824 23204 836
rect 23256 864 23262 876
rect 24213 867 24271 873
rect 24213 864 24225 867
rect 23256 836 24225 864
rect 23256 824 23262 836
rect 24213 833 24225 836
rect 24259 833 24271 867
rect 24213 827 24271 833
rect 24946 824 24952 876
rect 25004 864 25010 876
rect 26789 867 26847 873
rect 26789 864 26801 867
rect 25004 836 25544 864
rect 25004 824 25010 836
rect 23290 756 23296 808
rect 23348 756 23354 808
rect 23569 799 23627 805
rect 23569 765 23581 799
rect 23615 796 23627 799
rect 23658 796 23664 808
rect 23615 768 23664 796
rect 23615 765 23627 768
rect 23569 759 23627 765
rect 23658 756 23664 768
rect 23716 756 23722 808
rect 23753 799 23811 805
rect 23753 765 23765 799
rect 23799 765 23811 799
rect 23753 759 23811 765
rect 23477 731 23535 737
rect 23477 697 23489 731
rect 23523 728 23535 731
rect 23768 728 23796 759
rect 25222 756 25228 808
rect 25280 756 25286 808
rect 25516 805 25544 836
rect 25608 836 26801 864
rect 25501 799 25559 805
rect 25501 765 25513 799
rect 25547 765 25559 799
rect 25501 759 25559 765
rect 23523 700 23796 728
rect 23523 697 23535 700
rect 23477 691 23535 697
rect 24026 688 24032 740
rect 24084 728 24090 740
rect 24762 728 24768 740
rect 24084 700 24768 728
rect 24084 688 24090 700
rect 24762 688 24768 700
rect 24820 728 24826 740
rect 25608 728 25636 836
rect 26789 833 26801 836
rect 26835 833 26847 867
rect 26789 827 26847 833
rect 27338 824 27344 876
rect 27396 864 27402 876
rect 33321 867 33379 873
rect 27396 836 31754 864
rect 27396 824 27402 836
rect 25777 799 25835 805
rect 25777 765 25789 799
rect 25823 796 25835 799
rect 25866 796 25872 808
rect 25823 768 25872 796
rect 25823 765 25835 768
rect 25777 759 25835 765
rect 25866 756 25872 768
rect 25924 756 25930 808
rect 26329 799 26387 805
rect 26329 765 26341 799
rect 26375 765 26387 799
rect 26329 759 26387 765
rect 26344 728 26372 759
rect 27798 756 27804 808
rect 27856 756 27862 808
rect 28074 756 28080 808
rect 28132 756 28138 808
rect 28350 756 28356 808
rect 28408 756 28414 808
rect 28445 799 28503 805
rect 28445 765 28457 799
rect 28491 796 28503 799
rect 28905 799 28963 805
rect 28905 796 28917 799
rect 28491 768 28917 796
rect 28491 765 28503 768
rect 28445 759 28503 765
rect 28905 765 28917 768
rect 28951 765 28963 799
rect 28905 759 28963 765
rect 30374 756 30380 808
rect 30432 756 30438 808
rect 30650 756 30656 808
rect 30708 756 30714 808
rect 30926 756 30932 808
rect 30984 756 30990 808
rect 31021 799 31079 805
rect 31021 765 31033 799
rect 31067 796 31079 799
rect 31481 799 31539 805
rect 31481 796 31493 799
rect 31067 768 31493 796
rect 31067 765 31079 768
rect 31021 759 31079 765
rect 31481 765 31493 768
rect 31527 765 31539 799
rect 31481 759 31539 765
rect 24820 700 25636 728
rect 25792 700 26372 728
rect 24820 688 24826 700
rect 25593 663 25651 669
rect 25593 629 25605 663
rect 25639 660 25651 663
rect 25792 660 25820 700
rect 27890 688 27896 740
rect 27948 728 27954 740
rect 28629 731 28687 737
rect 28629 728 28641 731
rect 27948 700 28641 728
rect 27948 688 27954 700
rect 28629 697 28641 700
rect 28675 697 28687 731
rect 29825 731 29883 737
rect 29825 728 29837 731
rect 28629 691 28687 697
rect 28966 700 29837 728
rect 25639 632 25820 660
rect 25639 629 25651 632
rect 25593 623 25651 629
rect 25866 620 25872 672
rect 25924 660 25930 672
rect 28966 660 28994 700
rect 29825 697 29837 700
rect 29871 697 29883 731
rect 31726 728 31754 836
rect 33321 833 33333 867
rect 33367 864 33379 867
rect 33778 864 33784 876
rect 33367 836 33784 864
rect 33367 833 33379 836
rect 33321 827 33379 833
rect 33778 824 33784 836
rect 33836 824 33842 876
rect 33873 867 33931 873
rect 33873 833 33885 867
rect 33919 864 33931 867
rect 35897 867 35955 873
rect 33919 836 35572 864
rect 33919 833 33931 836
rect 33873 827 33931 833
rect 32950 756 32956 808
rect 33008 756 33014 808
rect 33413 799 33471 805
rect 33413 765 33425 799
rect 33459 796 33471 799
rect 33686 796 33692 808
rect 33459 768 33692 796
rect 33459 765 33471 768
rect 33413 759 33471 765
rect 33686 756 33692 768
rect 33744 756 33750 808
rect 33962 756 33968 808
rect 34020 796 34026 808
rect 35544 805 35572 836
rect 35897 833 35909 867
rect 35943 864 35955 867
rect 39761 867 39819 873
rect 35943 836 39436 864
rect 35943 833 35955 836
rect 35897 827 35955 833
rect 34057 799 34115 805
rect 34057 796 34069 799
rect 34020 768 34069 796
rect 34020 756 34026 768
rect 34057 765 34069 768
rect 34103 765 34115 799
rect 35529 799 35587 805
rect 34057 759 34115 765
rect 34348 768 35388 796
rect 32677 731 32735 737
rect 32677 728 32689 731
rect 29825 691 29883 697
rect 29932 700 31340 728
rect 31726 700 32689 728
rect 25924 632 28994 660
rect 25924 620 25930 632
rect 29546 620 29552 672
rect 29604 660 29610 672
rect 29932 660 29960 700
rect 29604 632 29960 660
rect 31312 660 31340 700
rect 32677 697 32689 700
rect 32723 728 32735 731
rect 34348 728 34376 768
rect 32723 700 34376 728
rect 32723 697 32735 700
rect 32677 691 32735 697
rect 35250 688 35256 740
rect 35308 688 35314 740
rect 35268 660 35296 688
rect 31312 632 35296 660
rect 35360 660 35388 768
rect 35529 765 35541 799
rect 35575 765 35587 799
rect 35529 759 35587 765
rect 35986 756 35992 808
rect 36044 796 36050 808
rect 36262 796 36268 808
rect 36044 768 36268 796
rect 36044 756 36050 768
rect 36262 756 36268 768
rect 36320 756 36326 808
rect 36446 756 36452 808
rect 36504 796 36510 808
rect 36633 799 36691 805
rect 36633 796 36645 799
rect 36504 768 36645 796
rect 36504 756 36510 768
rect 36633 765 36645 768
rect 36679 765 36691 799
rect 36633 759 36691 765
rect 37642 756 37648 808
rect 37700 796 37706 808
rect 38105 799 38163 805
rect 38105 796 38117 799
rect 37700 768 38117 796
rect 37700 756 37706 768
rect 38105 765 38117 768
rect 38151 765 38163 799
rect 38105 759 38163 765
rect 38473 799 38531 805
rect 38473 765 38485 799
rect 38519 765 38531 799
rect 38473 759 38531 765
rect 37458 688 37464 740
rect 37516 728 37522 740
rect 37553 731 37611 737
rect 37553 728 37565 731
rect 37516 700 37565 728
rect 37516 688 37522 700
rect 37553 697 37565 700
rect 37599 697 37611 731
rect 38488 728 38516 759
rect 38562 756 38568 808
rect 38620 796 38626 808
rect 38657 799 38715 805
rect 38657 796 38669 799
rect 38620 768 38669 796
rect 38620 756 38626 768
rect 38657 765 38669 768
rect 38703 765 38715 799
rect 38657 759 38715 765
rect 38930 756 38936 808
rect 38988 796 38994 808
rect 39209 799 39267 805
rect 39209 796 39221 799
rect 38988 768 39221 796
rect 38988 756 38994 768
rect 39209 765 39221 768
rect 39255 765 39267 799
rect 39209 759 39267 765
rect 39298 756 39304 808
rect 39356 756 39362 808
rect 39408 796 39436 836
rect 39761 833 39773 867
rect 39807 864 39819 867
rect 40034 864 40040 876
rect 39807 836 40040 864
rect 39807 833 39819 836
rect 39761 827 39819 833
rect 40034 824 40040 836
rect 40092 824 40098 876
rect 40144 805 40172 904
rect 40221 901 40233 935
rect 40267 932 40279 935
rect 40310 932 40316 944
rect 40267 904 40316 932
rect 40267 901 40279 904
rect 40221 895 40279 901
rect 40310 892 40316 904
rect 40368 932 40374 944
rect 40770 932 40776 944
rect 40368 904 40776 932
rect 40368 892 40374 904
rect 40770 892 40776 904
rect 40828 892 40834 944
rect 40880 864 40908 972
rect 41230 960 41236 1012
rect 41288 1000 41294 1012
rect 41325 1003 41383 1009
rect 41325 1000 41337 1003
rect 41288 972 41337 1000
rect 41288 960 41294 972
rect 41325 969 41337 972
rect 41371 969 41383 1003
rect 41325 963 41383 969
rect 41782 960 41788 1012
rect 41840 960 41846 1012
rect 40788 836 40908 864
rect 39853 799 39911 805
rect 39853 796 39865 799
rect 39408 768 39865 796
rect 39853 765 39865 768
rect 39899 765 39911 799
rect 39853 759 39911 765
rect 40129 799 40187 805
rect 40129 765 40141 799
rect 40175 765 40187 799
rect 40129 759 40187 765
rect 40402 756 40408 808
rect 40460 756 40466 808
rect 40494 756 40500 808
rect 40552 756 40558 808
rect 40678 756 40684 808
rect 40736 756 40742 808
rect 40788 790 40816 836
rect 41046 824 41052 876
rect 41104 864 41110 876
rect 41966 864 41972 876
rect 41104 836 41972 864
rect 41104 824 41110 836
rect 41966 824 41972 836
rect 42024 824 42030 876
rect 40949 801 41007 807
rect 40949 798 40961 801
rect 40880 790 40961 798
rect 40788 770 40961 790
rect 40788 762 40908 770
rect 40949 767 40961 770
rect 40995 767 41007 801
rect 40949 761 41007 767
rect 41233 799 41291 805
rect 41233 765 41245 799
rect 41279 765 41291 799
rect 41233 759 41291 765
rect 41248 728 41276 759
rect 41322 756 41328 808
rect 41380 796 41386 808
rect 42153 799 42211 805
rect 42153 796 42165 799
rect 41380 768 42165 796
rect 41380 756 41386 768
rect 42153 765 42165 768
rect 42199 765 42211 799
rect 42153 759 42211 765
rect 42334 756 42340 808
rect 42392 756 42398 808
rect 42521 731 42579 737
rect 42521 728 42533 731
rect 38488 700 41276 728
rect 41386 700 42533 728
rect 37553 691 37611 697
rect 38933 663 38991 669
rect 38933 660 38945 663
rect 35360 632 38945 660
rect 29604 620 29610 632
rect 38933 629 38945 632
rect 38979 629 38991 663
rect 38933 623 38991 629
rect 39022 620 39028 672
rect 39080 660 39086 672
rect 39945 663 40003 669
rect 39945 660 39957 663
rect 39080 632 39957 660
rect 39080 620 39086 632
rect 39945 629 39957 632
rect 39991 660 40003 663
rect 40402 660 40408 672
rect 39991 632 40408 660
rect 39991 629 40003 632
rect 39945 623 40003 629
rect 40402 620 40408 632
rect 40460 620 40466 672
rect 40770 620 40776 672
rect 40828 660 40834 672
rect 41386 660 41414 700
rect 42521 697 42533 700
rect 42567 697 42579 731
rect 42521 691 42579 697
rect 40828 632 41414 660
rect 40828 620 40834 632
rect 41506 620 41512 672
rect 41564 620 41570 672
rect 41782 620 41788 672
rect 41840 660 41846 672
rect 41969 663 42027 669
rect 41969 660 41981 663
rect 41840 632 41981 660
rect 41840 620 41846 632
rect 41969 629 41981 632
rect 42015 629 42027 663
rect 41969 623 42027 629
rect 460 570 43516 592
rect 460 518 1946 570
rect 1998 518 2010 570
rect 2062 518 2074 570
rect 2126 518 2138 570
rect 2190 518 2202 570
rect 2254 518 9946 570
rect 9998 518 10010 570
rect 10062 518 10074 570
rect 10126 518 10138 570
rect 10190 518 10202 570
rect 10254 518 17946 570
rect 17998 518 18010 570
rect 18062 518 18074 570
rect 18126 518 18138 570
rect 18190 518 18202 570
rect 18254 518 25946 570
rect 25998 518 26010 570
rect 26062 518 26074 570
rect 26126 518 26138 570
rect 26190 518 26202 570
rect 26254 518 33946 570
rect 33998 518 34010 570
rect 34062 518 34074 570
rect 34126 518 34138 570
rect 34190 518 34202 570
rect 34254 518 41946 570
rect 41998 518 42010 570
rect 42062 518 42074 570
rect 42126 518 42138 570
rect 42190 518 42202 570
rect 42254 518 43516 570
rect 460 496 43516 518
rect 25222 416 25228 468
rect 25280 456 25286 468
rect 27798 456 27804 468
rect 25280 428 27804 456
rect 25280 416 25286 428
rect 27798 416 27804 428
rect 27856 416 27862 468
rect 27982 416 27988 468
rect 28040 456 28046 468
rect 28626 456 28632 468
rect 28040 428 28632 456
rect 28040 416 28046 428
rect 28626 416 28632 428
rect 28684 416 28690 468
rect 33870 416 33876 468
rect 33928 456 33934 468
rect 34422 456 34428 468
rect 33928 428 34428 456
rect 33928 416 33934 428
rect 34422 416 34428 428
rect 34480 416 34486 468
rect 38194 416 38200 468
rect 38252 456 38258 468
rect 38838 456 38844 468
rect 38252 428 38844 456
rect 38252 416 38258 428
rect 38838 416 38844 428
rect 38896 416 38902 468
rect 39942 456 39948 468
rect 38948 428 39948 456
rect 24946 348 24952 400
rect 25004 388 25010 400
rect 27430 388 27436 400
rect 25004 360 27436 388
rect 25004 348 25010 360
rect 27430 348 27436 360
rect 27488 348 27494 400
rect 31294 348 31300 400
rect 31352 388 31358 400
rect 37458 388 37464 400
rect 31352 360 37464 388
rect 31352 348 31358 360
rect 37458 348 37464 360
rect 37516 388 37522 400
rect 38948 388 38976 428
rect 39942 416 39948 428
rect 40000 416 40006 468
rect 40402 416 40408 468
rect 40460 456 40466 468
rect 41046 456 41052 468
rect 40460 428 41052 456
rect 40460 416 40466 428
rect 41046 416 41052 428
rect 41104 416 41110 468
rect 37516 360 38976 388
rect 37516 348 37522 360
rect 39022 348 39028 400
rect 39080 388 39086 400
rect 40770 388 40776 400
rect 39080 360 40776 388
rect 39080 348 39086 360
rect 40770 348 40776 360
rect 40828 348 40834 400
rect 35250 280 35256 332
rect 35308 320 35314 332
rect 41506 320 41512 332
rect 35308 292 41512 320
rect 35308 280 35314 292
rect 41506 280 41512 292
rect 41564 280 41570 332
rect 40678 212 40684 264
rect 40736 252 40742 264
rect 41230 252 41236 264
rect 40736 224 41236 252
rect 40736 212 40742 224
rect 41230 212 41236 224
rect 41288 212 41294 264
rect 41782 252 41788 264
rect 41386 224 41788 252
rect 38286 144 38292 196
rect 38344 184 38350 196
rect 40954 184 40960 196
rect 38344 156 40960 184
rect 38344 144 38350 156
rect 40954 144 40960 156
rect 41012 144 41018 196
rect 39298 76 39304 128
rect 39356 116 39362 128
rect 41386 116 41414 224
rect 41782 212 41788 224
rect 41840 212 41846 264
rect 39356 88 41414 116
rect 39356 76 39362 88
rect 38562 8 38568 60
rect 38620 48 38626 60
rect 40218 48 40224 60
rect 38620 20 40224 48
rect 38620 8 38626 20
rect 40218 8 40224 20
rect 40276 8 40282 60
<< via1 >>
rect 31760 11568 31812 11620
rect 32680 11568 32732 11620
rect 10048 11500 10100 11552
rect 10416 11500 10468 11552
rect 18052 11500 18104 11552
rect 18696 11500 18748 11552
rect 25872 11500 25924 11552
rect 26056 11500 26108 11552
rect 30104 11500 30156 11552
rect 30748 11500 30800 11552
rect 31392 11500 31444 11552
rect 32128 11500 32180 11552
rect 32220 11500 32272 11552
rect 33508 11500 33560 11552
rect 1946 11398 1998 11450
rect 2010 11398 2062 11450
rect 2074 11398 2126 11450
rect 2138 11398 2190 11450
rect 2202 11398 2254 11450
rect 9946 11398 9998 11450
rect 10010 11398 10062 11450
rect 10074 11398 10126 11450
rect 10138 11398 10190 11450
rect 10202 11398 10254 11450
rect 17946 11398 17998 11450
rect 18010 11398 18062 11450
rect 18074 11398 18126 11450
rect 18138 11398 18190 11450
rect 18202 11398 18254 11450
rect 25946 11398 25998 11450
rect 26010 11398 26062 11450
rect 26074 11398 26126 11450
rect 26138 11398 26190 11450
rect 26202 11398 26254 11450
rect 33946 11398 33998 11450
rect 34010 11398 34062 11450
rect 34074 11398 34126 11450
rect 34138 11398 34190 11450
rect 34202 11398 34254 11450
rect 41946 11398 41998 11450
rect 42010 11398 42062 11450
rect 42074 11398 42126 11450
rect 42138 11398 42190 11450
rect 42202 11398 42254 11450
rect 25504 11296 25556 11348
rect 26884 11296 26936 11348
rect 24308 11203 24360 11212
rect 24308 11169 24317 11203
rect 24317 11169 24351 11203
rect 24351 11169 24360 11203
rect 24308 11160 24360 11169
rect 25964 11160 26016 11212
rect 26240 11160 26292 11212
rect 27436 11296 27488 11348
rect 28632 11296 28684 11348
rect 29368 11296 29420 11348
rect 27528 11160 27580 11212
rect 29920 11296 29972 11348
rect 30104 11339 30156 11348
rect 30104 11305 30113 11339
rect 30113 11305 30147 11339
rect 30147 11305 30156 11339
rect 30104 11296 30156 11305
rect 27160 11092 27212 11144
rect 28632 11160 28684 11212
rect 30932 11296 30984 11348
rect 31116 11296 31168 11348
rect 31852 11296 31904 11348
rect 31760 11271 31812 11280
rect 29092 11092 29144 11144
rect 30656 11203 30708 11212
rect 30656 11169 30665 11203
rect 30665 11169 30699 11203
rect 30699 11169 30708 11203
rect 30656 11160 30708 11169
rect 30840 11203 30892 11212
rect 30840 11169 30849 11203
rect 30849 11169 30883 11203
rect 30883 11169 30892 11203
rect 30840 11160 30892 11169
rect 31760 11237 31769 11271
rect 31769 11237 31803 11271
rect 31803 11237 31812 11271
rect 31760 11228 31812 11237
rect 29184 11024 29236 11076
rect 9128 10956 9180 11008
rect 9496 10956 9548 11008
rect 17132 10956 17184 11008
rect 17500 10956 17552 11008
rect 24216 10999 24268 11008
rect 24216 10965 24225 10999
rect 24225 10965 24259 10999
rect 24259 10965 24268 10999
rect 24216 10956 24268 10965
rect 25228 10956 25280 11008
rect 26424 10999 26476 11008
rect 26424 10965 26433 10999
rect 26433 10965 26467 10999
rect 26467 10965 26476 10999
rect 26424 10956 26476 10965
rect 27896 10999 27948 11008
rect 27896 10965 27905 10999
rect 27905 10965 27939 10999
rect 27939 10965 27948 10999
rect 27896 10956 27948 10965
rect 28172 10999 28224 11008
rect 28172 10965 28181 10999
rect 28181 10965 28215 10999
rect 28215 10965 28224 10999
rect 28172 10956 28224 10965
rect 28632 10999 28684 11008
rect 28632 10965 28641 10999
rect 28641 10965 28675 10999
rect 28675 10965 28684 10999
rect 28632 10956 28684 10965
rect 28724 10956 28776 11008
rect 32036 11160 32088 11212
rect 32588 11296 32640 11348
rect 32772 11296 32824 11348
rect 33784 11296 33836 11348
rect 33876 11339 33928 11348
rect 33876 11305 33885 11339
rect 33885 11305 33919 11339
rect 33919 11305 33928 11339
rect 33876 11296 33928 11305
rect 32220 11092 32272 11144
rect 32588 11203 32640 11212
rect 32588 11169 32597 11203
rect 32597 11169 32631 11203
rect 32631 11169 32640 11203
rect 32588 11160 32640 11169
rect 32772 11203 32824 11212
rect 32772 11169 32781 11203
rect 32781 11169 32815 11203
rect 32815 11169 32824 11203
rect 32772 11160 32824 11169
rect 32864 11203 32916 11212
rect 32864 11169 32873 11203
rect 32873 11169 32907 11203
rect 32907 11169 32916 11203
rect 32864 11160 32916 11169
rect 34336 11296 34388 11348
rect 33508 11135 33560 11144
rect 33508 11101 33517 11135
rect 33517 11101 33551 11135
rect 33551 11101 33560 11135
rect 33508 11092 33560 11101
rect 29552 10999 29604 11008
rect 29552 10965 29561 10999
rect 29561 10965 29595 10999
rect 29595 10965 29604 10999
rect 29552 10956 29604 10965
rect 29828 10999 29880 11008
rect 29828 10965 29837 10999
rect 29837 10965 29871 10999
rect 29871 10965 29880 10999
rect 29828 10956 29880 10965
rect 30472 10999 30524 11008
rect 30472 10965 30481 10999
rect 30481 10965 30515 10999
rect 30515 10965 30524 10999
rect 30472 10956 30524 10965
rect 31484 11024 31536 11076
rect 31852 10956 31904 11008
rect 31944 10956 31996 11008
rect 32772 10956 32824 11008
rect 33692 11024 33744 11076
rect 33140 10956 33192 11008
rect 33784 10956 33836 11008
rect 1306 10854 1358 10906
rect 1370 10854 1422 10906
rect 1434 10854 1486 10906
rect 1498 10854 1550 10906
rect 1562 10854 1614 10906
rect 9306 10854 9358 10906
rect 9370 10854 9422 10906
rect 9434 10854 9486 10906
rect 9498 10854 9550 10906
rect 9562 10854 9614 10906
rect 17306 10854 17358 10906
rect 17370 10854 17422 10906
rect 17434 10854 17486 10906
rect 17498 10854 17550 10906
rect 17562 10854 17614 10906
rect 25306 10854 25358 10906
rect 25370 10854 25422 10906
rect 25434 10854 25486 10906
rect 25498 10854 25550 10906
rect 25562 10854 25614 10906
rect 33306 10854 33358 10906
rect 33370 10854 33422 10906
rect 33434 10854 33486 10906
rect 33498 10854 33550 10906
rect 33562 10854 33614 10906
rect 41306 10854 41358 10906
rect 41370 10854 41422 10906
rect 41434 10854 41486 10906
rect 41498 10854 41550 10906
rect 41562 10854 41614 10906
rect 24308 10591 24360 10600
rect 24308 10557 24317 10591
rect 24317 10557 24351 10591
rect 24351 10557 24360 10591
rect 24308 10548 24360 10557
rect 25780 10752 25832 10804
rect 26332 10684 26384 10736
rect 26608 10616 26660 10668
rect 27160 10548 27212 10600
rect 27528 10591 27580 10600
rect 27528 10557 27537 10591
rect 27537 10557 27571 10591
rect 27571 10557 27580 10591
rect 27528 10548 27580 10557
rect 28816 10752 28868 10804
rect 30472 10752 30524 10804
rect 32220 10752 32272 10804
rect 29552 10684 29604 10736
rect 31208 10684 31260 10736
rect 30656 10548 30708 10600
rect 31668 10548 31720 10600
rect 32036 10616 32088 10668
rect 33232 10752 33284 10804
rect 33048 10480 33100 10532
rect 24492 10455 24544 10464
rect 24492 10421 24501 10455
rect 24501 10421 24535 10455
rect 24535 10421 24544 10455
rect 24492 10412 24544 10421
rect 24860 10455 24912 10464
rect 24860 10421 24869 10455
rect 24869 10421 24903 10455
rect 24903 10421 24912 10455
rect 24860 10412 24912 10421
rect 25136 10455 25188 10464
rect 25136 10421 25145 10455
rect 25145 10421 25179 10455
rect 25179 10421 25188 10455
rect 25136 10412 25188 10421
rect 27712 10455 27764 10464
rect 27712 10421 27721 10455
rect 27721 10421 27755 10455
rect 27755 10421 27764 10455
rect 27712 10412 27764 10421
rect 30012 10412 30064 10464
rect 33232 10412 33284 10464
rect 1946 10310 1998 10362
rect 2010 10310 2062 10362
rect 2074 10310 2126 10362
rect 2138 10310 2190 10362
rect 2202 10310 2254 10362
rect 9946 10310 9998 10362
rect 10010 10310 10062 10362
rect 10074 10310 10126 10362
rect 10138 10310 10190 10362
rect 10202 10310 10254 10362
rect 17946 10310 17998 10362
rect 18010 10310 18062 10362
rect 18074 10310 18126 10362
rect 18138 10310 18190 10362
rect 18202 10310 18254 10362
rect 25946 10310 25998 10362
rect 26010 10310 26062 10362
rect 26074 10310 26126 10362
rect 26138 10310 26190 10362
rect 26202 10310 26254 10362
rect 33946 10310 33998 10362
rect 34010 10310 34062 10362
rect 34074 10310 34126 10362
rect 34138 10310 34190 10362
rect 34202 10310 34254 10362
rect 41946 10310 41998 10362
rect 42010 10310 42062 10362
rect 42074 10310 42126 10362
rect 42138 10310 42190 10362
rect 42202 10310 42254 10362
rect 14740 10251 14792 10260
rect 14740 10217 14749 10251
rect 14749 10217 14783 10251
rect 14783 10217 14792 10251
rect 14740 10208 14792 10217
rect 16672 10251 16724 10260
rect 16672 10217 16681 10251
rect 16681 10217 16715 10251
rect 16715 10217 16724 10251
rect 16672 10208 16724 10217
rect 17224 10208 17276 10260
rect 18052 10208 18104 10260
rect 18696 10208 18748 10260
rect 19984 10208 20036 10260
rect 20996 10208 21048 10260
rect 21364 10208 21416 10260
rect 14464 10140 14516 10192
rect 15016 10140 15068 10192
rect 17776 10140 17828 10192
rect 18604 10140 18656 10192
rect 19800 10140 19852 10192
rect 20444 10140 20496 10192
rect 13452 10072 13504 10124
rect 18788 10072 18840 10124
rect 20352 10072 20404 10124
rect 20812 10072 20864 10124
rect 24308 10072 24360 10124
rect 25872 10208 25924 10260
rect 27988 10208 28040 10260
rect 26332 10072 26384 10124
rect 15660 10004 15712 10056
rect 18236 10004 18288 10056
rect 27160 10115 27212 10124
rect 27160 10081 27169 10115
rect 27169 10081 27203 10115
rect 27203 10081 27212 10115
rect 27160 10072 27212 10081
rect 27344 10115 27396 10124
rect 27344 10081 27353 10115
rect 27353 10081 27387 10115
rect 27387 10081 27396 10115
rect 27344 10072 27396 10081
rect 28540 10208 28592 10260
rect 30012 10183 30064 10192
rect 30012 10149 30021 10183
rect 30021 10149 30055 10183
rect 30055 10149 30064 10183
rect 30012 10140 30064 10149
rect 30840 10208 30892 10260
rect 31392 10208 31444 10260
rect 16580 9936 16632 9988
rect 20536 9936 20588 9988
rect 28264 10004 28316 10056
rect 28080 9936 28132 9988
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 30196 10004 30248 10056
rect 30840 10115 30892 10124
rect 30840 10081 30849 10115
rect 30849 10081 30883 10115
rect 30883 10081 30892 10115
rect 30840 10072 30892 10081
rect 32128 10140 32180 10192
rect 31116 10115 31168 10124
rect 31116 10081 31125 10115
rect 31125 10081 31159 10115
rect 31159 10081 31168 10115
rect 31116 10072 31168 10081
rect 31668 10115 31720 10124
rect 31668 10081 31677 10115
rect 31677 10081 31711 10115
rect 31711 10081 31720 10115
rect 31668 10072 31720 10081
rect 32956 10208 33008 10260
rect 14096 9868 14148 9920
rect 14648 9868 14700 9920
rect 16212 9868 16264 9920
rect 16304 9868 16356 9920
rect 16856 9911 16908 9920
rect 16856 9877 16865 9911
rect 16865 9877 16899 9911
rect 16899 9877 16908 9911
rect 16856 9868 16908 9877
rect 17040 9911 17092 9920
rect 17040 9877 17049 9911
rect 17049 9877 17083 9911
rect 17083 9877 17092 9911
rect 17040 9868 17092 9877
rect 17868 9868 17920 9920
rect 19248 9868 19300 9920
rect 19616 9868 19668 9920
rect 19892 9868 19944 9920
rect 20720 9911 20772 9920
rect 20720 9877 20729 9911
rect 20729 9877 20763 9911
rect 20763 9877 20772 9911
rect 20720 9868 20772 9877
rect 24676 9911 24728 9920
rect 24676 9877 24685 9911
rect 24685 9877 24719 9911
rect 24719 9877 24728 9911
rect 24676 9868 24728 9877
rect 26976 9911 27028 9920
rect 26976 9877 26985 9911
rect 26985 9877 27019 9911
rect 27019 9877 27028 9911
rect 26976 9868 27028 9877
rect 27252 9911 27304 9920
rect 27252 9877 27261 9911
rect 27261 9877 27295 9911
rect 27295 9877 27304 9911
rect 27252 9868 27304 9877
rect 27620 9868 27672 9920
rect 29000 9911 29052 9920
rect 29000 9877 29009 9911
rect 29009 9877 29043 9911
rect 29043 9877 29052 9911
rect 29000 9868 29052 9877
rect 29276 9911 29328 9920
rect 29276 9877 29285 9911
rect 29285 9877 29319 9911
rect 29319 9877 29328 9911
rect 29276 9868 29328 9877
rect 29552 9868 29604 9920
rect 31300 9936 31352 9988
rect 32680 9936 32732 9988
rect 30380 9868 30432 9920
rect 30748 9911 30800 9920
rect 30748 9877 30757 9911
rect 30757 9877 30791 9911
rect 30791 9877 30800 9911
rect 30748 9868 30800 9877
rect 31116 9868 31168 9920
rect 32404 9868 32456 9920
rect 1306 9766 1358 9818
rect 1370 9766 1422 9818
rect 1434 9766 1486 9818
rect 1498 9766 1550 9818
rect 1562 9766 1614 9818
rect 9306 9766 9358 9818
rect 9370 9766 9422 9818
rect 9434 9766 9486 9818
rect 9498 9766 9550 9818
rect 9562 9766 9614 9818
rect 17306 9766 17358 9818
rect 17370 9766 17422 9818
rect 17434 9766 17486 9818
rect 17498 9766 17550 9818
rect 17562 9766 17614 9818
rect 25306 9766 25358 9818
rect 25370 9766 25422 9818
rect 25434 9766 25486 9818
rect 25498 9766 25550 9818
rect 25562 9766 25614 9818
rect 33306 9766 33358 9818
rect 33370 9766 33422 9818
rect 33434 9766 33486 9818
rect 33498 9766 33550 9818
rect 33562 9766 33614 9818
rect 41306 9766 41358 9818
rect 41370 9766 41422 9818
rect 41434 9766 41486 9818
rect 41498 9766 41550 9818
rect 41562 9766 41614 9818
rect 12992 9596 13044 9648
rect 13636 9596 13688 9648
rect 14372 9664 14424 9716
rect 11060 9528 11112 9580
rect 13452 9528 13504 9580
rect 13820 9528 13872 9580
rect 8760 9460 8812 9512
rect 15568 9596 15620 9648
rect 16672 9664 16724 9716
rect 17224 9664 17276 9716
rect 17592 9664 17644 9716
rect 17868 9664 17920 9716
rect 15752 9596 15804 9648
rect 16120 9596 16172 9648
rect 14280 9528 14332 9580
rect 14740 9528 14792 9580
rect 15200 9528 15252 9580
rect 15844 9528 15896 9580
rect 14096 9503 14148 9512
rect 14096 9469 14105 9503
rect 14105 9469 14139 9503
rect 14139 9469 14148 9503
rect 14096 9460 14148 9469
rect 16580 9528 16632 9580
rect 13268 9392 13320 9444
rect 16028 9503 16080 9512
rect 16028 9469 16037 9503
rect 16037 9469 16071 9503
rect 16071 9469 16080 9503
rect 16028 9460 16080 9469
rect 16212 9460 16264 9512
rect 16672 9460 16724 9512
rect 16856 9460 16908 9512
rect 14740 9435 14792 9444
rect 14740 9401 14749 9435
rect 14749 9401 14783 9435
rect 14783 9401 14792 9435
rect 14740 9392 14792 9401
rect 15476 9392 15528 9444
rect 16948 9392 17000 9444
rect 17500 9503 17552 9512
rect 17500 9469 17509 9503
rect 17509 9469 17543 9503
rect 17543 9469 17552 9503
rect 17500 9460 17552 9469
rect 18052 9571 18104 9580
rect 18052 9537 18061 9571
rect 18061 9537 18095 9571
rect 18095 9537 18104 9571
rect 18052 9528 18104 9537
rect 18420 9639 18472 9648
rect 18420 9605 18429 9639
rect 18429 9605 18463 9639
rect 18463 9605 18472 9639
rect 18420 9596 18472 9605
rect 18880 9596 18932 9648
rect 19156 9639 19208 9648
rect 19156 9605 19165 9639
rect 19165 9605 19199 9639
rect 19199 9605 19208 9639
rect 19156 9596 19208 9605
rect 21548 9664 21600 9716
rect 18696 9528 18748 9580
rect 19708 9596 19760 9648
rect 18972 9460 19024 9512
rect 19432 9460 19484 9512
rect 19616 9503 19668 9512
rect 19616 9469 19625 9503
rect 19625 9469 19659 9503
rect 19659 9469 19668 9503
rect 19616 9460 19668 9469
rect 19984 9528 20036 9580
rect 22192 9596 22244 9648
rect 22744 9596 22796 9648
rect 23572 9596 23624 9648
rect 32864 9664 32916 9716
rect 33324 9664 33376 9716
rect 38752 9664 38804 9716
rect 40500 9664 40552 9716
rect 24492 9596 24544 9648
rect 24768 9596 24820 9648
rect 21088 9528 21140 9580
rect 18696 9392 18748 9444
rect 20076 9392 20128 9444
rect 20168 9392 20220 9444
rect 20720 9503 20772 9512
rect 20720 9469 20729 9503
rect 20729 9469 20763 9503
rect 20763 9469 20772 9503
rect 20720 9460 20772 9469
rect 21364 9571 21416 9580
rect 21364 9537 21373 9571
rect 21373 9537 21407 9571
rect 21407 9537 21416 9571
rect 21364 9528 21416 9537
rect 21640 9528 21692 9580
rect 12716 9324 12768 9376
rect 13636 9324 13688 9376
rect 15384 9324 15436 9376
rect 15844 9324 15896 9376
rect 17868 9324 17920 9376
rect 18144 9367 18196 9376
rect 18144 9333 18153 9367
rect 18153 9333 18187 9367
rect 18187 9333 18196 9367
rect 18144 9324 18196 9333
rect 18604 9367 18656 9376
rect 18604 9333 18613 9367
rect 18613 9333 18647 9367
rect 18647 9333 18656 9367
rect 18604 9324 18656 9333
rect 19340 9324 19392 9376
rect 19524 9324 19576 9376
rect 19984 9324 20036 9376
rect 20812 9392 20864 9444
rect 20904 9392 20956 9444
rect 22928 9528 22980 9580
rect 23020 9528 23072 9580
rect 24032 9528 24084 9580
rect 24124 9460 24176 9512
rect 28080 9460 28132 9512
rect 29644 9596 29696 9648
rect 22560 9435 22612 9444
rect 22560 9401 22569 9435
rect 22569 9401 22603 9435
rect 22603 9401 22612 9435
rect 22560 9392 22612 9401
rect 25412 9435 25464 9444
rect 25412 9401 25421 9435
rect 25421 9401 25455 9435
rect 25455 9401 25464 9435
rect 25412 9392 25464 9401
rect 21732 9367 21784 9376
rect 21732 9333 21741 9367
rect 21741 9333 21775 9367
rect 21775 9333 21784 9367
rect 21732 9324 21784 9333
rect 23756 9324 23808 9376
rect 23848 9324 23900 9376
rect 24676 9324 24728 9376
rect 28356 9367 28408 9376
rect 28356 9333 28365 9367
rect 28365 9333 28399 9367
rect 28399 9333 28408 9367
rect 28356 9324 28408 9333
rect 1946 9222 1998 9274
rect 2010 9222 2062 9274
rect 2074 9222 2126 9274
rect 2138 9222 2190 9274
rect 2202 9222 2254 9274
rect 9946 9222 9998 9274
rect 10010 9222 10062 9274
rect 10074 9222 10126 9274
rect 10138 9222 10190 9274
rect 10202 9222 10254 9274
rect 33946 9222 33998 9274
rect 34010 9222 34062 9274
rect 34074 9222 34126 9274
rect 34138 9222 34190 9274
rect 34202 9222 34254 9274
rect 41946 9222 41998 9274
rect 42010 9222 42062 9274
rect 42074 9222 42126 9274
rect 42138 9222 42190 9274
rect 42202 9222 42254 9274
rect 10140 9052 10192 9104
rect 12256 9120 12308 9172
rect 10876 9027 10928 9036
rect 10876 8993 10885 9027
rect 10885 8993 10919 9027
rect 10919 8993 10928 9027
rect 10876 8984 10928 8993
rect 12072 9052 12124 9104
rect 11980 8984 12032 9036
rect 12440 9027 12492 9036
rect 12440 8993 12449 9027
rect 12449 8993 12483 9027
rect 12483 8993 12492 9027
rect 12440 8984 12492 8993
rect 12992 9095 13044 9104
rect 12992 9061 13001 9095
rect 13001 9061 13035 9095
rect 13035 9061 13044 9095
rect 12992 9052 13044 9061
rect 15660 9120 15712 9172
rect 16396 9120 16448 9172
rect 16488 9120 16540 9172
rect 18880 9120 18932 9172
rect 18972 9120 19024 9172
rect 19064 9120 19116 9172
rect 14372 9052 14424 9104
rect 14464 9095 14516 9104
rect 14464 9061 14473 9095
rect 14473 9061 14507 9095
rect 14507 9061 14516 9095
rect 14464 9052 14516 9061
rect 11612 8916 11664 8968
rect 12808 8916 12860 8968
rect 10876 8848 10928 8900
rect 11980 8848 12032 8900
rect 10508 8780 10560 8832
rect 11888 8823 11940 8832
rect 11888 8789 11897 8823
rect 11897 8789 11931 8823
rect 11931 8789 11940 8823
rect 11888 8780 11940 8789
rect 12072 8823 12124 8832
rect 12072 8789 12081 8823
rect 12081 8789 12115 8823
rect 12115 8789 12124 8823
rect 12072 8780 12124 8789
rect 13636 8848 13688 8900
rect 14280 8984 14332 9036
rect 14648 9027 14700 9036
rect 14648 8993 14657 9027
rect 14657 8993 14691 9027
rect 14691 8993 14700 9027
rect 14648 8984 14700 8993
rect 14188 8780 14240 8832
rect 15568 9052 15620 9104
rect 17776 9095 17828 9104
rect 17776 9061 17785 9095
rect 17785 9061 17819 9095
rect 17819 9061 17828 9095
rect 17776 9052 17828 9061
rect 18420 9095 18472 9104
rect 18420 9061 18429 9095
rect 18429 9061 18463 9095
rect 18463 9061 18472 9095
rect 18420 9052 18472 9061
rect 15200 9027 15252 9036
rect 15200 8993 15209 9027
rect 15209 8993 15243 9027
rect 15243 8993 15252 9027
rect 15200 8984 15252 8993
rect 15476 8984 15528 9036
rect 16764 8984 16816 9036
rect 17224 9027 17276 9036
rect 17224 8993 17233 9027
rect 17233 8993 17267 9027
rect 17267 8993 17276 9027
rect 17224 8984 17276 8993
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 17500 8984 17552 9036
rect 18144 8984 18196 9036
rect 19984 9120 20036 9172
rect 19800 9052 19852 9104
rect 20352 9095 20404 9104
rect 20352 9061 20361 9095
rect 20361 9061 20395 9095
rect 20395 9061 20404 9095
rect 20352 9052 20404 9061
rect 19248 9027 19300 9036
rect 19248 8993 19257 9027
rect 19257 8993 19291 9027
rect 19291 8993 19300 9027
rect 19248 8984 19300 8993
rect 19432 8984 19484 9036
rect 19892 9027 19944 9036
rect 19892 8993 19901 9027
rect 19901 8993 19935 9027
rect 19935 8993 19944 9027
rect 19892 8984 19944 8993
rect 20904 9052 20956 9104
rect 20996 9095 21048 9104
rect 20996 9061 21005 9095
rect 21005 9061 21039 9095
rect 21039 9061 21048 9095
rect 20996 9052 21048 9061
rect 22376 9120 22428 9172
rect 20536 9027 20588 9036
rect 20536 8993 20545 9027
rect 20545 8993 20579 9027
rect 20579 8993 20588 9027
rect 20536 8984 20588 8993
rect 21088 8984 21140 9036
rect 21640 9052 21692 9104
rect 22192 9052 22244 9104
rect 21732 8984 21784 9036
rect 22560 9052 22612 9104
rect 23020 9052 23072 9104
rect 23756 9027 23808 9036
rect 23756 8993 23765 9027
rect 23765 8993 23799 9027
rect 23799 8993 23808 9027
rect 23756 8984 23808 8993
rect 25964 9120 26016 9172
rect 24032 9052 24084 9104
rect 24676 9052 24728 9104
rect 24768 9052 24820 9104
rect 26608 9052 26660 9104
rect 15936 8916 15988 8968
rect 17408 8916 17460 8968
rect 17776 8916 17828 8968
rect 16028 8780 16080 8832
rect 16212 8780 16264 8832
rect 17224 8848 17276 8900
rect 17132 8780 17184 8832
rect 20260 8916 20312 8968
rect 22008 8848 22060 8900
rect 23480 8916 23532 8968
rect 23112 8848 23164 8900
rect 23848 8848 23900 8900
rect 25872 8984 25924 9036
rect 24676 8959 24728 8968
rect 24676 8925 24685 8959
rect 24685 8925 24719 8959
rect 24719 8925 24728 8959
rect 24676 8916 24728 8925
rect 25044 8916 25096 8968
rect 27804 9120 27856 9172
rect 28080 8916 28132 8968
rect 19800 8780 19852 8832
rect 20352 8780 20404 8832
rect 23388 8780 23440 8832
rect 23572 8823 23624 8832
rect 23572 8789 23581 8823
rect 23581 8789 23615 8823
rect 23615 8789 23624 8823
rect 23572 8780 23624 8789
rect 26884 8848 26936 8900
rect 26240 8780 26292 8832
rect 26332 8823 26384 8832
rect 26332 8789 26341 8823
rect 26341 8789 26375 8823
rect 26375 8789 26384 8823
rect 26332 8780 26384 8789
rect 26792 8823 26844 8832
rect 26792 8789 26801 8823
rect 26801 8789 26835 8823
rect 26835 8789 26844 8823
rect 26792 8780 26844 8789
rect 1306 8678 1358 8730
rect 1370 8678 1422 8730
rect 1434 8678 1486 8730
rect 1498 8678 1550 8730
rect 1562 8678 1614 8730
rect 9306 8678 9358 8730
rect 9370 8678 9422 8730
rect 9434 8678 9486 8730
rect 9498 8678 9550 8730
rect 9562 8678 9614 8730
rect 41306 8678 41358 8730
rect 41370 8678 41422 8730
rect 41434 8678 41486 8730
rect 41498 8678 41550 8730
rect 41562 8678 41614 8730
rect 6460 8619 6512 8628
rect 6460 8585 6469 8619
rect 6469 8585 6503 8619
rect 6503 8585 6512 8619
rect 6460 8576 6512 8585
rect 7564 8619 7616 8628
rect 7564 8585 7573 8619
rect 7573 8585 7607 8619
rect 7607 8585 7616 8619
rect 7564 8576 7616 8585
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 9864 8576 9916 8628
rect 10600 8576 10652 8628
rect 9036 8508 9088 8560
rect 10508 8508 10560 8560
rect 13912 8576 13964 8628
rect 10140 8483 10192 8492
rect 10140 8449 10149 8483
rect 10149 8449 10183 8483
rect 10183 8449 10192 8483
rect 10140 8440 10192 8449
rect 10692 8483 10744 8492
rect 10692 8449 10701 8483
rect 10701 8449 10735 8483
rect 10735 8449 10744 8483
rect 10692 8440 10744 8449
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 6828 8372 6880 8424
rect 8024 8372 8076 8424
rect 9496 8372 9548 8424
rect 9680 8415 9732 8424
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 11336 8508 11388 8560
rect 12532 8508 12584 8560
rect 15292 8576 15344 8628
rect 16396 8576 16448 8628
rect 17592 8576 17644 8628
rect 11612 8483 11664 8492
rect 11612 8449 11621 8483
rect 11621 8449 11655 8483
rect 11655 8449 11664 8483
rect 11612 8440 11664 8449
rect 12164 8440 12216 8492
rect 9680 8372 9732 8381
rect 11428 8372 11480 8424
rect 11888 8372 11940 8424
rect 12624 8415 12676 8424
rect 12624 8381 12633 8415
rect 12633 8381 12667 8415
rect 12667 8381 12676 8415
rect 12624 8372 12676 8381
rect 13820 8440 13872 8492
rect 14372 8440 14424 8492
rect 14924 8508 14976 8560
rect 15016 8440 15068 8492
rect 16948 8508 17000 8560
rect 18512 8576 18564 8628
rect 19156 8576 19208 8628
rect 19708 8576 19760 8628
rect 21916 8576 21968 8628
rect 22744 8576 22796 8628
rect 5264 8304 5316 8356
rect 6644 8347 6696 8356
rect 6644 8313 6653 8347
rect 6653 8313 6687 8347
rect 6687 8313 6696 8347
rect 6644 8304 6696 8313
rect 6920 8304 6972 8356
rect 8576 8347 8628 8356
rect 8576 8313 8585 8347
rect 8585 8313 8619 8347
rect 8619 8313 8628 8347
rect 8576 8304 8628 8313
rect 5448 8236 5500 8288
rect 6000 8236 6052 8288
rect 6368 8236 6420 8288
rect 10692 8304 10744 8356
rect 14740 8415 14792 8424
rect 14740 8381 14749 8415
rect 14749 8381 14783 8415
rect 14783 8381 14792 8415
rect 14740 8372 14792 8381
rect 15384 8415 15436 8424
rect 15384 8381 15393 8415
rect 15393 8381 15427 8415
rect 15427 8381 15436 8415
rect 15384 8372 15436 8381
rect 16120 8440 16172 8492
rect 16212 8440 16264 8492
rect 13268 8304 13320 8356
rect 13452 8347 13504 8356
rect 13452 8313 13461 8347
rect 13461 8313 13495 8347
rect 13495 8313 13504 8347
rect 13452 8304 13504 8313
rect 14004 8304 14056 8356
rect 10416 8236 10468 8288
rect 15844 8236 15896 8288
rect 16028 8304 16080 8356
rect 16304 8304 16356 8356
rect 16488 8415 16540 8424
rect 16488 8381 16497 8415
rect 16497 8381 16531 8415
rect 16531 8381 16540 8415
rect 16488 8372 16540 8381
rect 16580 8415 16632 8424
rect 16580 8381 16589 8415
rect 16589 8381 16623 8415
rect 16623 8381 16632 8415
rect 16580 8372 16632 8381
rect 17684 8483 17736 8492
rect 17684 8449 17693 8483
rect 17693 8449 17727 8483
rect 17727 8449 17736 8483
rect 17684 8440 17736 8449
rect 20260 8508 20312 8560
rect 17316 8236 17368 8288
rect 17684 8304 17736 8356
rect 17868 8372 17920 8424
rect 20352 8440 20404 8492
rect 21456 8440 21508 8492
rect 22008 8508 22060 8560
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 18604 8372 18656 8424
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 20444 8415 20496 8424
rect 20444 8381 20453 8415
rect 20453 8381 20487 8415
rect 20487 8381 20496 8415
rect 20444 8372 20496 8381
rect 20720 8415 20772 8424
rect 20720 8381 20729 8415
rect 20729 8381 20763 8415
rect 20763 8381 20772 8415
rect 20720 8372 20772 8381
rect 21180 8372 21232 8424
rect 21364 8372 21416 8424
rect 21732 8415 21784 8424
rect 21732 8381 21741 8415
rect 21741 8381 21775 8415
rect 21775 8381 21784 8415
rect 21732 8372 21784 8381
rect 21824 8415 21876 8424
rect 21824 8381 21833 8415
rect 21833 8381 21867 8415
rect 21867 8381 21876 8415
rect 21824 8372 21876 8381
rect 19892 8304 19944 8356
rect 20168 8304 20220 8356
rect 20996 8236 21048 8288
rect 21180 8236 21232 8288
rect 23020 8415 23072 8424
rect 23020 8381 23029 8415
rect 23029 8381 23063 8415
rect 23063 8381 23072 8415
rect 23020 8372 23072 8381
rect 25412 8576 25464 8628
rect 25780 8576 25832 8628
rect 23940 8440 23992 8492
rect 26148 8508 26200 8560
rect 25872 8440 25924 8492
rect 24124 8372 24176 8424
rect 24400 8347 24452 8356
rect 24400 8313 24409 8347
rect 24409 8313 24443 8347
rect 24443 8313 24452 8347
rect 24400 8304 24452 8313
rect 24676 8304 24728 8356
rect 24952 8415 25004 8424
rect 24952 8381 24961 8415
rect 24961 8381 24995 8415
rect 24995 8381 25004 8415
rect 24952 8372 25004 8381
rect 25044 8415 25096 8424
rect 25044 8381 25053 8415
rect 25053 8381 25087 8415
rect 25087 8381 25096 8415
rect 25044 8372 25096 8381
rect 25504 8415 25556 8424
rect 25504 8381 25513 8415
rect 25513 8381 25547 8415
rect 25547 8381 25556 8415
rect 25504 8372 25556 8381
rect 26516 8372 26568 8424
rect 26608 8372 26660 8424
rect 27068 8372 27120 8424
rect 27252 8304 27304 8356
rect 31852 8304 31904 8356
rect 23940 8236 23992 8288
rect 1946 8134 1998 8186
rect 2010 8134 2062 8186
rect 2074 8134 2126 8186
rect 2138 8134 2190 8186
rect 2202 8134 2254 8186
rect 9946 8134 9998 8186
rect 10010 8134 10062 8186
rect 10074 8134 10126 8186
rect 10138 8134 10190 8186
rect 10202 8134 10254 8186
rect 33946 8134 33998 8186
rect 34010 8134 34062 8186
rect 34074 8134 34126 8186
rect 34138 8134 34190 8186
rect 34202 8134 34254 8186
rect 41946 8134 41998 8186
rect 42010 8134 42062 8186
rect 42074 8134 42126 8186
rect 42138 8134 42190 8186
rect 42202 8134 42254 8186
rect 4252 8032 4304 8084
rect 5080 8032 5132 8084
rect 5540 8075 5592 8084
rect 5540 8041 5549 8075
rect 5549 8041 5583 8075
rect 5583 8041 5592 8075
rect 5540 8032 5592 8041
rect 6184 8032 6236 8084
rect 6552 8032 6604 8084
rect 7288 8032 7340 8084
rect 7472 8075 7524 8084
rect 7472 8041 7481 8075
rect 7481 8041 7515 8075
rect 7515 8041 7524 8075
rect 7472 8032 7524 8041
rect 8116 8032 8168 8084
rect 4344 7964 4396 8016
rect 6000 7964 6052 8016
rect 6460 7964 6512 8016
rect 2780 7692 2832 7744
rect 6092 7896 6144 7948
rect 6828 7964 6880 8016
rect 6644 7896 6696 7948
rect 7564 7964 7616 8016
rect 8392 7964 8444 8016
rect 5172 7760 5224 7812
rect 6828 7871 6880 7880
rect 6828 7837 6837 7871
rect 6837 7837 6871 7871
rect 6871 7837 6880 7871
rect 6828 7828 6880 7837
rect 8576 7939 8628 7948
rect 8576 7905 8585 7939
rect 8585 7905 8619 7939
rect 8619 7905 8628 7939
rect 8576 7896 8628 7905
rect 9220 7964 9272 8016
rect 10324 8032 10376 8084
rect 9496 7964 9548 8016
rect 10968 8075 11020 8084
rect 10968 8041 10977 8075
rect 10977 8041 11011 8075
rect 11011 8041 11020 8075
rect 10968 8032 11020 8041
rect 11244 8032 11296 8084
rect 14004 8032 14056 8084
rect 14556 8032 14608 8084
rect 18604 8032 18656 8084
rect 18696 8032 18748 8084
rect 19524 8032 19576 8084
rect 19800 8032 19852 8084
rect 23204 8032 23256 8084
rect 23480 8032 23532 8084
rect 25044 8032 25096 8084
rect 29184 8032 29236 8084
rect 34980 8032 35032 8084
rect 17132 7964 17184 8016
rect 17224 7964 17276 8016
rect 17960 7964 18012 8016
rect 18880 7964 18932 8016
rect 20260 7964 20312 8016
rect 21088 7964 21140 8016
rect 24676 7964 24728 8016
rect 30104 7964 30156 8016
rect 36084 7964 36136 8016
rect 9956 7828 10008 7880
rect 10140 7871 10192 7880
rect 10140 7837 10149 7871
rect 10149 7837 10183 7871
rect 10183 7837 10192 7871
rect 10140 7828 10192 7837
rect 10324 7828 10376 7880
rect 16396 7896 16448 7948
rect 16488 7896 16540 7948
rect 20628 7896 20680 7948
rect 20812 7896 20864 7948
rect 11336 7828 11388 7880
rect 11888 7828 11940 7880
rect 14740 7828 14792 7880
rect 15108 7828 15160 7880
rect 18696 7828 18748 7880
rect 19892 7828 19944 7880
rect 22468 7828 22520 7880
rect 5356 7692 5408 7744
rect 5816 7692 5868 7744
rect 6460 7735 6512 7744
rect 6460 7701 6469 7735
rect 6469 7701 6503 7735
rect 6503 7701 6512 7735
rect 6460 7692 6512 7701
rect 7196 7692 7248 7744
rect 8208 7692 8260 7744
rect 11060 7692 11112 7744
rect 1306 7590 1358 7642
rect 1370 7590 1422 7642
rect 1434 7590 1486 7642
rect 1498 7590 1550 7642
rect 1562 7590 1614 7642
rect 9306 7590 9358 7642
rect 9370 7590 9422 7642
rect 9434 7590 9486 7642
rect 9498 7590 9550 7642
rect 9562 7590 9614 7642
rect 13544 7760 13596 7812
rect 19156 7760 19208 7812
rect 29368 7828 29420 7880
rect 35256 7828 35308 7880
rect 29920 7760 29972 7812
rect 36452 7760 36504 7812
rect 11796 7692 11848 7744
rect 17500 7692 17552 7744
rect 21456 7692 21508 7744
rect 12900 7624 12952 7676
rect 13360 7624 13412 7676
rect 13452 7624 13504 7676
rect 15936 7624 15988 7676
rect 16304 7624 16356 7676
rect 14602 7556 14654 7608
rect 4528 7488 4580 7540
rect 5724 7488 5776 7540
rect 6000 7488 6052 7540
rect 6736 7488 6788 7540
rect 6368 7420 6420 7472
rect 4252 7395 4304 7404
rect 4252 7361 4261 7395
rect 4261 7361 4295 7395
rect 4295 7361 4304 7395
rect 4252 7352 4304 7361
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 4988 7395 5040 7404
rect 4988 7361 4997 7395
rect 4997 7361 5031 7395
rect 5031 7361 5040 7395
rect 4988 7352 5040 7361
rect 5540 7395 5592 7404
rect 5540 7361 5549 7395
rect 5549 7361 5583 7395
rect 5583 7361 5592 7395
rect 5540 7352 5592 7361
rect 5724 7352 5776 7404
rect 4160 7284 4212 7336
rect 3056 7148 3108 7200
rect 4620 7216 4672 7268
rect 4436 7148 4488 7200
rect 5448 7284 5500 7336
rect 6276 7327 6328 7336
rect 6276 7293 6285 7327
rect 6285 7293 6319 7327
rect 6319 7293 6328 7327
rect 6276 7284 6328 7293
rect 6552 7352 6604 7404
rect 7380 7488 7432 7540
rect 9128 7488 9180 7540
rect 7472 7395 7524 7404
rect 7472 7361 7481 7395
rect 7481 7361 7515 7395
rect 7515 7361 7524 7395
rect 7472 7352 7524 7361
rect 8668 7352 8720 7404
rect 10048 7420 10100 7472
rect 11152 7488 11204 7540
rect 12348 7488 12400 7540
rect 15154 7488 15206 7540
rect 13452 7420 13504 7472
rect 6460 7216 6512 7268
rect 7380 7284 7432 7336
rect 8208 7284 8260 7336
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 10692 7352 10744 7404
rect 13544 7352 13596 7404
rect 10140 7284 10192 7336
rect 10968 7284 11020 7336
rect 11060 7284 11112 7336
rect 16626 7556 16678 7608
rect 15568 7488 15620 7540
rect 19754 7556 19806 7608
rect 21594 7556 21646 7608
rect 23572 7692 23624 7744
rect 29552 7692 29604 7744
rect 36176 7692 36228 7744
rect 23802 7556 23854 7608
rect 24952 7556 25004 7608
rect 25826 7556 25878 7608
rect 28402 7556 28454 7608
rect 30840 7556 30892 7608
rect 41306 7590 41358 7642
rect 41370 7590 41422 7642
rect 41434 7590 41486 7642
rect 41498 7590 41550 7642
rect 41562 7590 41614 7642
rect 17730 7488 17782 7540
rect 17960 7488 18012 7540
rect 20122 7488 20174 7540
rect 22008 7488 22060 7540
rect 25274 7488 25326 7540
rect 27298 7488 27350 7540
rect 28954 7488 29006 7540
rect 36360 7488 36412 7540
rect 8116 7148 8168 7200
rect 8300 7191 8352 7200
rect 8300 7157 8309 7191
rect 8309 7157 8343 7191
rect 8343 7157 8352 7191
rect 8300 7148 8352 7157
rect 9036 7148 9088 7200
rect 10140 7148 10192 7200
rect 10692 7148 10744 7200
rect 33324 7395 33376 7404
rect 33324 7361 33333 7395
rect 33333 7361 33367 7395
rect 33367 7361 33376 7395
rect 33324 7352 33376 7361
rect 32312 7284 32364 7336
rect 37648 7148 37700 7200
rect 38384 7148 38436 7200
rect 1946 7046 1998 7098
rect 2010 7046 2062 7098
rect 2074 7046 2126 7098
rect 2138 7046 2190 7098
rect 2202 7046 2254 7098
rect 9946 7046 9998 7098
rect 10010 7046 10062 7098
rect 10074 7046 10126 7098
rect 10138 7046 10190 7098
rect 10202 7046 10254 7098
rect 33946 7046 33998 7098
rect 34010 7046 34062 7098
rect 34074 7046 34126 7098
rect 34138 7046 34190 7098
rect 34202 7046 34254 7098
rect 41946 7046 41998 7098
rect 42010 7046 42062 7098
rect 42074 7046 42126 7098
rect 42138 7046 42190 7098
rect 42202 7046 42254 7098
rect 4528 6987 4580 6996
rect 4528 6953 4537 6987
rect 4537 6953 4571 6987
rect 4571 6953 4580 6987
rect 4528 6944 4580 6953
rect 6000 6987 6052 6996
rect 6000 6953 6009 6987
rect 6009 6953 6043 6987
rect 6043 6953 6052 6987
rect 6000 6944 6052 6953
rect 6276 6944 6328 6996
rect 12348 6944 12400 6996
rect 9312 6876 9364 6928
rect 11244 6876 11296 6928
rect 3884 6740 3936 6792
rect 4620 6740 4672 6792
rect 4896 6783 4948 6792
rect 4896 6749 4905 6783
rect 4905 6749 4939 6783
rect 4939 6749 4948 6783
rect 4896 6740 4948 6749
rect 3332 6672 3384 6724
rect 5632 6808 5684 6860
rect 7012 6851 7064 6860
rect 5080 6740 5132 6792
rect 5724 6783 5776 6792
rect 5724 6749 5733 6783
rect 5733 6749 5767 6783
rect 5767 6749 5776 6783
rect 5724 6740 5776 6749
rect 6276 6783 6328 6792
rect 6276 6749 6285 6783
rect 6285 6749 6319 6783
rect 6319 6749 6328 6783
rect 6276 6740 6328 6749
rect 3608 6604 3660 6656
rect 4160 6647 4212 6656
rect 4160 6613 4169 6647
rect 4169 6613 4203 6647
rect 4203 6613 4212 6647
rect 4160 6604 4212 6613
rect 4804 6604 4856 6656
rect 7012 6817 7021 6851
rect 7021 6817 7055 6851
rect 7055 6817 7064 6851
rect 7012 6808 7064 6817
rect 7104 6783 7156 6792
rect 7104 6749 7113 6783
rect 7113 6749 7147 6783
rect 7147 6749 7156 6783
rect 7104 6740 7156 6749
rect 6828 6672 6880 6724
rect 7840 6808 7892 6860
rect 8760 6851 8812 6860
rect 8760 6817 8769 6851
rect 8769 6817 8803 6851
rect 8803 6817 8812 6851
rect 8760 6808 8812 6817
rect 6644 6604 6696 6656
rect 8852 6783 8904 6792
rect 8852 6749 8861 6783
rect 8861 6749 8895 6783
rect 8895 6749 8904 6783
rect 8852 6740 8904 6749
rect 7748 6672 7800 6724
rect 9496 6851 9548 6860
rect 9496 6817 9505 6851
rect 9505 6817 9539 6851
rect 9539 6817 9548 6851
rect 9496 6808 9548 6817
rect 9128 6740 9180 6792
rect 9956 6808 10008 6860
rect 11152 6851 11204 6860
rect 11152 6817 11161 6851
rect 11161 6817 11195 6851
rect 11195 6817 11204 6851
rect 12900 6876 12952 6928
rect 36084 6876 36136 6928
rect 36452 6876 36504 6928
rect 11152 6808 11204 6817
rect 32864 6851 32916 6860
rect 32864 6817 32873 6851
rect 32873 6817 32907 6851
rect 32907 6817 32916 6851
rect 32864 6808 32916 6817
rect 10140 6783 10192 6792
rect 10140 6749 10149 6783
rect 10149 6749 10183 6783
rect 10183 6749 10192 6783
rect 10140 6740 10192 6749
rect 11704 6740 11756 6792
rect 32496 6740 32548 6792
rect 34612 6851 34664 6860
rect 34612 6817 34621 6851
rect 34621 6817 34655 6851
rect 34655 6817 34664 6851
rect 34612 6808 34664 6817
rect 35624 6740 35676 6792
rect 10416 6672 10468 6724
rect 8944 6604 8996 6656
rect 9864 6604 9916 6656
rect 10508 6604 10560 6656
rect 1306 6502 1358 6554
rect 1370 6502 1422 6554
rect 1434 6502 1486 6554
rect 1498 6502 1550 6554
rect 1562 6502 1614 6554
rect 9306 6502 9358 6554
rect 9370 6502 9422 6554
rect 9434 6502 9486 6554
rect 9498 6502 9550 6554
rect 9562 6502 9614 6554
rect 5632 6443 5684 6452
rect 5632 6409 5641 6443
rect 5641 6409 5675 6443
rect 5675 6409 5684 6443
rect 5632 6400 5684 6409
rect 7840 6443 7892 6452
rect 7840 6409 7849 6443
rect 7849 6409 7883 6443
rect 7883 6409 7892 6443
rect 7840 6400 7892 6409
rect 8668 6400 8720 6452
rect 8852 6400 8904 6452
rect 11336 6400 11388 6452
rect 9772 6332 9824 6384
rect 10508 6332 10560 6384
rect 10784 6332 10836 6384
rect 8944 6239 8996 6248
rect 8944 6205 8953 6239
rect 8953 6205 8987 6239
rect 8987 6205 8996 6239
rect 8944 6196 8996 6205
rect 6368 6128 6420 6180
rect 7380 6171 7432 6180
rect 7380 6137 7389 6171
rect 7389 6137 7423 6171
rect 7423 6137 7432 6171
rect 7380 6128 7432 6137
rect 7472 6128 7524 6180
rect 9588 6128 9640 6180
rect 5540 6060 5592 6112
rect 6828 6060 6880 6112
rect 7748 6060 7800 6112
rect 9220 6060 9272 6112
rect 9956 6060 10008 6112
rect 11520 6332 11572 6384
rect 13084 6604 13136 6656
rect 31484 6604 31536 6656
rect 41306 6502 41358 6554
rect 41370 6502 41422 6554
rect 41434 6502 41486 6554
rect 41498 6502 41550 6554
rect 41562 6502 41614 6554
rect 37924 6400 37976 6452
rect 39856 6400 39908 6452
rect 10784 6239 10836 6248
rect 10784 6205 10793 6239
rect 10793 6205 10827 6239
rect 10827 6205 10836 6239
rect 10784 6196 10836 6205
rect 11520 6060 11572 6112
rect 1946 5958 1998 6010
rect 2010 5958 2062 6010
rect 2074 5958 2126 6010
rect 2138 5958 2190 6010
rect 2202 5958 2254 6010
rect 9946 5958 9998 6010
rect 10010 5958 10062 6010
rect 10074 5958 10126 6010
rect 10138 5958 10190 6010
rect 10202 5958 10254 6010
rect 9772 5899 9824 5908
rect 9772 5865 9781 5899
rect 9781 5865 9815 5899
rect 9815 5865 9824 5899
rect 9772 5856 9824 5865
rect 10416 5856 10468 5908
rect 10508 5899 10560 5908
rect 10508 5865 10517 5899
rect 10517 5865 10551 5899
rect 10551 5865 10560 5899
rect 10508 5856 10560 5865
rect 35992 6264 36044 6316
rect 34888 6239 34940 6248
rect 34888 6205 34897 6239
rect 34897 6205 34931 6239
rect 34931 6205 34940 6239
rect 34888 6196 34940 6205
rect 35624 6239 35676 6248
rect 35624 6205 35633 6239
rect 35633 6205 35667 6239
rect 35667 6205 35676 6239
rect 35624 6196 35676 6205
rect 32864 6103 32916 6112
rect 32864 6069 32873 6103
rect 32873 6069 32907 6103
rect 32907 6069 32916 6103
rect 32864 6060 32916 6069
rect 37004 6060 37056 6112
rect 33946 5958 33998 6010
rect 34010 5958 34062 6010
rect 34074 5958 34126 6010
rect 34138 5958 34190 6010
rect 34202 5958 34254 6010
rect 41946 5958 41998 6010
rect 42010 5958 42062 6010
rect 42074 5958 42126 6010
rect 42138 5958 42190 6010
rect 42202 5958 42254 6010
rect 9864 5788 9916 5840
rect 11336 5788 11388 5840
rect 12072 5788 12124 5840
rect 8944 5720 8996 5772
rect 11888 5720 11940 5772
rect 8576 5584 8628 5636
rect 9588 5584 9640 5636
rect 9128 5516 9180 5568
rect 1306 5414 1358 5466
rect 1370 5414 1422 5466
rect 1434 5414 1486 5466
rect 1498 5414 1550 5466
rect 1562 5414 1614 5466
rect 9306 5414 9358 5466
rect 9370 5414 9422 5466
rect 9434 5414 9486 5466
rect 9498 5414 9550 5466
rect 9562 5414 9614 5466
rect 41306 5414 41358 5466
rect 41370 5414 41422 5466
rect 41434 5414 41486 5466
rect 41498 5414 41550 5466
rect 41562 5414 41614 5466
rect 32128 5176 32180 5228
rect 32588 5108 32640 5160
rect 35992 5151 36044 5160
rect 35992 5117 36001 5151
rect 36001 5117 36035 5151
rect 36035 5117 36044 5151
rect 35992 5108 36044 5117
rect 31944 5040 31996 5092
rect 1946 4870 1998 4922
rect 2010 4870 2062 4922
rect 2074 4870 2126 4922
rect 2138 4870 2190 4922
rect 2202 4870 2254 4922
rect 1306 4326 1358 4378
rect 1370 4326 1422 4378
rect 1434 4326 1486 4378
rect 1498 4326 1550 4378
rect 1562 4326 1614 4378
rect 9306 4326 9358 4378
rect 9370 4326 9422 4378
rect 9434 4326 9486 4378
rect 9498 4326 9550 4378
rect 9562 4326 9614 4378
rect 29920 4360 29972 4412
rect 33692 4972 33744 5024
rect 37280 4972 37332 5024
rect 33946 4870 33998 4922
rect 34010 4870 34062 4922
rect 34074 4870 34126 4922
rect 34138 4870 34190 4922
rect 34202 4870 34254 4922
rect 41946 4870 41998 4922
rect 42010 4870 42062 4922
rect 42074 4870 42126 4922
rect 42138 4870 42190 4922
rect 42202 4870 42254 4922
rect 32772 4675 32824 4684
rect 32772 4641 32781 4675
rect 32781 4641 32815 4675
rect 32815 4641 32824 4675
rect 32772 4632 32824 4641
rect 32956 4632 33008 4684
rect 33232 4675 33284 4684
rect 33232 4641 33241 4675
rect 33241 4641 33275 4675
rect 33275 4641 33284 4675
rect 33232 4632 33284 4641
rect 35164 4675 35216 4684
rect 35164 4641 35173 4675
rect 35173 4641 35207 4675
rect 35207 4641 35216 4675
rect 35164 4632 35216 4641
rect 35900 4564 35952 4616
rect 32956 4428 33008 4480
rect 34336 4471 34388 4480
rect 34336 4437 34345 4471
rect 34345 4437 34379 4471
rect 34379 4437 34388 4471
rect 34336 4428 34388 4437
rect 34888 4428 34940 4480
rect 35624 4471 35676 4480
rect 35624 4437 35633 4471
rect 35633 4437 35667 4471
rect 35667 4437 35676 4471
rect 35624 4428 35676 4437
rect 41306 4326 41358 4378
rect 41370 4326 41422 4378
rect 41434 4326 41486 4378
rect 41498 4326 41550 4378
rect 41562 4326 41614 4378
rect 9864 4156 9916 4208
rect 10876 4156 10928 4208
rect 32864 4088 32916 4140
rect 36084 4224 36136 4276
rect 36912 4224 36964 4276
rect 33048 4156 33100 4208
rect 34520 4199 34572 4208
rect 34520 4165 34529 4199
rect 34529 4165 34563 4199
rect 34563 4165 34572 4199
rect 34520 4156 34572 4165
rect 32680 4020 32732 4072
rect 33416 4063 33468 4072
rect 33416 4029 33425 4063
rect 33425 4029 33459 4063
rect 33459 4029 33468 4063
rect 33416 4020 33468 4029
rect 33508 4063 33560 4072
rect 33508 4029 33517 4063
rect 33517 4029 33551 4063
rect 33551 4029 33560 4063
rect 35348 4088 35400 4140
rect 37924 4088 37976 4140
rect 33508 4020 33560 4029
rect 33784 4020 33836 4072
rect 34428 4020 34480 4072
rect 35900 4063 35952 4072
rect 35900 4029 35909 4063
rect 35909 4029 35943 4063
rect 35943 4029 35952 4063
rect 35900 4020 35952 4029
rect 33876 3952 33928 4004
rect 34796 3952 34848 4004
rect 35808 3952 35860 4004
rect 37740 3952 37792 4004
rect 32036 3884 32088 3936
rect 32680 3884 32732 3936
rect 32956 3884 33008 3936
rect 34612 3884 34664 3936
rect 34704 3927 34756 3936
rect 34704 3893 34713 3927
rect 34713 3893 34747 3927
rect 34747 3893 34756 3927
rect 34704 3884 34756 3893
rect 35164 3927 35216 3936
rect 35164 3893 35173 3927
rect 35173 3893 35207 3927
rect 35207 3893 35216 3927
rect 35164 3884 35216 3893
rect 35440 3927 35492 3936
rect 35440 3893 35449 3927
rect 35449 3893 35483 3927
rect 35483 3893 35492 3927
rect 35440 3884 35492 3893
rect 35900 3884 35952 3936
rect 36360 3884 36412 3936
rect 36728 3927 36780 3936
rect 36728 3893 36737 3927
rect 36737 3893 36771 3927
rect 36771 3893 36780 3927
rect 36728 3884 36780 3893
rect 1946 3782 1998 3834
rect 2010 3782 2062 3834
rect 2074 3782 2126 3834
rect 2138 3782 2190 3834
rect 2202 3782 2254 3834
rect 9946 3782 9998 3834
rect 10010 3782 10062 3834
rect 10074 3782 10126 3834
rect 10138 3782 10190 3834
rect 10202 3782 10254 3834
rect 28356 3816 28408 3868
rect 31852 3816 31904 3868
rect 33946 3782 33998 3834
rect 34010 3782 34062 3834
rect 34074 3782 34126 3834
rect 34138 3782 34190 3834
rect 34202 3782 34254 3834
rect 41946 3782 41998 3834
rect 42010 3782 42062 3834
rect 42074 3782 42126 3834
rect 42138 3782 42190 3834
rect 42202 3782 42254 3834
rect 30472 3680 30524 3732
rect 32864 3680 32916 3732
rect 31300 3612 31352 3664
rect 37096 3680 37148 3732
rect 34704 3612 34756 3664
rect 36452 3612 36504 3664
rect 37832 3612 37884 3664
rect 32956 3587 33008 3596
rect 32956 3553 32965 3587
rect 32965 3553 32999 3587
rect 32999 3553 33008 3587
rect 32956 3544 33008 3553
rect 33600 3544 33652 3596
rect 34060 3544 34112 3596
rect 34152 3544 34204 3596
rect 31116 3476 31168 3528
rect 34336 3476 34388 3528
rect 29828 3408 29880 3460
rect 33784 3408 33836 3460
rect 30380 3340 30432 3392
rect 33324 3340 33376 3392
rect 34060 3340 34112 3392
rect 34796 3587 34848 3596
rect 34796 3553 34805 3587
rect 34805 3553 34839 3587
rect 34839 3553 34848 3587
rect 34796 3544 34848 3553
rect 35348 3587 35400 3596
rect 35348 3553 35357 3587
rect 35357 3553 35391 3587
rect 35391 3553 35400 3587
rect 35348 3544 35400 3553
rect 35440 3544 35492 3596
rect 35808 3544 35860 3596
rect 36544 3544 36596 3596
rect 34612 3476 34664 3528
rect 35532 3476 35584 3528
rect 35256 3408 35308 3460
rect 36084 3476 36136 3528
rect 36176 3408 36228 3460
rect 36728 3408 36780 3460
rect 37372 3544 37424 3596
rect 38568 3544 38620 3596
rect 37648 3476 37700 3528
rect 37188 3408 37240 3460
rect 34612 3383 34664 3392
rect 34612 3349 34621 3383
rect 34621 3349 34655 3383
rect 34655 3349 34664 3383
rect 34612 3340 34664 3349
rect 35808 3340 35860 3392
rect 37464 3340 37516 3392
rect 1306 3238 1358 3290
rect 1370 3238 1422 3290
rect 1434 3238 1486 3290
rect 1498 3238 1550 3290
rect 1562 3238 1614 3290
rect 9306 3238 9358 3290
rect 9370 3238 9422 3290
rect 9434 3238 9486 3290
rect 9498 3238 9550 3290
rect 9562 3238 9614 3290
rect 41306 3238 41358 3290
rect 41370 3238 41422 3290
rect 41434 3238 41486 3290
rect 41498 3238 41550 3290
rect 41562 3238 41614 3290
rect 28080 3000 28132 3052
rect 29828 3043 29880 3052
rect 29828 3009 29837 3043
rect 29837 3009 29871 3043
rect 29871 3009 29880 3043
rect 29828 3000 29880 3009
rect 32220 3068 32272 3120
rect 33784 3179 33836 3188
rect 33784 3145 33793 3179
rect 33793 3145 33827 3179
rect 33827 3145 33836 3179
rect 33784 3136 33836 3145
rect 36360 3136 36412 3188
rect 36544 3136 36596 3188
rect 39028 3136 39080 3188
rect 28172 2932 28224 2984
rect 28448 2975 28500 2984
rect 28448 2941 28457 2975
rect 28457 2941 28491 2975
rect 28491 2941 28500 2975
rect 28448 2932 28500 2941
rect 28724 2975 28776 2984
rect 28724 2941 28733 2975
rect 28733 2941 28767 2975
rect 28767 2941 28776 2975
rect 28724 2932 28776 2941
rect 32036 3000 32088 3052
rect 30380 2975 30432 2984
rect 30380 2941 30389 2975
rect 30389 2941 30423 2975
rect 30423 2941 30432 2975
rect 30380 2932 30432 2941
rect 30656 2975 30708 2984
rect 30656 2941 30665 2975
rect 30665 2941 30699 2975
rect 30699 2941 30708 2975
rect 30656 2932 30708 2941
rect 31668 2932 31720 2984
rect 31852 2932 31904 2984
rect 32404 3000 32456 3052
rect 33324 3000 33376 3052
rect 33968 3068 34020 3120
rect 36084 3068 36136 3120
rect 37188 3068 37240 3120
rect 34888 3000 34940 3052
rect 36360 3000 36412 3052
rect 24768 2864 24820 2916
rect 26332 2864 26384 2916
rect 29092 2864 29144 2916
rect 31484 2864 31536 2916
rect 33232 2975 33284 2984
rect 33232 2941 33241 2975
rect 33241 2941 33275 2975
rect 33275 2941 33284 2975
rect 33232 2932 33284 2941
rect 34612 2932 34664 2984
rect 34980 2932 35032 2984
rect 35624 2975 35676 2984
rect 35624 2941 35633 2975
rect 35633 2941 35667 2975
rect 35667 2941 35676 2975
rect 35624 2932 35676 2941
rect 35808 2932 35860 2984
rect 25964 2839 26016 2848
rect 25964 2805 25973 2839
rect 25973 2805 26007 2839
rect 26007 2805 26016 2839
rect 25964 2796 26016 2805
rect 27988 2839 28040 2848
rect 27988 2805 27997 2839
rect 27997 2805 28031 2839
rect 28031 2805 28040 2839
rect 27988 2796 28040 2805
rect 30380 2796 30432 2848
rect 30564 2796 30616 2848
rect 31300 2796 31352 2848
rect 32956 2796 33008 2848
rect 35072 2864 35124 2916
rect 37464 3043 37516 3052
rect 37464 3009 37473 3043
rect 37473 3009 37507 3043
rect 37507 3009 37516 3043
rect 37464 3000 37516 3009
rect 37188 2975 37240 2984
rect 37188 2941 37197 2975
rect 37197 2941 37231 2975
rect 37231 2941 37240 2975
rect 37188 2932 37240 2941
rect 38016 3068 38068 3120
rect 38108 2932 38160 2984
rect 38200 2864 38252 2916
rect 34336 2796 34388 2848
rect 37740 2796 37792 2848
rect 38016 2796 38068 2848
rect 38844 2839 38896 2848
rect 38844 2805 38853 2839
rect 38853 2805 38887 2839
rect 38887 2805 38896 2839
rect 38844 2796 38896 2805
rect 1946 2694 1998 2746
rect 2010 2694 2062 2746
rect 2074 2694 2126 2746
rect 2138 2694 2190 2746
rect 2202 2694 2254 2746
rect 9946 2694 9998 2746
rect 10010 2694 10062 2746
rect 10074 2694 10126 2746
rect 10138 2694 10190 2746
rect 10202 2694 10254 2746
rect 33946 2694 33998 2746
rect 34010 2694 34062 2746
rect 34074 2694 34126 2746
rect 34138 2694 34190 2746
rect 34202 2694 34254 2746
rect 41946 2694 41998 2746
rect 42010 2694 42062 2746
rect 42074 2694 42126 2746
rect 42138 2694 42190 2746
rect 42202 2694 42254 2746
rect 27620 2592 27672 2644
rect 24860 2524 24912 2576
rect 27988 2524 28040 2576
rect 29828 2592 29880 2644
rect 31300 2592 31352 2644
rect 31392 2592 31444 2644
rect 34520 2592 34572 2644
rect 30472 2524 30524 2576
rect 25136 2456 25188 2508
rect 27712 2499 27764 2508
rect 27712 2465 27721 2499
rect 27721 2465 27755 2499
rect 27755 2465 27764 2499
rect 27712 2456 27764 2465
rect 29000 2499 29052 2508
rect 29000 2465 29009 2499
rect 29009 2465 29043 2499
rect 29043 2465 29052 2499
rect 29000 2456 29052 2465
rect 29092 2456 29144 2508
rect 24308 2388 24360 2440
rect 26884 2388 26936 2440
rect 30564 2456 30616 2508
rect 31576 2524 31628 2576
rect 32956 2524 33008 2576
rect 39120 2592 39172 2644
rect 31024 2499 31076 2508
rect 31024 2465 31033 2499
rect 31033 2465 31067 2499
rect 31067 2465 31076 2499
rect 31024 2456 31076 2465
rect 31484 2499 31536 2508
rect 31484 2465 31493 2499
rect 31493 2465 31527 2499
rect 31527 2465 31536 2499
rect 31484 2456 31536 2465
rect 30472 2388 30524 2440
rect 31668 2388 31720 2440
rect 32128 2388 32180 2440
rect 33600 2388 33652 2440
rect 31484 2320 31536 2372
rect 36544 2524 36596 2576
rect 34704 2456 34756 2508
rect 35900 2499 35952 2508
rect 35900 2465 35909 2499
rect 35909 2465 35943 2499
rect 35943 2465 35952 2499
rect 35900 2456 35952 2465
rect 34796 2388 34848 2440
rect 37280 2499 37332 2508
rect 37280 2465 37289 2499
rect 37289 2465 37323 2499
rect 37323 2465 37332 2499
rect 37280 2456 37332 2465
rect 37464 2499 37516 2508
rect 37464 2465 37473 2499
rect 37473 2465 37507 2499
rect 37507 2465 37516 2499
rect 37464 2456 37516 2465
rect 37556 2456 37608 2508
rect 38108 2499 38160 2508
rect 38108 2465 38117 2499
rect 38117 2465 38151 2499
rect 38151 2465 38160 2499
rect 38108 2456 38160 2465
rect 38844 2524 38896 2576
rect 38476 2456 38528 2508
rect 40684 2456 40736 2508
rect 34612 2320 34664 2372
rect 26056 2295 26108 2304
rect 26056 2261 26065 2295
rect 26065 2261 26099 2295
rect 26099 2261 26108 2295
rect 26056 2252 26108 2261
rect 31024 2252 31076 2304
rect 31852 2252 31904 2304
rect 32128 2252 32180 2304
rect 35164 2252 35216 2304
rect 36820 2320 36872 2372
rect 38568 2388 38620 2440
rect 38660 2320 38712 2372
rect 39120 2388 39172 2440
rect 39580 2320 39632 2372
rect 39212 2252 39264 2304
rect 39672 2295 39724 2304
rect 39672 2261 39681 2295
rect 39681 2261 39715 2295
rect 39715 2261 39724 2295
rect 39672 2252 39724 2261
rect 39764 2252 39816 2304
rect 40500 2295 40552 2304
rect 40500 2261 40509 2295
rect 40509 2261 40543 2295
rect 40543 2261 40552 2295
rect 40500 2252 40552 2261
rect 1306 2150 1358 2202
rect 1370 2150 1422 2202
rect 1434 2150 1486 2202
rect 1498 2150 1550 2202
rect 1562 2150 1614 2202
rect 9306 2150 9358 2202
rect 9370 2150 9422 2202
rect 9434 2150 9486 2202
rect 9498 2150 9550 2202
rect 9562 2150 9614 2202
rect 17306 2150 17358 2202
rect 17370 2150 17422 2202
rect 17434 2150 17486 2202
rect 17498 2150 17550 2202
rect 17562 2150 17614 2202
rect 25306 2150 25358 2202
rect 25370 2150 25422 2202
rect 25434 2150 25486 2202
rect 25498 2150 25550 2202
rect 25562 2150 25614 2202
rect 33306 2150 33358 2202
rect 33370 2150 33422 2202
rect 33434 2150 33486 2202
rect 33498 2150 33550 2202
rect 33562 2150 33614 2202
rect 41306 2150 41358 2202
rect 41370 2150 41422 2202
rect 41434 2150 41486 2202
rect 41498 2150 41550 2202
rect 41562 2150 41614 2202
rect 28172 2048 28224 2100
rect 28448 2048 28500 2100
rect 32772 2048 32824 2100
rect 25964 1980 26016 2032
rect 26424 1980 26476 2032
rect 29092 1980 29144 2032
rect 31668 1980 31720 2032
rect 24584 1912 24636 1964
rect 26056 1912 26108 1964
rect 28724 1912 28776 1964
rect 25044 1887 25096 1896
rect 25044 1853 25053 1887
rect 25053 1853 25087 1887
rect 25087 1853 25096 1887
rect 25044 1844 25096 1853
rect 25596 1844 25648 1896
rect 26792 1887 26844 1896
rect 26792 1853 26801 1887
rect 26801 1853 26835 1887
rect 26835 1853 26844 1887
rect 26792 1844 26844 1853
rect 28264 1887 28316 1896
rect 28264 1853 28273 1887
rect 28273 1853 28307 1887
rect 28307 1853 28316 1887
rect 28264 1844 28316 1853
rect 28540 1887 28592 1896
rect 28540 1853 28549 1887
rect 28549 1853 28583 1887
rect 28583 1853 28592 1887
rect 28540 1844 28592 1853
rect 28632 1844 28684 1896
rect 23756 1776 23808 1828
rect 27896 1819 27948 1828
rect 27896 1785 27905 1819
rect 27905 1785 27939 1819
rect 27939 1785 27948 1819
rect 27896 1776 27948 1785
rect 27068 1708 27120 1760
rect 29920 1776 29972 1828
rect 30288 1887 30340 1896
rect 30288 1853 30297 1887
rect 30297 1853 30331 1887
rect 30331 1853 30340 1887
rect 30288 1844 30340 1853
rect 30380 1887 30432 1896
rect 30380 1853 30389 1887
rect 30389 1853 30423 1887
rect 30423 1853 30432 1887
rect 30380 1844 30432 1853
rect 30840 1912 30892 1964
rect 31944 1912 31996 1964
rect 34520 2048 34572 2100
rect 36728 2048 36780 2100
rect 35164 1980 35216 2032
rect 33048 1955 33100 1964
rect 33048 1921 33057 1955
rect 33057 1921 33091 1955
rect 33091 1921 33100 1955
rect 33048 1912 33100 1921
rect 33324 1955 33376 1964
rect 33324 1921 33333 1955
rect 33333 1921 33367 1955
rect 33367 1921 33376 1955
rect 33324 1912 33376 1921
rect 31392 1819 31444 1828
rect 31392 1785 31401 1819
rect 31401 1785 31435 1819
rect 31435 1785 31444 1819
rect 31392 1776 31444 1785
rect 31852 1887 31904 1896
rect 31852 1853 31861 1887
rect 31861 1853 31895 1887
rect 31895 1853 31904 1887
rect 31852 1844 31904 1853
rect 34428 1912 34480 1964
rect 34612 1955 34664 1964
rect 34612 1921 34621 1955
rect 34621 1921 34655 1955
rect 34655 1921 34664 1955
rect 34612 1912 34664 1921
rect 33968 1844 34020 1896
rect 33784 1776 33836 1828
rect 35532 1887 35584 1896
rect 35532 1853 35541 1887
rect 35541 1853 35575 1887
rect 35575 1853 35584 1887
rect 35532 1844 35584 1853
rect 36636 1912 36688 1964
rect 38476 1980 38528 2032
rect 39580 2091 39632 2100
rect 39580 2057 39589 2091
rect 39589 2057 39623 2091
rect 39623 2057 39632 2091
rect 39580 2048 39632 2057
rect 40224 2048 40276 2100
rect 38752 1980 38804 2032
rect 39488 1980 39540 2032
rect 39764 1980 39816 2032
rect 35716 1844 35768 1896
rect 37556 1776 37608 1828
rect 29276 1708 29328 1760
rect 37832 1887 37884 1896
rect 37832 1853 37841 1887
rect 37841 1853 37875 1887
rect 37875 1853 37884 1887
rect 37832 1844 37884 1853
rect 38384 1844 38436 1896
rect 38660 1889 38712 1896
rect 38660 1855 38669 1889
rect 38669 1855 38703 1889
rect 38703 1855 38712 1889
rect 38660 1844 38712 1855
rect 39304 1844 39356 1896
rect 39396 1844 39448 1896
rect 40132 1844 40184 1896
rect 40868 1844 40920 1896
rect 38568 1708 38620 1760
rect 38752 1751 38804 1760
rect 38752 1717 38761 1751
rect 38761 1717 38795 1751
rect 38795 1717 38804 1751
rect 38752 1708 38804 1717
rect 39212 1708 39264 1760
rect 39856 1776 39908 1828
rect 40408 1708 40460 1760
rect 40776 1708 40828 1760
rect 1946 1606 1998 1658
rect 2010 1606 2062 1658
rect 2074 1606 2126 1658
rect 2138 1606 2190 1658
rect 2202 1606 2254 1658
rect 9946 1606 9998 1658
rect 10010 1606 10062 1658
rect 10074 1606 10126 1658
rect 10138 1606 10190 1658
rect 10202 1606 10254 1658
rect 17946 1606 17998 1658
rect 18010 1606 18062 1658
rect 18074 1606 18126 1658
rect 18138 1606 18190 1658
rect 18202 1606 18254 1658
rect 25946 1606 25998 1658
rect 26010 1606 26062 1658
rect 26074 1606 26126 1658
rect 26138 1606 26190 1658
rect 26202 1606 26254 1658
rect 33946 1606 33998 1658
rect 34010 1606 34062 1658
rect 34074 1606 34126 1658
rect 34138 1606 34190 1658
rect 34202 1606 34254 1658
rect 41946 1606 41998 1658
rect 42010 1606 42062 1658
rect 42074 1606 42126 1658
rect 42138 1606 42190 1658
rect 42202 1606 42254 1658
rect 25136 1547 25188 1556
rect 25136 1513 25145 1547
rect 25145 1513 25179 1547
rect 25179 1513 25188 1547
rect 25136 1504 25188 1513
rect 26792 1504 26844 1556
rect 30104 1504 30156 1556
rect 23572 1411 23624 1420
rect 23572 1377 23581 1411
rect 23581 1377 23615 1411
rect 23615 1377 23624 1411
rect 23572 1368 23624 1377
rect 25228 1411 25280 1420
rect 25228 1377 25237 1411
rect 25237 1377 25271 1411
rect 25271 1377 25280 1411
rect 25228 1368 25280 1377
rect 25688 1411 25740 1420
rect 25688 1377 25697 1411
rect 25697 1377 25731 1411
rect 25731 1377 25740 1411
rect 25688 1368 25740 1377
rect 25780 1368 25832 1420
rect 26424 1436 26476 1488
rect 29368 1436 29420 1488
rect 34060 1504 34112 1556
rect 39212 1504 39264 1556
rect 21548 1300 21600 1352
rect 22560 1300 22612 1352
rect 23480 1300 23532 1352
rect 25964 1300 26016 1352
rect 27436 1411 27488 1420
rect 27436 1377 27445 1411
rect 27445 1377 27479 1411
rect 27479 1377 27488 1411
rect 27436 1368 27488 1377
rect 27988 1411 28040 1420
rect 27988 1377 27997 1411
rect 27997 1377 28031 1411
rect 28031 1377 28040 1411
rect 27988 1368 28040 1377
rect 29276 1411 29328 1420
rect 29276 1377 29285 1411
rect 29285 1377 29319 1411
rect 29319 1377 29328 1411
rect 29276 1368 29328 1377
rect 25780 1232 25832 1284
rect 26516 1232 26568 1284
rect 30840 1411 30892 1420
rect 30840 1377 30849 1411
rect 30849 1377 30883 1411
rect 30883 1377 30892 1411
rect 30840 1368 30892 1377
rect 31024 1368 31076 1420
rect 32036 1368 32088 1420
rect 30748 1343 30800 1352
rect 30748 1309 30757 1343
rect 30757 1309 30791 1343
rect 30791 1309 30800 1343
rect 30748 1300 30800 1309
rect 23756 1164 23808 1216
rect 31208 1232 31260 1284
rect 32772 1300 32824 1352
rect 36360 1436 36412 1488
rect 34244 1368 34296 1420
rect 34060 1300 34112 1352
rect 34336 1300 34388 1352
rect 36728 1436 36780 1488
rect 36912 1436 36964 1488
rect 36636 1411 36688 1420
rect 36636 1377 36645 1411
rect 36645 1377 36679 1411
rect 36679 1377 36688 1411
rect 36636 1368 36688 1377
rect 36820 1368 36872 1420
rect 36268 1300 36320 1352
rect 37556 1368 37608 1420
rect 37924 1368 37976 1420
rect 38200 1368 38252 1420
rect 39764 1436 39816 1488
rect 39120 1411 39172 1420
rect 39120 1377 39129 1411
rect 39129 1377 39163 1411
rect 39163 1377 39172 1411
rect 39120 1368 39172 1377
rect 40040 1504 40092 1556
rect 41144 1436 41196 1488
rect 40040 1411 40092 1420
rect 40040 1377 40049 1411
rect 40049 1377 40083 1411
rect 40083 1377 40092 1411
rect 40040 1368 40092 1377
rect 40500 1411 40552 1420
rect 40500 1377 40509 1411
rect 40509 1377 40543 1411
rect 40543 1377 40552 1411
rect 40500 1368 40552 1377
rect 35716 1232 35768 1284
rect 38660 1343 38712 1352
rect 38660 1309 38669 1343
rect 38669 1309 38703 1343
rect 38703 1309 38712 1343
rect 38660 1300 38712 1309
rect 40132 1300 40184 1352
rect 40408 1232 40460 1284
rect 40960 1232 41012 1284
rect 36360 1164 36412 1216
rect 36728 1207 36780 1216
rect 36728 1173 36737 1207
rect 36737 1173 36771 1207
rect 36771 1173 36780 1207
rect 36728 1164 36780 1173
rect 36820 1164 36872 1216
rect 39304 1164 39356 1216
rect 39948 1164 40000 1216
rect 41328 1232 41380 1284
rect 41972 1207 42024 1216
rect 41972 1173 41981 1207
rect 41981 1173 42015 1207
rect 42015 1173 42024 1207
rect 41972 1164 42024 1173
rect 1306 1062 1358 1114
rect 1370 1062 1422 1114
rect 1434 1062 1486 1114
rect 1498 1062 1550 1114
rect 1562 1062 1614 1114
rect 9306 1062 9358 1114
rect 9370 1062 9422 1114
rect 9434 1062 9486 1114
rect 9498 1062 9550 1114
rect 9562 1062 9614 1114
rect 17306 1062 17358 1114
rect 17370 1062 17422 1114
rect 17434 1062 17486 1114
rect 17498 1062 17550 1114
rect 17562 1062 17614 1114
rect 25306 1062 25358 1114
rect 25370 1062 25422 1114
rect 25434 1062 25486 1114
rect 25498 1062 25550 1114
rect 25562 1062 25614 1114
rect 33306 1062 33358 1114
rect 33370 1062 33422 1114
rect 33434 1062 33486 1114
rect 33498 1062 33550 1114
rect 33562 1062 33614 1114
rect 41306 1062 41358 1114
rect 41370 1062 41422 1114
rect 41434 1062 41486 1114
rect 41498 1062 41550 1114
rect 41562 1062 41614 1114
rect 23572 960 23624 1012
rect 25044 960 25096 1012
rect 25688 960 25740 1012
rect 27712 960 27764 1012
rect 27988 960 28040 1012
rect 30288 960 30340 1012
rect 31208 1003 31260 1012
rect 31208 969 31217 1003
rect 31217 969 31251 1003
rect 31251 969 31260 1003
rect 31208 960 31260 969
rect 32220 960 32272 1012
rect 36360 1003 36412 1012
rect 36360 969 36369 1003
rect 36369 969 36403 1003
rect 36403 969 36412 1003
rect 36360 960 36412 969
rect 38660 960 38712 1012
rect 23480 892 23532 944
rect 29000 892 29052 944
rect 30840 892 30892 944
rect 34612 892 34664 944
rect 36728 892 36780 944
rect 23204 824 23256 876
rect 24952 824 25004 876
rect 23296 799 23348 808
rect 23296 765 23305 799
rect 23305 765 23339 799
rect 23339 765 23348 799
rect 23296 756 23348 765
rect 23664 756 23716 808
rect 25228 799 25280 808
rect 25228 765 25237 799
rect 25237 765 25271 799
rect 25271 765 25280 799
rect 25228 756 25280 765
rect 24032 688 24084 740
rect 24768 688 24820 740
rect 27344 824 27396 876
rect 25872 756 25924 808
rect 27804 799 27856 808
rect 27804 765 27813 799
rect 27813 765 27847 799
rect 27847 765 27856 799
rect 27804 756 27856 765
rect 28080 799 28132 808
rect 28080 765 28089 799
rect 28089 765 28123 799
rect 28123 765 28132 799
rect 28080 756 28132 765
rect 28356 799 28408 808
rect 28356 765 28365 799
rect 28365 765 28399 799
rect 28399 765 28408 799
rect 28356 756 28408 765
rect 30380 799 30432 808
rect 30380 765 30389 799
rect 30389 765 30423 799
rect 30423 765 30432 799
rect 30380 756 30432 765
rect 30656 799 30708 808
rect 30656 765 30665 799
rect 30665 765 30699 799
rect 30699 765 30708 799
rect 30656 756 30708 765
rect 30932 799 30984 808
rect 30932 765 30941 799
rect 30941 765 30975 799
rect 30975 765 30984 799
rect 30932 756 30984 765
rect 27896 688 27948 740
rect 25872 620 25924 672
rect 33784 824 33836 876
rect 32956 799 33008 808
rect 32956 765 32965 799
rect 32965 765 32999 799
rect 32999 765 33008 799
rect 32956 756 33008 765
rect 33692 756 33744 808
rect 33968 756 34020 808
rect 29552 620 29604 672
rect 35256 731 35308 740
rect 35256 697 35265 731
rect 35265 697 35299 731
rect 35299 697 35308 731
rect 35256 688 35308 697
rect 35992 756 36044 808
rect 36268 799 36320 808
rect 36268 765 36277 799
rect 36277 765 36311 799
rect 36311 765 36320 799
rect 36268 756 36320 765
rect 36452 756 36504 808
rect 37648 756 37700 808
rect 37464 688 37516 740
rect 38568 756 38620 808
rect 38936 756 38988 808
rect 39304 799 39356 808
rect 39304 765 39313 799
rect 39313 765 39347 799
rect 39347 765 39356 799
rect 39304 756 39356 765
rect 40040 824 40092 876
rect 40316 892 40368 944
rect 40776 892 40828 944
rect 41236 960 41288 1012
rect 41788 1003 41840 1012
rect 41788 969 41797 1003
rect 41797 969 41831 1003
rect 41831 969 41840 1003
rect 41788 960 41840 969
rect 40408 799 40460 808
rect 40408 765 40417 799
rect 40417 765 40451 799
rect 40451 765 40460 799
rect 40408 756 40460 765
rect 40500 799 40552 808
rect 40500 765 40509 799
rect 40509 765 40543 799
rect 40543 765 40552 799
rect 40500 756 40552 765
rect 40684 799 40736 808
rect 40684 765 40693 799
rect 40693 765 40727 799
rect 40727 765 40736 799
rect 40684 756 40736 765
rect 41052 867 41104 876
rect 41052 833 41061 867
rect 41061 833 41095 867
rect 41095 833 41104 867
rect 41052 824 41104 833
rect 41972 824 42024 876
rect 41328 756 41380 808
rect 42340 799 42392 808
rect 42340 765 42349 799
rect 42349 765 42383 799
rect 42383 765 42392 799
rect 42340 756 42392 765
rect 39028 620 39080 672
rect 40408 620 40460 672
rect 40776 663 40828 672
rect 40776 629 40785 663
rect 40785 629 40819 663
rect 40819 629 40828 663
rect 40776 620 40828 629
rect 41512 663 41564 672
rect 41512 629 41521 663
rect 41521 629 41555 663
rect 41555 629 41564 663
rect 41512 620 41564 629
rect 41788 620 41840 672
rect 1946 518 1998 570
rect 2010 518 2062 570
rect 2074 518 2126 570
rect 2138 518 2190 570
rect 2202 518 2254 570
rect 9946 518 9998 570
rect 10010 518 10062 570
rect 10074 518 10126 570
rect 10138 518 10190 570
rect 10202 518 10254 570
rect 17946 518 17998 570
rect 18010 518 18062 570
rect 18074 518 18126 570
rect 18138 518 18190 570
rect 18202 518 18254 570
rect 25946 518 25998 570
rect 26010 518 26062 570
rect 26074 518 26126 570
rect 26138 518 26190 570
rect 26202 518 26254 570
rect 33946 518 33998 570
rect 34010 518 34062 570
rect 34074 518 34126 570
rect 34138 518 34190 570
rect 34202 518 34254 570
rect 41946 518 41998 570
rect 42010 518 42062 570
rect 42074 518 42126 570
rect 42138 518 42190 570
rect 42202 518 42254 570
rect 25228 416 25280 468
rect 27804 416 27856 468
rect 27988 416 28040 468
rect 28632 416 28684 468
rect 33876 416 33928 468
rect 34428 416 34480 468
rect 38200 416 38252 468
rect 38844 416 38896 468
rect 24952 348 25004 400
rect 27436 348 27488 400
rect 31300 348 31352 400
rect 37464 348 37516 400
rect 39948 416 40000 468
rect 40408 416 40460 468
rect 41052 416 41104 468
rect 39028 348 39080 400
rect 40776 348 40828 400
rect 35256 280 35308 332
rect 41512 280 41564 332
rect 40684 212 40736 264
rect 41236 212 41288 264
rect 38292 144 38344 196
rect 40960 144 41012 196
rect 39304 76 39356 128
rect 41788 212 41840 264
rect 38568 8 38620 60
rect 40224 8 40276 60
<< metal2 >>
rect 5078 11600 5134 12000
rect 5354 11600 5410 12000
rect 5630 11600 5686 12000
rect 5906 11600 5962 12000
rect 6182 11600 6238 12000
rect 6458 11600 6514 12000
rect 6734 11600 6790 12000
rect 7010 11600 7066 12000
rect 7286 11600 7342 12000
rect 7562 11600 7618 12000
rect 7838 11600 7894 12000
rect 8114 11600 8170 12000
rect 8390 11600 8446 12000
rect 8666 11600 8722 12000
rect 8942 11600 8998 12000
rect 9218 11600 9274 12000
rect 9494 11600 9550 12000
rect 9770 11600 9826 12000
rect 10046 11600 10102 12000
rect 10322 11600 10378 12000
rect 10598 11600 10654 12000
rect 10874 11600 10930 12000
rect 11150 11600 11206 12000
rect 11426 11600 11482 12000
rect 11702 11600 11758 12000
rect 11978 11600 12034 12000
rect 12254 11600 12310 12000
rect 12530 11600 12586 12000
rect 12806 11600 12862 12000
rect 13082 11600 13138 12000
rect 13358 11600 13414 12000
rect 13634 11600 13690 12000
rect 13910 11600 13966 12000
rect 14186 11600 14242 12000
rect 14462 11600 14518 12000
rect 14738 11600 14794 12000
rect 15014 11600 15070 12000
rect 15290 11600 15346 12000
rect 15566 11600 15622 12000
rect 15842 11600 15898 12000
rect 16118 11600 16174 12000
rect 16394 11600 16450 12000
rect 16670 11600 16726 12000
rect 16946 11600 17002 12000
rect 17222 11600 17278 12000
rect 17498 11600 17554 12000
rect 17774 11600 17830 12000
rect 18050 11600 18106 12000
rect 18326 11600 18382 12000
rect 18602 11600 18658 12000
rect 18878 11600 18934 12000
rect 19154 11600 19210 12000
rect 19430 11600 19486 12000
rect 19706 11600 19762 12000
rect 19982 11600 20038 12000
rect 20258 11600 20314 12000
rect 20534 11600 20590 12000
rect 20810 11600 20866 12000
rect 21086 11600 21142 12000
rect 21362 11600 21418 12000
rect 21638 11600 21694 12000
rect 21914 11600 21970 12000
rect 22190 11600 22246 12000
rect 22466 11600 22522 12000
rect 22742 11600 22798 12000
rect 23018 11600 23074 12000
rect 23294 11600 23350 12000
rect 23570 11600 23626 12000
rect 23846 11600 23902 12000
rect 24122 11600 24178 12000
rect 24398 11600 24454 12000
rect 24674 11600 24730 12000
rect 24950 11600 25006 12000
rect 25226 11600 25282 12000
rect 25502 11600 25558 12000
rect 25778 11600 25834 12000
rect 26054 11600 26110 12000
rect 26330 11600 26386 12000
rect 26606 11600 26662 12000
rect 26882 11600 26938 12000
rect 27158 11600 27214 12000
rect 27434 11600 27490 12000
rect 27710 11600 27766 12000
rect 27986 11600 28042 12000
rect 28262 11600 28318 12000
rect 28538 11600 28594 12000
rect 28814 11600 28870 12000
rect 29090 11600 29146 12000
rect 29366 11600 29422 12000
rect 29642 11600 29698 12000
rect 29918 11600 29974 12000
rect 30194 11600 30250 12000
rect 30470 11600 30526 12000
rect 30746 11600 30802 12000
rect 31022 11600 31078 12000
rect 31298 11600 31354 12000
rect 31574 11600 31630 12000
rect 31760 11620 31812 11626
rect 1946 11452 2254 11461
rect 1946 11450 1952 11452
rect 2008 11450 2032 11452
rect 2088 11450 2112 11452
rect 2168 11450 2192 11452
rect 2248 11450 2254 11452
rect 2008 11398 2010 11450
rect 2190 11398 2192 11450
rect 1946 11396 1952 11398
rect 2008 11396 2032 11398
rect 2088 11396 2112 11398
rect 2168 11396 2192 11398
rect 2248 11396 2254 11398
rect 1946 11387 2254 11396
rect 1306 10908 1614 10917
rect 1306 10906 1312 10908
rect 1368 10906 1392 10908
rect 1448 10906 1472 10908
rect 1528 10906 1552 10908
rect 1608 10906 1614 10908
rect 1368 10854 1370 10906
rect 1550 10854 1552 10906
rect 1306 10852 1312 10854
rect 1368 10852 1392 10854
rect 1448 10852 1472 10854
rect 1528 10852 1552 10854
rect 1608 10852 1614 10854
rect 1306 10843 1614 10852
rect 1946 10364 2254 10373
rect 1946 10362 1952 10364
rect 2008 10362 2032 10364
rect 2088 10362 2112 10364
rect 2168 10362 2192 10364
rect 2248 10362 2254 10364
rect 2008 10310 2010 10362
rect 2190 10310 2192 10362
rect 1946 10308 1952 10310
rect 2008 10308 2032 10310
rect 2088 10308 2112 10310
rect 2168 10308 2192 10310
rect 2248 10308 2254 10310
rect 1946 10299 2254 10308
rect 1306 9820 1614 9829
rect 1306 9818 1312 9820
rect 1368 9818 1392 9820
rect 1448 9818 1472 9820
rect 1528 9818 1552 9820
rect 1608 9818 1614 9820
rect 1368 9766 1370 9818
rect 1550 9766 1552 9818
rect 1306 9764 1312 9766
rect 1368 9764 1392 9766
rect 1448 9764 1472 9766
rect 1528 9764 1552 9766
rect 1608 9764 1614 9766
rect 1306 9755 1614 9764
rect 1946 9276 2254 9285
rect 1946 9274 1952 9276
rect 2008 9274 2032 9276
rect 2088 9274 2112 9276
rect 2168 9274 2192 9276
rect 2248 9274 2254 9276
rect 2008 9222 2010 9274
rect 2190 9222 2192 9274
rect 1946 9220 1952 9222
rect 2008 9220 2032 9222
rect 2088 9220 2112 9222
rect 2168 9220 2192 9222
rect 2248 9220 2254 9222
rect 1946 9211 2254 9220
rect 1306 8732 1614 8741
rect 1306 8730 1312 8732
rect 1368 8730 1392 8732
rect 1448 8730 1472 8732
rect 1528 8730 1552 8732
rect 1608 8730 1614 8732
rect 1368 8678 1370 8730
rect 1550 8678 1552 8730
rect 1306 8676 1312 8678
rect 1368 8676 1392 8678
rect 1448 8676 1472 8678
rect 1528 8676 1552 8678
rect 1608 8676 1614 8678
rect 1306 8667 1614 8676
rect 1946 8188 2254 8197
rect 1946 8186 1952 8188
rect 2008 8186 2032 8188
rect 2088 8186 2112 8188
rect 2168 8186 2192 8188
rect 2248 8186 2254 8188
rect 2008 8134 2010 8186
rect 2190 8134 2192 8186
rect 1946 8132 1952 8134
rect 2008 8132 2032 8134
rect 2088 8132 2112 8134
rect 2168 8132 2192 8134
rect 2248 8132 2254 8134
rect 1946 8123 2254 8132
rect 5092 8090 5120 11600
rect 5264 8356 5316 8362
rect 5264 8298 5316 8304
rect 5170 8256 5226 8265
rect 5170 8191 5226 8200
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 5080 8084 5132 8090
rect 5080 8026 5132 8032
rect 2780 7744 2832 7750
rect 2780 7686 2832 7692
rect 1306 7644 1614 7653
rect 1306 7642 1312 7644
rect 1368 7642 1392 7644
rect 1448 7642 1472 7644
rect 1528 7642 1552 7644
rect 1608 7642 1614 7644
rect 1368 7590 1370 7642
rect 1550 7590 1552 7642
rect 1306 7588 1312 7590
rect 1368 7588 1392 7590
rect 1448 7588 1472 7590
rect 1528 7588 1552 7590
rect 1608 7588 1614 7590
rect 1306 7579 1614 7588
rect 1946 7100 2254 7109
rect 1946 7098 1952 7100
rect 2008 7098 2032 7100
rect 2088 7098 2112 7100
rect 2168 7098 2192 7100
rect 2248 7098 2254 7100
rect 2008 7046 2010 7098
rect 2190 7046 2192 7098
rect 1946 7044 1952 7046
rect 2008 7044 2032 7046
rect 2088 7044 2112 7046
rect 2168 7044 2192 7046
rect 2248 7044 2254 7046
rect 1946 7035 2254 7044
rect 1306 6556 1614 6565
rect 1306 6554 1312 6556
rect 1368 6554 1392 6556
rect 1448 6554 1472 6556
rect 1528 6554 1552 6556
rect 1608 6554 1614 6556
rect 1368 6502 1370 6554
rect 1550 6502 1552 6554
rect 1306 6500 1312 6502
rect 1368 6500 1392 6502
rect 1448 6500 1472 6502
rect 1528 6500 1552 6502
rect 1608 6500 1614 6502
rect 1306 6491 1614 6500
rect 1946 6012 2254 6021
rect 1946 6010 1952 6012
rect 2008 6010 2032 6012
rect 2088 6010 2112 6012
rect 2168 6010 2192 6012
rect 2248 6010 2254 6012
rect 2008 5958 2010 6010
rect 2190 5958 2192 6010
rect 1946 5956 1952 5958
rect 2008 5956 2032 5958
rect 2088 5956 2112 5958
rect 2168 5956 2192 5958
rect 2248 5956 2254 5958
rect 1946 5947 2254 5956
rect 1306 5468 1614 5477
rect 1306 5466 1312 5468
rect 1368 5466 1392 5468
rect 1448 5466 1472 5468
rect 1528 5466 1552 5468
rect 1608 5466 1614 5468
rect 1368 5414 1370 5466
rect 1550 5414 1552 5466
rect 1306 5412 1312 5414
rect 1368 5412 1392 5414
rect 1448 5412 1472 5414
rect 1528 5412 1552 5414
rect 1608 5412 1614 5414
rect 1306 5403 1614 5412
rect 1946 4924 2254 4933
rect 1946 4922 1952 4924
rect 2008 4922 2032 4924
rect 2088 4922 2112 4924
rect 2168 4922 2192 4924
rect 2248 4922 2254 4924
rect 2008 4870 2010 4922
rect 2190 4870 2192 4922
rect 1946 4868 1952 4870
rect 2008 4868 2032 4870
rect 2088 4868 2112 4870
rect 2168 4868 2192 4870
rect 2248 4868 2254 4870
rect 1946 4859 2254 4868
rect 1306 4380 1614 4389
rect 1306 4378 1312 4380
rect 1368 4378 1392 4380
rect 1448 4378 1472 4380
rect 1528 4378 1552 4380
rect 1608 4378 1614 4380
rect 1368 4326 1370 4378
rect 1550 4326 1552 4378
rect 1306 4324 1312 4326
rect 1368 4324 1392 4326
rect 1448 4324 1472 4326
rect 1528 4324 1552 4326
rect 1608 4324 1614 4326
rect 1306 4315 1614 4324
rect 1946 3836 2254 3845
rect 1946 3834 1952 3836
rect 2008 3834 2032 3836
rect 2088 3834 2112 3836
rect 2168 3834 2192 3836
rect 2248 3834 2254 3836
rect 2008 3782 2010 3834
rect 2190 3782 2192 3834
rect 1946 3780 1952 3782
rect 2008 3780 2032 3782
rect 2088 3780 2112 3782
rect 2168 3780 2192 3782
rect 2248 3780 2254 3782
rect 1946 3771 2254 3780
rect 1306 3292 1614 3301
rect 1306 3290 1312 3292
rect 1368 3290 1392 3292
rect 1448 3290 1472 3292
rect 1528 3290 1552 3292
rect 1608 3290 1614 3292
rect 1368 3238 1370 3290
rect 1550 3238 1552 3290
rect 1306 3236 1312 3238
rect 1368 3236 1392 3238
rect 1448 3236 1472 3238
rect 1528 3236 1552 3238
rect 1608 3236 1614 3238
rect 1306 3227 1614 3236
rect 1946 2748 2254 2757
rect 1946 2746 1952 2748
rect 2008 2746 2032 2748
rect 2088 2746 2112 2748
rect 2168 2746 2192 2748
rect 2248 2746 2254 2748
rect 2008 2694 2010 2746
rect 2190 2694 2192 2746
rect 1946 2692 1952 2694
rect 2008 2692 2032 2694
rect 2088 2692 2112 2694
rect 2168 2692 2192 2694
rect 2248 2692 2254 2694
rect 1946 2683 2254 2692
rect 1306 2204 1614 2213
rect 1306 2202 1312 2204
rect 1368 2202 1392 2204
rect 1448 2202 1472 2204
rect 1528 2202 1552 2204
rect 1608 2202 1614 2204
rect 1368 2150 1370 2202
rect 1550 2150 1552 2202
rect 1306 2148 1312 2150
rect 1368 2148 1392 2150
rect 1448 2148 1472 2150
rect 1528 2148 1552 2150
rect 1608 2148 1614 2150
rect 1306 2139 1614 2148
rect 1946 1660 2254 1669
rect 1946 1658 1952 1660
rect 2008 1658 2032 1660
rect 2088 1658 2112 1660
rect 2168 1658 2192 1660
rect 2248 1658 2254 1660
rect 2008 1606 2010 1658
rect 2190 1606 2192 1658
rect 1946 1604 1952 1606
rect 2008 1604 2032 1606
rect 2088 1604 2112 1606
rect 2168 1604 2192 1606
rect 2248 1604 2254 1606
rect 1946 1595 2254 1604
rect 1306 1116 1614 1125
rect 1306 1114 1312 1116
rect 1368 1114 1392 1116
rect 1448 1114 1472 1116
rect 1528 1114 1552 1116
rect 1608 1114 1614 1116
rect 1368 1062 1370 1114
rect 1550 1062 1552 1114
rect 1306 1060 1312 1062
rect 1368 1060 1392 1062
rect 1448 1060 1472 1062
rect 1528 1060 1552 1062
rect 1608 1060 1614 1062
rect 1306 1051 1614 1060
rect 1946 572 2254 581
rect 1946 570 1952 572
rect 2008 570 2032 572
rect 2088 570 2112 572
rect 2168 570 2192 572
rect 2248 570 2254 572
rect 2008 518 2010 570
rect 2190 518 2192 570
rect 1946 516 1952 518
rect 2008 516 2032 518
rect 2088 516 2112 518
rect 2168 516 2192 518
rect 2248 516 2254 518
rect 1946 507 2254 516
rect 2792 400 2820 7686
rect 4264 7410 4292 8026
rect 4344 8016 4396 8022
rect 4344 7958 4396 7964
rect 4894 7984 4950 7993
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4160 7336 4212 7342
rect 4160 7278 4212 7284
rect 3056 7200 3108 7206
rect 3056 7142 3108 7148
rect 3068 400 3096 7142
rect 3884 6792 3936 6798
rect 3884 6734 3936 6740
rect 3332 6724 3384 6730
rect 3332 6666 3384 6672
rect 3344 400 3372 6666
rect 3608 6656 3660 6662
rect 3608 6598 3660 6604
rect 3620 400 3648 6598
rect 3896 400 3924 6734
rect 4172 6662 4200 7278
rect 4160 6656 4212 6662
rect 4160 6598 4212 6604
rect 4356 2774 4384 7958
rect 4894 7919 4950 7928
rect 4528 7540 4580 7546
rect 4528 7482 4580 7488
rect 4436 7200 4488 7206
rect 4436 7142 4488 7148
rect 4172 2746 4384 2774
rect 4172 400 4200 2746
rect 4448 400 4476 7142
rect 4540 7002 4568 7482
rect 4908 7410 4936 7919
rect 5184 7818 5212 8191
rect 5172 7812 5224 7818
rect 5172 7754 5224 7760
rect 4986 7440 5042 7449
rect 4896 7404 4948 7410
rect 4986 7375 4988 7384
rect 4896 7346 4948 7352
rect 5040 7375 5042 7384
rect 4988 7346 5040 7352
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4528 6996 4580 7002
rect 4528 6938 4580 6944
rect 4632 6798 4660 7210
rect 4620 6792 4672 6798
rect 4896 6792 4948 6798
rect 4620 6734 4672 6740
rect 4894 6760 4896 6769
rect 5080 6792 5132 6798
rect 4948 6760 4950 6769
rect 5080 6734 5132 6740
rect 4894 6695 4950 6704
rect 4804 6656 4856 6662
rect 4804 6598 4856 6604
rect 4816 2774 4844 6598
rect 5092 2774 5120 6734
rect 4724 2746 4844 2774
rect 5000 2746 5120 2774
rect 4724 400 4752 2746
rect 5000 400 5028 2746
rect 5276 400 5304 8298
rect 5368 7750 5396 11600
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5356 7744 5408 7750
rect 5356 7686 5408 7692
rect 5460 7342 5488 8230
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5552 7410 5580 8026
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5448 7336 5500 7342
rect 5448 7278 5500 7284
rect 5644 6866 5672 11600
rect 5920 7970 5948 11600
rect 6000 8288 6052 8294
rect 6000 8230 6052 8236
rect 6012 8022 6040 8230
rect 6196 8090 6224 11600
rect 6472 8634 6500 11600
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6184 8084 6236 8090
rect 6184 8026 6236 8032
rect 5736 7942 5948 7970
rect 6000 8016 6052 8022
rect 6000 7958 6052 7964
rect 6092 7948 6144 7954
rect 5736 7546 5764 7942
rect 6092 7890 6144 7896
rect 5816 7744 5868 7750
rect 5816 7686 5868 7692
rect 5724 7540 5776 7546
rect 5724 7482 5776 7488
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5644 6458 5672 6802
rect 5736 6798 5764 7346
rect 5724 6792 5776 6798
rect 5724 6734 5776 6740
rect 5632 6452 5684 6458
rect 5632 6394 5684 6400
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5552 400 5580 6054
rect 5828 400 5856 7686
rect 6000 7540 6052 7546
rect 6000 7482 6052 7488
rect 6012 7002 6040 7482
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6104 400 6132 7890
rect 6380 7478 6408 8230
rect 6472 8022 6500 8570
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 6460 8016 6512 8022
rect 6460 7958 6512 7964
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6368 7472 6420 7478
rect 6368 7414 6420 7420
rect 6276 7336 6328 7342
rect 6276 7278 6328 7284
rect 6288 7002 6316 7278
rect 6472 7274 6500 7686
rect 6564 7410 6592 8026
rect 6656 7954 6684 8298
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6748 7546 6776 11600
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 8022 6868 8366
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 6828 8016 6880 8022
rect 6828 7958 6880 7964
rect 6828 7880 6880 7886
rect 6826 7848 6828 7857
rect 6880 7848 6882 7857
rect 6826 7783 6882 7792
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 6552 7404 6604 7410
rect 6552 7346 6604 7352
rect 6460 7268 6512 7274
rect 6460 7210 6512 7216
rect 6276 6996 6328 7002
rect 6276 6938 6328 6944
rect 6276 6792 6328 6798
rect 6276 6734 6328 6740
rect 6288 6225 6316 6734
rect 6828 6724 6880 6730
rect 6828 6666 6880 6672
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6274 6216 6330 6225
rect 6274 6151 6330 6160
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6380 400 6408 6122
rect 6656 400 6684 6598
rect 6840 6118 6868 6666
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6932 400 6960 8298
rect 7024 6866 7052 11600
rect 7300 8090 7328 11600
rect 7576 8634 7604 11600
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7378 8528 7434 8537
rect 7378 8463 7434 8472
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7012 6860 7064 6866
rect 7012 6802 7064 6808
rect 7104 6792 7156 6798
rect 7104 6734 7156 6740
rect 7116 6361 7144 6734
rect 7102 6352 7158 6361
rect 7102 6287 7158 6296
rect 7208 400 7236 7686
rect 7392 7546 7420 8463
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7484 7410 7512 8026
rect 7576 8022 7604 8570
rect 7564 8016 7616 8022
rect 7564 7958 7616 7964
rect 7472 7404 7524 7410
rect 7472 7346 7524 7352
rect 7380 7336 7432 7342
rect 7380 7278 7432 7284
rect 7392 6186 7420 7278
rect 7852 6866 7880 11600
rect 8024 8424 8076 8430
rect 8024 8366 8076 8372
rect 7840 6860 7892 6866
rect 7840 6802 7892 6808
rect 7748 6724 7800 6730
rect 7748 6666 7800 6672
rect 7380 6180 7432 6186
rect 7380 6122 7432 6128
rect 7472 6180 7524 6186
rect 7472 6122 7524 6128
rect 7484 400 7512 6122
rect 7760 6118 7788 6666
rect 7852 6458 7880 6802
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7748 6112 7800 6118
rect 7748 6054 7800 6060
rect 7760 400 7788 6054
rect 8036 400 8064 8366
rect 8128 8090 8156 11600
rect 8404 8634 8432 11600
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8116 8084 8168 8090
rect 8116 8026 8168 8032
rect 8404 8022 8432 8570
rect 8576 8356 8628 8362
rect 8576 8298 8628 8304
rect 8392 8016 8444 8022
rect 8392 7958 8444 7964
rect 8588 7954 8616 8298
rect 8576 7948 8628 7954
rect 8576 7890 8628 7896
rect 8208 7744 8260 7750
rect 8208 7686 8260 7692
rect 8220 7342 8248 7686
rect 8680 7410 8708 11600
rect 8760 9512 8812 9518
rect 8760 9454 8812 9460
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8208 7336 8260 7342
rect 8114 7304 8170 7313
rect 8208 7278 8260 7284
rect 8114 7239 8170 7248
rect 8128 7206 8156 7239
rect 8116 7200 8168 7206
rect 8116 7142 8168 7148
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8312 400 8340 7142
rect 8680 6458 8708 7346
rect 8772 6866 8800 9454
rect 8760 6860 8812 6866
rect 8760 6802 8812 6808
rect 8852 6792 8904 6798
rect 8852 6734 8904 6740
rect 8864 6458 8892 6734
rect 8956 6662 8984 11600
rect 9128 11008 9180 11014
rect 9128 10950 9180 10956
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 9048 7206 9076 8502
rect 9140 7546 9168 10950
rect 9232 8634 9260 11600
rect 9508 11014 9536 11600
rect 9496 11008 9548 11014
rect 9496 10950 9548 10956
rect 9306 10908 9614 10917
rect 9306 10906 9312 10908
rect 9368 10906 9392 10908
rect 9448 10906 9472 10908
rect 9528 10906 9552 10908
rect 9608 10906 9614 10908
rect 9368 10854 9370 10906
rect 9550 10854 9552 10906
rect 9306 10852 9312 10854
rect 9368 10852 9392 10854
rect 9448 10852 9472 10854
rect 9528 10852 9552 10854
rect 9608 10852 9614 10854
rect 9306 10843 9614 10852
rect 9306 9820 9614 9829
rect 9306 9818 9312 9820
rect 9368 9818 9392 9820
rect 9448 9818 9472 9820
rect 9528 9818 9552 9820
rect 9608 9818 9614 9820
rect 9368 9766 9370 9818
rect 9550 9766 9552 9818
rect 9306 9764 9312 9766
rect 9368 9764 9392 9766
rect 9448 9764 9472 9766
rect 9528 9764 9552 9766
rect 9608 9764 9614 9766
rect 9306 9755 9614 9764
rect 9784 8809 9812 11600
rect 10060 11558 10088 11600
rect 10048 11552 10100 11558
rect 10048 11494 10100 11500
rect 9946 11452 10254 11461
rect 9946 11450 9952 11452
rect 10008 11450 10032 11452
rect 10088 11450 10112 11452
rect 10168 11450 10192 11452
rect 10248 11450 10254 11452
rect 10008 11398 10010 11450
rect 10190 11398 10192 11450
rect 9946 11396 9952 11398
rect 10008 11396 10032 11398
rect 10088 11396 10112 11398
rect 10168 11396 10192 11398
rect 10248 11396 10254 11398
rect 9946 11387 10254 11396
rect 9946 10364 10254 10373
rect 9946 10362 9952 10364
rect 10008 10362 10032 10364
rect 10088 10362 10112 10364
rect 10168 10362 10192 10364
rect 10248 10362 10254 10364
rect 10008 10310 10010 10362
rect 10190 10310 10192 10362
rect 9946 10308 9952 10310
rect 10008 10308 10032 10310
rect 10088 10308 10112 10310
rect 10168 10308 10192 10310
rect 10248 10308 10254 10310
rect 9946 10299 10254 10308
rect 9946 9276 10254 9285
rect 9946 9274 9952 9276
rect 10008 9274 10032 9276
rect 10088 9274 10112 9276
rect 10168 9274 10192 9276
rect 10248 9274 10254 9276
rect 10008 9222 10010 9274
rect 10190 9222 10192 9274
rect 9946 9220 9952 9222
rect 10008 9220 10032 9222
rect 10088 9220 10112 9222
rect 10168 9220 10192 9222
rect 10248 9220 10254 9222
rect 9946 9211 10254 9220
rect 10140 9104 10192 9110
rect 10140 9046 10192 9052
rect 9770 8800 9826 8809
rect 9306 8732 9614 8741
rect 9770 8735 9826 8744
rect 9306 8730 9312 8732
rect 9368 8730 9392 8732
rect 9448 8730 9472 8732
rect 9528 8730 9552 8732
rect 9608 8730 9614 8732
rect 9368 8678 9370 8730
rect 9550 8678 9552 8730
rect 9306 8676 9312 8678
rect 9368 8676 9392 8678
rect 9448 8676 9472 8678
rect 9528 8676 9552 8678
rect 9608 8676 9614 8678
rect 9306 8667 9614 8676
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9232 8022 9260 8570
rect 9496 8424 9548 8430
rect 9680 8424 9732 8430
rect 9496 8366 9548 8372
rect 9600 8372 9680 8378
rect 9600 8366 9732 8372
rect 9508 8022 9536 8366
rect 9600 8350 9720 8366
rect 9220 8016 9272 8022
rect 9220 7958 9272 7964
rect 9496 8016 9548 8022
rect 9496 7958 9548 7964
rect 9600 7834 9628 8350
rect 9678 8120 9734 8129
rect 9678 8055 9734 8064
rect 9692 7834 9720 8055
rect 9600 7806 9720 7834
rect 9876 7732 9904 8570
rect 10152 8498 10180 9046
rect 10140 8492 10192 8498
rect 10140 8434 10192 8440
rect 9946 8188 10254 8197
rect 9946 8186 9952 8188
rect 10008 8186 10032 8188
rect 10088 8186 10112 8188
rect 10168 8186 10192 8188
rect 10248 8186 10254 8188
rect 10008 8134 10010 8186
rect 10190 8134 10192 8186
rect 9946 8132 9952 8134
rect 10008 8132 10032 8134
rect 10088 8132 10112 8134
rect 10168 8132 10192 8134
rect 10248 8132 10254 8134
rect 9946 8123 10254 8132
rect 10336 8090 10364 11600
rect 10416 11552 10468 11558
rect 10416 11494 10468 11500
rect 10428 8412 10456 11494
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10520 8566 10548 8774
rect 10612 8634 10640 11600
rect 10888 9330 10916 11600
rect 11164 9738 11192 11600
rect 10796 9302 10916 9330
rect 10980 9710 11192 9738
rect 10690 9072 10746 9081
rect 10690 9007 10746 9016
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10508 8560 10560 8566
rect 10560 8508 10640 8514
rect 10508 8502 10640 8508
rect 10520 8486 10640 8502
rect 10704 8498 10732 9007
rect 10428 8384 10548 8412
rect 10416 8288 10468 8294
rect 10416 8230 10468 8236
rect 10324 8084 10376 8090
rect 10324 8026 10376 8032
rect 10428 7970 10456 8230
rect 9968 7942 10456 7970
rect 9968 7886 9996 7942
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 10140 7880 10192 7886
rect 10140 7822 10192 7828
rect 10324 7880 10376 7886
rect 10324 7822 10376 7828
rect 9876 7704 10088 7732
rect 9306 7644 9614 7653
rect 9306 7642 9312 7644
rect 9368 7642 9392 7644
rect 9448 7642 9472 7644
rect 9528 7642 9552 7644
rect 9608 7642 9614 7644
rect 9368 7590 9370 7642
rect 9550 7590 9552 7642
rect 9306 7588 9312 7590
rect 9368 7588 9392 7590
rect 9448 7588 9472 7590
rect 9528 7588 9552 7590
rect 9608 7588 9614 7590
rect 9306 7579 9614 7588
rect 9128 7540 9180 7546
rect 9128 7482 9180 7488
rect 10060 7478 10088 7704
rect 10152 7585 10180 7822
rect 10138 7576 10194 7585
rect 10138 7511 10194 7520
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 10140 7336 10192 7342
rect 10140 7278 10192 7284
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8668 6452 8720 6458
rect 8668 6394 8720 6400
rect 8852 6452 8904 6458
rect 8852 6394 8904 6400
rect 8944 6248 8996 6254
rect 8944 6190 8996 6196
rect 8956 5778 8984 6190
rect 8944 5772 8996 5778
rect 8944 5714 8996 5720
rect 8576 5636 8628 5642
rect 8576 5578 8628 5584
rect 8588 400 8616 5578
rect 9048 5250 9076 7142
rect 9324 6934 9352 7278
rect 10152 7206 10180 7278
rect 10140 7200 10192 7206
rect 10140 7142 10192 7148
rect 9946 7100 10254 7109
rect 9946 7098 9952 7100
rect 10008 7098 10032 7100
rect 10088 7098 10112 7100
rect 10168 7098 10192 7100
rect 10248 7098 10254 7100
rect 10008 7046 10010 7098
rect 10190 7046 10192 7098
rect 9946 7044 9952 7046
rect 10008 7044 10032 7046
rect 10088 7044 10112 7046
rect 10168 7044 10192 7046
rect 10248 7044 10254 7046
rect 9946 7035 10254 7044
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9494 6896 9550 6905
rect 9494 6831 9496 6840
rect 9548 6831 9550 6840
rect 9956 6860 10008 6866
rect 9496 6802 9548 6808
rect 9956 6802 10008 6808
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 5574 9168 6734
rect 9864 6656 9916 6662
rect 9864 6598 9916 6604
rect 9306 6556 9614 6565
rect 9306 6554 9312 6556
rect 9368 6554 9392 6556
rect 9448 6554 9472 6556
rect 9528 6554 9552 6556
rect 9608 6554 9614 6556
rect 9368 6502 9370 6554
rect 9550 6502 9552 6554
rect 9306 6500 9312 6502
rect 9368 6500 9392 6502
rect 9448 6500 9472 6502
rect 9528 6500 9552 6502
rect 9608 6500 9614 6502
rect 9306 6491 9614 6500
rect 9770 6488 9826 6497
rect 9770 6423 9826 6432
rect 9784 6390 9812 6423
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9588 6180 9640 6186
rect 9588 6122 9640 6128
rect 9220 6112 9272 6118
rect 9220 6054 9272 6060
rect 9128 5568 9180 5574
rect 9128 5510 9180 5516
rect 8864 5222 9076 5250
rect 8864 400 8892 5222
rect 9140 400 9168 5510
rect 9232 898 9260 6054
rect 9600 5642 9628 6122
rect 9784 5914 9812 6326
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 9876 5846 9904 6598
rect 9968 6118 9996 6802
rect 10140 6792 10192 6798
rect 10140 6734 10192 6740
rect 10152 6633 10180 6734
rect 10138 6624 10194 6633
rect 10138 6559 10194 6568
rect 9956 6112 10008 6118
rect 9956 6054 10008 6060
rect 9946 6012 10254 6021
rect 9946 6010 9952 6012
rect 10008 6010 10032 6012
rect 10088 6010 10112 6012
rect 10168 6010 10192 6012
rect 10248 6010 10254 6012
rect 10008 5958 10010 6010
rect 10190 5958 10192 6010
rect 9946 5956 9952 5958
rect 10008 5956 10032 5958
rect 10088 5956 10112 5958
rect 10168 5956 10192 5958
rect 10248 5956 10254 5958
rect 9946 5947 10254 5956
rect 9864 5840 9916 5846
rect 9864 5782 9916 5788
rect 9588 5636 9640 5642
rect 9588 5578 9640 5584
rect 9306 5468 9614 5477
rect 9306 5466 9312 5468
rect 9368 5466 9392 5468
rect 9448 5466 9472 5468
rect 9528 5466 9552 5468
rect 9608 5466 9614 5468
rect 9368 5414 9370 5466
rect 9550 5414 9552 5466
rect 9306 5412 9312 5414
rect 9368 5412 9392 5414
rect 9448 5412 9472 5414
rect 9528 5412 9552 5414
rect 9608 5412 9614 5414
rect 9306 5403 9614 5412
rect 9306 4380 9614 4389
rect 9306 4378 9312 4380
rect 9368 4378 9392 4380
rect 9448 4378 9472 4380
rect 9528 4378 9552 4380
rect 9608 4378 9614 4380
rect 9368 4326 9370 4378
rect 9550 4326 9552 4378
rect 9306 4324 9312 4326
rect 9368 4324 9392 4326
rect 9448 4324 9472 4326
rect 9528 4324 9552 4326
rect 9608 4324 9614 4326
rect 9306 4315 9614 4324
rect 9864 4208 9916 4214
rect 9864 4150 9916 4156
rect 9678 4040 9734 4049
rect 9678 3975 9734 3984
rect 9306 3292 9614 3301
rect 9306 3290 9312 3292
rect 9368 3290 9392 3292
rect 9448 3290 9472 3292
rect 9528 3290 9552 3292
rect 9608 3290 9614 3292
rect 9368 3238 9370 3290
rect 9550 3238 9552 3290
rect 9306 3236 9312 3238
rect 9368 3236 9392 3238
rect 9448 3236 9472 3238
rect 9528 3236 9552 3238
rect 9608 3236 9614 3238
rect 9306 3227 9614 3236
rect 9306 2204 9614 2213
rect 9306 2202 9312 2204
rect 9368 2202 9392 2204
rect 9448 2202 9472 2204
rect 9528 2202 9552 2204
rect 9608 2202 9614 2204
rect 9368 2150 9370 2202
rect 9550 2150 9552 2202
rect 9306 2148 9312 2150
rect 9368 2148 9392 2150
rect 9448 2148 9472 2150
rect 9528 2148 9552 2150
rect 9608 2148 9614 2150
rect 9306 2139 9614 2148
rect 9306 1116 9614 1125
rect 9306 1114 9312 1116
rect 9368 1114 9392 1116
rect 9448 1114 9472 1116
rect 9528 1114 9552 1116
rect 9608 1114 9614 1116
rect 9368 1062 9370 1114
rect 9550 1062 9552 1114
rect 9306 1060 9312 1062
rect 9368 1060 9392 1062
rect 9448 1060 9472 1062
rect 9528 1060 9552 1062
rect 9608 1060 9614 1062
rect 9306 1051 9614 1060
rect 9232 870 9444 898
rect 9416 400 9444 870
rect 9692 400 9720 3975
rect 9876 456 9904 4150
rect 9946 3836 10254 3845
rect 9946 3834 9952 3836
rect 10008 3834 10032 3836
rect 10088 3834 10112 3836
rect 10168 3834 10192 3836
rect 10248 3834 10254 3836
rect 10008 3782 10010 3834
rect 10190 3782 10192 3834
rect 9946 3780 9952 3782
rect 10008 3780 10032 3782
rect 10088 3780 10112 3782
rect 10168 3780 10192 3782
rect 10248 3780 10254 3782
rect 9946 3771 10254 3780
rect 9946 2748 10254 2757
rect 9946 2746 9952 2748
rect 10008 2746 10032 2748
rect 10088 2746 10112 2748
rect 10168 2746 10192 2748
rect 10248 2746 10254 2748
rect 10008 2694 10010 2746
rect 10190 2694 10192 2746
rect 9946 2692 9952 2694
rect 10008 2692 10032 2694
rect 10088 2692 10112 2694
rect 10168 2692 10192 2694
rect 10248 2692 10254 2694
rect 9946 2683 10254 2692
rect 9946 1660 10254 1669
rect 9946 1658 9952 1660
rect 10008 1658 10032 1660
rect 10088 1658 10112 1660
rect 10168 1658 10192 1660
rect 10248 1658 10254 1660
rect 10008 1606 10010 1658
rect 10190 1606 10192 1658
rect 9946 1604 9952 1606
rect 10008 1604 10032 1606
rect 10088 1604 10112 1606
rect 10168 1604 10192 1606
rect 10248 1604 10254 1606
rect 9946 1595 10254 1604
rect 9946 572 10254 581
rect 9946 570 9952 572
rect 10008 570 10032 572
rect 10088 570 10112 572
rect 10168 570 10192 572
rect 10248 570 10254 572
rect 10008 518 10010 570
rect 10190 518 10192 570
rect 9946 516 9952 518
rect 10008 516 10032 518
rect 10088 516 10112 518
rect 10168 516 10192 518
rect 10248 516 10254 518
rect 9946 507 10254 516
rect 10336 456 10364 7822
rect 10414 7032 10470 7041
rect 10414 6967 10470 6976
rect 10428 6730 10456 6967
rect 10416 6724 10468 6730
rect 10416 6666 10468 6672
rect 10428 5914 10456 6666
rect 10520 6662 10548 8384
rect 10508 6656 10560 6662
rect 10508 6598 10560 6604
rect 10508 6384 10560 6390
rect 10508 6326 10560 6332
rect 10520 5914 10548 6326
rect 10416 5908 10468 5914
rect 10416 5850 10468 5856
rect 10508 5908 10560 5914
rect 10508 5850 10560 5856
rect 10612 2774 10640 8486
rect 10692 8492 10744 8498
rect 10692 8434 10744 8440
rect 10690 8392 10746 8401
rect 10690 8327 10692 8336
rect 10744 8327 10746 8336
rect 10692 8298 10744 8304
rect 10690 8256 10746 8265
rect 10690 8191 10746 8200
rect 10704 7585 10732 8191
rect 10690 7576 10746 7585
rect 10690 7511 10746 7520
rect 10692 7404 10744 7410
rect 10692 7346 10744 7352
rect 10704 7206 10732 7346
rect 10692 7200 10744 7206
rect 10692 7142 10744 7148
rect 10796 6390 10824 9302
rect 10874 9208 10930 9217
rect 10874 9143 10930 9152
rect 10888 9042 10916 9143
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10876 8900 10928 8906
rect 10876 8842 10928 8848
rect 10784 6384 10836 6390
rect 10784 6326 10836 6332
rect 10784 6248 10836 6254
rect 10784 6190 10836 6196
rect 9876 428 9996 456
rect 9968 400 9996 428
rect 10244 428 10364 456
rect 10520 2746 10640 2774
rect 10244 400 10272 428
rect 10520 400 10548 2746
rect 10796 400 10824 6190
rect 10888 4214 10916 8842
rect 10980 8090 11008 9710
rect 11440 9674 11468 11600
rect 11440 9646 11560 9674
rect 11060 9580 11112 9586
rect 11060 9522 11112 9528
rect 11072 8498 11100 9522
rect 11336 8560 11388 8566
rect 11336 8502 11388 8508
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 10968 8084 11020 8090
rect 10968 8026 11020 8032
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 10980 7342 11008 8026
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 11072 7342 11100 7686
rect 11152 7540 11204 7546
rect 11152 7482 11204 7488
rect 10968 7336 11020 7342
rect 10968 7278 11020 7284
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 11072 400 11100 7278
rect 11164 6866 11192 7482
rect 11256 6934 11284 8026
rect 11348 7886 11376 8502
rect 11428 8424 11480 8430
rect 11428 8366 11480 8372
rect 11336 7880 11388 7886
rect 11336 7822 11388 7828
rect 11334 7576 11390 7585
rect 11334 7511 11390 7520
rect 11244 6928 11296 6934
rect 11244 6870 11296 6876
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 11348 6458 11376 7511
rect 11336 6452 11388 6458
rect 11336 6394 11388 6400
rect 11336 5840 11388 5846
rect 11336 5782 11388 5788
rect 11348 400 11376 5782
rect 11440 2774 11468 8366
rect 11532 8072 11560 9646
rect 11612 8968 11664 8974
rect 11612 8910 11664 8916
rect 11624 8498 11652 8910
rect 11612 8492 11664 8498
rect 11612 8434 11664 8440
rect 11532 8044 11652 8072
rect 11518 7984 11574 7993
rect 11518 7919 11574 7928
rect 11532 6390 11560 7919
rect 11624 7041 11652 8044
rect 11610 7032 11666 7041
rect 11610 6967 11666 6976
rect 11716 6798 11744 11600
rect 11992 9042 12020 11600
rect 12268 9178 12296 11600
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12072 9104 12124 9110
rect 12072 9046 12124 9052
rect 11980 9036 12032 9042
rect 11980 8978 12032 8984
rect 11980 8900 12032 8906
rect 11980 8842 12032 8848
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8430 11928 8774
rect 11888 8424 11940 8430
rect 11888 8366 11940 8372
rect 11888 7880 11940 7886
rect 11888 7822 11940 7828
rect 11796 7744 11848 7750
rect 11796 7686 11848 7692
rect 11704 6792 11756 6798
rect 11704 6734 11756 6740
rect 11520 6384 11572 6390
rect 11520 6326 11572 6332
rect 11808 6202 11836 7686
rect 11900 7313 11928 7822
rect 11886 7304 11942 7313
rect 11886 7239 11942 7248
rect 11886 7032 11942 7041
rect 11886 6967 11942 6976
rect 11532 6174 11836 6202
rect 11532 6118 11560 6174
rect 11520 6112 11572 6118
rect 11520 6054 11572 6060
rect 11900 5778 11928 6967
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11992 2774 12020 8842
rect 12084 8838 12112 9046
rect 12440 9036 12492 9042
rect 12440 8978 12492 8984
rect 12072 8832 12124 8838
rect 12072 8774 12124 8780
rect 12084 5846 12112 8774
rect 12164 8492 12216 8498
rect 12164 8434 12216 8440
rect 12072 5840 12124 5846
rect 12072 5782 12124 5788
rect 11440 2746 11652 2774
rect 11624 400 11652 2746
rect 11900 2746 12020 2774
rect 11900 400 11928 2746
rect 12176 400 12204 8434
rect 12254 8120 12310 8129
rect 12254 8055 12310 8064
rect 12268 7313 12296 8055
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12254 7304 12310 7313
rect 12254 7239 12310 7248
rect 12360 7002 12388 7482
rect 12452 7041 12480 8978
rect 12544 8566 12572 11600
rect 12716 9376 12768 9382
rect 12716 9318 12768 9324
rect 12622 8664 12678 8673
rect 12622 8599 12678 8608
rect 12532 8560 12584 8566
rect 12532 8502 12584 8508
rect 12636 8430 12664 8599
rect 12624 8424 12676 8430
rect 12624 8366 12676 8372
rect 12438 7032 12494 7041
rect 12348 6996 12400 7002
rect 12438 6967 12494 6976
rect 12348 6938 12400 6944
rect 12438 1320 12494 1329
rect 12438 1255 12494 1264
rect 12452 400 12480 1255
rect 12728 400 12756 9318
rect 12820 8974 12848 11600
rect 12992 9648 13044 9654
rect 12992 9590 13044 9596
rect 13004 9110 13032 9590
rect 12992 9104 13044 9110
rect 12992 9046 13044 9052
rect 12808 8968 12860 8974
rect 12808 8910 12860 8916
rect 12900 7676 12952 7682
rect 12900 7618 12952 7624
rect 12912 6934 12940 7618
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 13096 6662 13124 11600
rect 13268 9444 13320 9450
rect 13268 9386 13320 9392
rect 13174 8392 13230 8401
rect 13280 8362 13308 9386
rect 13174 8327 13230 8336
rect 13268 8356 13320 8362
rect 13188 7290 13216 8327
rect 13268 8298 13320 8304
rect 13372 7682 13400 11600
rect 13452 10124 13504 10130
rect 13452 10066 13504 10072
rect 13464 9586 13492 10066
rect 13648 9654 13676 11600
rect 13636 9648 13688 9654
rect 13636 9590 13688 9596
rect 13452 9580 13504 9586
rect 13452 9522 13504 9528
rect 13820 9580 13872 9586
rect 13820 9522 13872 9528
rect 13636 9376 13688 9382
rect 13636 9318 13688 9324
rect 13648 8906 13676 9318
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13832 8498 13860 9522
rect 13924 8634 13952 11600
rect 14096 9920 14148 9926
rect 14096 9862 14148 9868
rect 14002 9616 14058 9625
rect 14002 9551 14058 9560
rect 14016 9081 14044 9551
rect 14108 9518 14136 9862
rect 14096 9512 14148 9518
rect 14094 9480 14096 9489
rect 14148 9480 14150 9489
rect 14094 9415 14150 9424
rect 14002 9072 14058 9081
rect 14002 9007 14058 9016
rect 14200 8838 14228 11600
rect 14476 10282 14504 11600
rect 14384 10254 14504 10282
rect 14752 10266 14780 11600
rect 14740 10260 14792 10266
rect 14384 9722 14412 10254
rect 14740 10202 14792 10208
rect 14464 10192 14516 10198
rect 14464 10134 14516 10140
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14280 9580 14332 9586
rect 14280 9522 14332 9528
rect 14292 9042 14320 9522
rect 14370 9208 14426 9217
rect 14370 9143 14426 9152
rect 14384 9110 14412 9143
rect 14476 9110 14504 10134
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14372 9104 14424 9110
rect 14372 9046 14424 9052
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 14660 9042 14688 9862
rect 14752 9586 14780 10202
rect 15028 10198 15056 11600
rect 15016 10192 15068 10198
rect 15016 10134 15068 10140
rect 14740 9580 14792 9586
rect 14740 9522 14792 9528
rect 15200 9580 15252 9586
rect 15200 9522 15252 9528
rect 14740 9444 14792 9450
rect 14740 9386 14792 9392
rect 14752 9081 14780 9386
rect 14738 9072 14794 9081
rect 14280 9036 14332 9042
rect 14280 8978 14332 8984
rect 14648 9036 14700 9042
rect 14738 9007 14794 9016
rect 14922 9072 14978 9081
rect 15212 9042 15240 9522
rect 14922 9007 14978 9016
rect 15200 9036 15252 9042
rect 14648 8978 14700 8984
rect 14660 8945 14688 8978
rect 14646 8936 14702 8945
rect 14646 8871 14702 8880
rect 14188 8832 14240 8838
rect 14188 8774 14240 8780
rect 13912 8628 13964 8634
rect 13912 8570 13964 8576
rect 14936 8566 14964 9007
rect 15200 8978 15252 8984
rect 15106 8664 15162 8673
rect 15304 8634 15332 11600
rect 15580 9654 15608 11600
rect 15660 10056 15712 10062
rect 15660 9998 15712 10004
rect 15568 9648 15620 9654
rect 15568 9590 15620 9596
rect 15476 9444 15528 9450
rect 15476 9386 15528 9392
rect 15384 9376 15436 9382
rect 15384 9318 15436 9324
rect 15106 8599 15162 8608
rect 15292 8628 15344 8634
rect 14924 8560 14976 8566
rect 14924 8502 14976 8508
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 14372 8492 14424 8498
rect 15016 8492 15068 8498
rect 14424 8452 14504 8480
rect 14372 8434 14424 8440
rect 14476 8412 14504 8452
rect 15016 8434 15068 8440
rect 14740 8424 14792 8430
rect 13450 8392 13506 8401
rect 14476 8384 14740 8412
rect 14740 8366 14792 8372
rect 13450 8327 13452 8336
rect 13504 8327 13506 8336
rect 14004 8356 14056 8362
rect 13452 8298 13504 8304
rect 14004 8298 14056 8304
rect 14016 8090 14044 8298
rect 14752 8265 14780 8366
rect 14554 8256 14610 8265
rect 14554 8191 14610 8200
rect 14738 8256 14794 8265
rect 14738 8191 14794 8200
rect 14568 8090 14596 8191
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14556 8084 14608 8090
rect 14556 8026 14608 8032
rect 14740 7880 14792 7886
rect 14186 7848 14242 7857
rect 13544 7812 13596 7818
rect 15028 7857 15056 8434
rect 15120 7886 15148 8599
rect 15292 8570 15344 8576
rect 15396 8430 15424 9318
rect 15488 9042 15516 9386
rect 15580 9110 15608 9590
rect 15672 9353 15700 9998
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15658 9344 15714 9353
rect 15658 9279 15714 9288
rect 15660 9172 15712 9178
rect 15660 9114 15712 9120
rect 15568 9104 15620 9110
rect 15568 9046 15620 9052
rect 15476 9036 15528 9042
rect 15476 8978 15528 8984
rect 15672 8616 15700 9114
rect 15580 8588 15700 8616
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15396 8265 15424 8366
rect 15382 8256 15438 8265
rect 15382 8191 15438 8200
rect 15108 7880 15160 7886
rect 14740 7822 14792 7828
rect 15014 7848 15070 7857
rect 14186 7783 14242 7792
rect 13544 7754 13596 7760
rect 13360 7676 13412 7682
rect 13360 7618 13412 7624
rect 13452 7676 13504 7682
rect 13452 7618 13504 7624
rect 13464 7478 13492 7618
rect 13452 7472 13504 7478
rect 13452 7414 13504 7420
rect 13556 7410 13584 7754
rect 14200 7562 14228 7783
rect 14602 7608 14654 7614
rect 14200 7534 14274 7562
rect 14602 7550 14654 7556
rect 14752 7562 14780 7822
rect 15108 7822 15160 7828
rect 15014 7783 15070 7792
rect 15290 7712 15346 7721
rect 15290 7647 15346 7656
rect 15304 7562 15332 7647
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 14246 7344 14274 7534
rect 14416 7372 14472 7381
rect 14614 7344 14642 7550
rect 14752 7534 14826 7562
rect 14798 7344 14826 7534
rect 15154 7540 15206 7546
rect 15304 7534 15378 7562
rect 15580 7546 15608 8588
rect 15658 8528 15714 8537
rect 15658 8463 15714 8472
rect 15672 7562 15700 8463
rect 15764 8412 15792 9590
rect 15856 9586 15884 11600
rect 16132 9654 16160 11600
rect 16212 9920 16264 9926
rect 16212 9862 16264 9868
rect 16304 9920 16356 9926
rect 16304 9862 16356 9868
rect 16120 9648 16172 9654
rect 16120 9590 16172 9596
rect 15844 9580 15896 9586
rect 15844 9522 15896 9528
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 15844 9376 15896 9382
rect 16040 9353 16068 9454
rect 15844 9318 15896 9324
rect 16026 9344 16082 9353
rect 15856 8945 15884 9318
rect 16026 9279 16082 9288
rect 15936 8968 15988 8974
rect 15842 8936 15898 8945
rect 15936 8910 15988 8916
rect 15842 8871 15898 8880
rect 15948 8537 15976 8910
rect 16028 8832 16080 8838
rect 16028 8774 16080 8780
rect 15934 8528 15990 8537
rect 15934 8463 15990 8472
rect 15764 8384 15976 8412
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15856 7562 15884 8230
rect 15948 8106 15976 8384
rect 16040 8362 16068 8774
rect 16132 8498 16160 9590
rect 16224 9518 16252 9862
rect 16212 9512 16264 9518
rect 16210 9480 16212 9489
rect 16264 9480 16266 9489
rect 16210 9415 16266 9424
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 16224 8498 16252 8774
rect 16316 8514 16344 9862
rect 16408 9178 16436 11600
rect 16684 10266 16712 11600
rect 16672 10260 16724 10266
rect 16672 10202 16724 10208
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16592 9586 16620 9930
rect 16684 9722 16712 10202
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16580 9580 16632 9586
rect 16580 9522 16632 9528
rect 16486 9208 16542 9217
rect 16396 9172 16448 9178
rect 16486 9143 16488 9152
rect 16396 9114 16448 9120
rect 16540 9143 16542 9152
rect 16488 9114 16540 9120
rect 16408 8634 16436 9114
rect 16592 8673 16620 9522
rect 16868 9518 16896 9862
rect 16672 9512 16724 9518
rect 16672 9454 16724 9460
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16684 8809 16712 9454
rect 16960 9450 16988 11600
rect 17132 11008 17184 11014
rect 17132 10950 17184 10956
rect 17040 9920 17092 9926
rect 17040 9862 17092 9868
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16670 8800 16726 8809
rect 16670 8735 16726 8744
rect 16578 8664 16634 8673
rect 16396 8628 16448 8634
rect 16776 8650 16804 8978
rect 16578 8599 16634 8608
rect 16684 8622 16804 8650
rect 16396 8570 16448 8576
rect 16684 8514 16712 8622
rect 16960 8566 16988 9386
rect 17052 8945 17080 9862
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 17144 8838 17172 10950
rect 17236 10266 17264 11600
rect 17512 11014 17540 11600
rect 17500 11008 17552 11014
rect 17500 10950 17552 10956
rect 17306 10908 17614 10917
rect 17306 10906 17312 10908
rect 17368 10906 17392 10908
rect 17448 10906 17472 10908
rect 17528 10906 17552 10908
rect 17608 10906 17614 10908
rect 17368 10854 17370 10906
rect 17550 10854 17552 10906
rect 17306 10852 17312 10854
rect 17368 10852 17392 10854
rect 17448 10852 17472 10854
rect 17528 10852 17552 10854
rect 17608 10852 17614 10854
rect 17306 10843 17614 10852
rect 17788 10282 17816 11600
rect 18064 11558 18092 11600
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18340 11506 18368 11600
rect 18340 11478 18552 11506
rect 17946 11452 18254 11461
rect 17946 11450 17952 11452
rect 18008 11450 18032 11452
rect 18088 11450 18112 11452
rect 18168 11450 18192 11452
rect 18248 11450 18254 11452
rect 18008 11398 18010 11450
rect 18190 11398 18192 11450
rect 17946 11396 17952 11398
rect 18008 11396 18032 11398
rect 18088 11396 18112 11398
rect 18168 11396 18192 11398
rect 18248 11396 18254 11398
rect 17946 11387 18254 11396
rect 17946 10364 18254 10373
rect 17946 10362 17952 10364
rect 18008 10362 18032 10364
rect 18088 10362 18112 10364
rect 18168 10362 18192 10364
rect 18248 10362 18254 10364
rect 18008 10310 18010 10362
rect 18190 10310 18192 10362
rect 17946 10308 17952 10310
rect 18008 10308 18032 10310
rect 18088 10308 18112 10310
rect 18168 10308 18192 10310
rect 18248 10308 18254 10310
rect 17946 10299 18254 10308
rect 17224 10260 17276 10266
rect 17224 10202 17276 10208
rect 17696 10254 17816 10282
rect 18052 10260 18104 10266
rect 17236 9722 17264 10202
rect 17306 9820 17614 9829
rect 17306 9818 17312 9820
rect 17368 9818 17392 9820
rect 17448 9818 17472 9820
rect 17528 9818 17552 9820
rect 17608 9818 17614 9820
rect 17368 9766 17370 9818
rect 17550 9766 17552 9818
rect 17306 9764 17312 9766
rect 17368 9764 17392 9766
rect 17448 9764 17472 9766
rect 17528 9764 17552 9766
rect 17608 9764 17614 9766
rect 17306 9755 17614 9764
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17592 9716 17644 9722
rect 17592 9658 17644 9664
rect 17500 9512 17552 9518
rect 17498 9480 17500 9489
rect 17552 9480 17554 9489
rect 17498 9415 17554 9424
rect 17222 9208 17278 9217
rect 17222 9143 17278 9152
rect 17236 9042 17264 9143
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 17500 9036 17552 9042
rect 17604 9024 17632 9658
rect 17552 8996 17632 9024
rect 17500 8978 17552 8984
rect 17328 8945 17356 8978
rect 17408 8968 17460 8974
rect 17314 8936 17370 8945
rect 17224 8900 17276 8906
rect 17408 8910 17460 8916
rect 17314 8871 17370 8880
rect 17224 8842 17276 8848
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16212 8492 16264 8498
rect 16316 8486 16712 8514
rect 16948 8560 17000 8566
rect 16948 8502 17000 8508
rect 16212 8434 16264 8440
rect 16028 8356 16080 8362
rect 16028 8298 16080 8304
rect 16224 8265 16252 8434
rect 16488 8424 16540 8430
rect 16486 8392 16488 8401
rect 16580 8424 16632 8430
rect 16540 8392 16542 8401
rect 16304 8356 16356 8362
rect 16356 8316 16436 8344
rect 16580 8366 16632 8372
rect 16486 8327 16542 8336
rect 16304 8298 16356 8304
rect 16210 8256 16266 8265
rect 16210 8191 16266 8200
rect 16408 8106 16436 8316
rect 15948 8078 16252 8106
rect 16408 8078 16528 8106
rect 15936 7676 15988 7682
rect 15988 7636 16114 7664
rect 15936 7618 15988 7624
rect 15154 7482 15206 7488
rect 15166 7344 15194 7482
rect 15350 7344 15378 7534
rect 15568 7540 15620 7546
rect 15672 7534 15746 7562
rect 15856 7534 15930 7562
rect 15568 7482 15620 7488
rect 15718 7344 15746 7534
rect 15902 7344 15930 7534
rect 16086 7344 16114 7636
rect 16224 7562 16252 8078
rect 16500 7954 16528 8078
rect 16396 7948 16448 7954
rect 16396 7890 16448 7896
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 16302 7712 16358 7721
rect 16302 7647 16304 7656
rect 16356 7647 16358 7656
rect 16408 7664 16436 7890
rect 16592 7721 16620 8366
rect 16684 7993 16712 8486
rect 16762 8120 16818 8129
rect 16762 8055 16818 8064
rect 16670 7984 16726 7993
rect 16670 7919 16726 7928
rect 16578 7712 16634 7721
rect 16408 7636 16482 7664
rect 16578 7647 16634 7656
rect 16304 7618 16356 7624
rect 16224 7534 16298 7562
rect 16270 7344 16298 7534
rect 16454 7344 16482 7636
rect 16626 7608 16678 7614
rect 16626 7550 16678 7556
rect 16776 7562 16804 8055
rect 17236 8022 17264 8842
rect 17316 8288 17368 8294
rect 17316 8230 17368 8236
rect 17132 8016 17184 8022
rect 17132 7958 17184 7964
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 16992 7576 17048 7585
rect 16638 7344 16666 7550
rect 16776 7534 16850 7562
rect 16822 7344 16850 7534
rect 16992 7511 17048 7520
rect 17144 7528 17172 7958
rect 17328 7562 17356 8230
rect 17420 7834 17448 8910
rect 17512 8265 17540 8978
rect 17696 8786 17724 10254
rect 18052 10202 18104 10208
rect 17776 10192 17828 10198
rect 17776 10134 17828 10140
rect 17788 9110 17816 10134
rect 17868 9920 17920 9926
rect 17868 9862 17920 9868
rect 17880 9722 17908 9862
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17866 9616 17922 9625
rect 18064 9586 18092 10202
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 17866 9551 17922 9560
rect 18052 9580 18104 9586
rect 17880 9466 17908 9551
rect 18052 9522 18104 9528
rect 18248 9466 18276 9998
rect 18420 9648 18472 9654
rect 18420 9590 18472 9596
rect 17880 9438 18000 9466
rect 18248 9438 18368 9466
rect 17868 9376 17920 9382
rect 17868 9318 17920 9324
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17776 8968 17828 8974
rect 17776 8910 17828 8916
rect 17604 8758 17724 8786
rect 17604 8634 17632 8758
rect 17682 8664 17738 8673
rect 17592 8628 17644 8634
rect 17682 8599 17738 8608
rect 17592 8570 17644 8576
rect 17696 8498 17724 8599
rect 17684 8492 17736 8498
rect 17684 8434 17736 8440
rect 17682 8392 17738 8401
rect 17682 8327 17684 8336
rect 17736 8327 17738 8336
rect 17684 8298 17736 8304
rect 17498 8256 17554 8265
rect 17498 8191 17554 8200
rect 17788 8129 17816 8910
rect 17880 8430 17908 9318
rect 17868 8424 17920 8430
rect 17868 8366 17920 8372
rect 17774 8120 17830 8129
rect 17774 8055 17830 8064
rect 17880 7993 17908 8366
rect 17972 8242 18000 9438
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18156 9042 18184 9318
rect 18144 9036 18196 9042
rect 18144 8978 18196 8984
rect 18156 8537 18184 8978
rect 18340 8922 18368 9438
rect 18432 9110 18460 9590
rect 18420 9104 18472 9110
rect 18420 9046 18472 9052
rect 18340 8894 18460 8922
rect 18142 8528 18198 8537
rect 18142 8463 18198 8472
rect 17972 8214 18276 8242
rect 17960 8016 18012 8022
rect 17866 7984 17922 7993
rect 17960 7958 18012 7964
rect 17866 7919 17922 7928
rect 17420 7806 17908 7834
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17512 7562 17540 7686
rect 17880 7585 17908 7806
rect 17866 7576 17922 7585
rect 17328 7534 17402 7562
rect 17512 7534 17586 7562
rect 17006 7344 17034 7511
rect 17144 7500 17212 7528
rect 13858 7304 13914 7313
rect 14416 7307 14472 7316
rect 13188 7262 13702 7290
rect 17184 7276 17212 7500
rect 17374 7344 17402 7534
rect 17558 7344 17586 7534
rect 17730 7540 17782 7546
rect 17972 7546 18000 7958
rect 18248 7562 18276 8214
rect 18432 7562 18460 8894
rect 18524 8634 18552 11478
rect 18616 10198 18644 11600
rect 18696 11552 18748 11558
rect 18696 11494 18748 11500
rect 18708 10266 18736 11494
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18604 10192 18656 10198
rect 18604 10134 18656 10140
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18708 9450 18736 9522
rect 18696 9444 18748 9450
rect 18696 9386 18748 9392
rect 18604 9376 18656 9382
rect 18604 9318 18656 9324
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18616 8430 18644 9318
rect 18604 8424 18656 8430
rect 18604 8366 18656 8372
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 17866 7511 17922 7520
rect 17960 7540 18012 7546
rect 17730 7482 17782 7488
rect 18248 7534 18322 7562
rect 18432 7534 18506 7562
rect 17960 7482 18012 7488
rect 17742 7344 17770 7482
rect 18294 7344 18322 7534
rect 18478 7344 18506 7534
rect 18616 7528 18644 8026
rect 18708 7886 18736 8026
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18800 7562 18828 10066
rect 18892 9654 18920 11600
rect 19168 9654 19196 11600
rect 19248 9920 19300 9926
rect 19248 9862 19300 9868
rect 18880 9648 18932 9654
rect 18880 9590 18932 9596
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 18972 9512 19024 9518
rect 18972 9454 19024 9460
rect 18984 9178 19012 9454
rect 18880 9172 18932 9178
rect 18880 9114 18932 9120
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 19064 9172 19116 9178
rect 19064 9114 19116 9120
rect 18892 8022 18920 9114
rect 18880 8016 18932 8022
rect 19076 7993 19104 9114
rect 19168 8634 19196 9590
rect 19260 9042 19288 9862
rect 19444 9518 19472 11600
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 19628 9518 19656 9862
rect 19720 9654 19748 11600
rect 19996 10266 20024 11600
rect 19984 10260 20036 10266
rect 19984 10202 20036 10208
rect 19800 10192 19852 10198
rect 19800 10134 19852 10140
rect 19708 9648 19760 9654
rect 19708 9590 19760 9596
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 19616 9512 19668 9518
rect 19616 9454 19668 9460
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19524 9376 19576 9382
rect 19524 9318 19576 9324
rect 19248 9036 19300 9042
rect 19248 8978 19300 8984
rect 19260 8945 19288 8978
rect 19246 8936 19302 8945
rect 19246 8871 19302 8880
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19352 8514 19380 9318
rect 19432 9036 19484 9042
rect 19432 8978 19484 8984
rect 19444 8945 19472 8978
rect 19430 8936 19486 8945
rect 19430 8871 19486 8880
rect 19430 8528 19486 8537
rect 19352 8486 19430 8514
rect 19430 8463 19486 8472
rect 19444 8430 19472 8463
rect 19432 8424 19484 8430
rect 19536 8401 19564 9318
rect 19432 8366 19484 8372
rect 19522 8392 19578 8401
rect 19522 8327 19578 8336
rect 19628 8276 19656 9454
rect 19720 8634 19748 9590
rect 19812 9110 19840 10134
rect 19892 9920 19944 9926
rect 19892 9862 19944 9868
rect 19800 9104 19852 9110
rect 19800 9046 19852 9052
rect 19904 9042 19932 9862
rect 19996 9586 20024 10202
rect 20272 9738 20300 11600
rect 20548 10282 20576 11600
rect 20456 10254 20576 10282
rect 20456 10198 20484 10254
rect 20444 10192 20496 10198
rect 20444 10134 20496 10140
rect 20824 10130 20852 11600
rect 20996 10260 21048 10266
rect 20996 10202 21048 10208
rect 20352 10124 20404 10130
rect 20352 10066 20404 10072
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20180 9710 20300 9738
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 20180 9450 20208 9710
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 19984 9376 20036 9382
rect 19984 9318 20036 9324
rect 19996 9178 20024 9318
rect 19984 9172 20036 9178
rect 19984 9114 20036 9120
rect 19892 9036 19944 9042
rect 19892 8978 19944 8984
rect 19996 8945 20024 9114
rect 19982 8936 20038 8945
rect 19982 8871 20038 8880
rect 19800 8832 19852 8838
rect 19800 8774 19852 8780
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19444 8248 19656 8276
rect 18880 7958 18932 7964
rect 19062 7984 19118 7993
rect 19062 7919 19118 7928
rect 18970 7848 19026 7857
rect 18970 7783 19026 7792
rect 19156 7812 19208 7818
rect 18984 7562 19012 7783
rect 19156 7754 19208 7760
rect 19168 7562 19196 7754
rect 18800 7534 18874 7562
rect 18984 7534 19058 7562
rect 19168 7534 19242 7562
rect 18616 7500 18684 7528
rect 18656 7276 18684 7500
rect 18846 7344 18874 7534
rect 19030 7344 19058 7534
rect 19214 7344 19242 7534
rect 19444 7528 19472 8248
rect 19812 8090 19840 8774
rect 19892 8356 19944 8362
rect 19892 8298 19944 8304
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19800 8084 19852 8090
rect 19800 8026 19852 8032
rect 19536 7562 19564 8026
rect 19904 7886 19932 8298
rect 19892 7880 19944 7886
rect 19892 7822 19944 7828
rect 20088 7698 20116 9386
rect 20180 8362 20208 9386
rect 20364 9110 20392 10066
rect 20536 9988 20588 9994
rect 20536 9930 20588 9936
rect 20352 9104 20404 9110
rect 20352 9046 20404 9052
rect 20442 9072 20498 9081
rect 20548 9042 20576 9930
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20732 9518 20760 9862
rect 20720 9512 20772 9518
rect 20720 9454 20772 9460
rect 20442 9007 20498 9016
rect 20536 9036 20588 9042
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20272 8566 20300 8910
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20260 8560 20312 8566
rect 20260 8502 20312 8508
rect 20364 8498 20392 8774
rect 20456 8514 20484 9007
rect 20536 8978 20588 8984
rect 20548 8945 20576 8978
rect 20534 8936 20590 8945
rect 20534 8871 20590 8880
rect 20732 8650 20760 9454
rect 20812 9444 20864 9450
rect 20812 9386 20864 9392
rect 20904 9444 20956 9450
rect 20904 9386 20956 9392
rect 20640 8622 20760 8650
rect 20352 8492 20404 8498
rect 20456 8486 20576 8514
rect 20352 8434 20404 8440
rect 20444 8424 20496 8430
rect 20442 8392 20444 8401
rect 20496 8392 20498 8401
rect 20168 8356 20220 8362
rect 20442 8327 20498 8336
rect 20168 8298 20220 8304
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 19996 7670 20116 7698
rect 19754 7608 19806 7614
rect 19536 7534 19604 7562
rect 19996 7562 20024 7670
rect 19754 7550 19806 7556
rect 19306 7500 19472 7528
rect 19306 7449 19334 7500
rect 19292 7440 19348 7449
rect 19292 7375 19348 7384
rect 19378 7304 19434 7313
rect 13858 7239 13914 7248
rect 19576 7276 19604 7534
rect 19766 7344 19794 7550
rect 19950 7534 20024 7562
rect 20272 7562 20300 7958
rect 20548 7562 20576 8486
rect 20640 8242 20668 8622
rect 20720 8424 20772 8430
rect 20718 8392 20720 8401
rect 20772 8392 20774 8401
rect 20718 8327 20774 8336
rect 20640 8214 20760 8242
rect 20732 8129 20760 8214
rect 20718 8120 20774 8129
rect 20718 8055 20774 8064
rect 20824 7954 20852 9386
rect 20916 9110 20944 9386
rect 21008 9110 21036 10202
rect 21100 9586 21128 11600
rect 21376 10266 21404 11600
rect 21364 10260 21416 10266
rect 21364 10202 21416 10208
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21270 9344 21326 9353
rect 21270 9279 21326 9288
rect 20904 9104 20956 9110
rect 20904 9046 20956 9052
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 21088 9036 21140 9042
rect 21088 8978 21140 8984
rect 20902 8800 20958 8809
rect 20902 8735 20958 8744
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20812 7948 20864 7954
rect 20812 7890 20864 7896
rect 20122 7540 20174 7546
rect 19950 7344 19978 7534
rect 20272 7534 20340 7562
rect 20122 7482 20174 7488
rect 20134 7344 20162 7482
rect 20312 7276 20340 7534
rect 20502 7534 20576 7562
rect 20640 7562 20668 7890
rect 20916 7562 20944 8735
rect 20996 8288 21048 8294
rect 20996 8230 21048 8236
rect 20640 7534 20708 7562
rect 20502 7344 20530 7534
rect 20680 7276 20708 7534
rect 20824 7534 20944 7562
rect 21008 7562 21036 8230
rect 21100 8022 21128 8978
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21192 8294 21220 8366
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21178 7848 21234 7857
rect 21178 7783 21234 7792
rect 21192 7596 21220 7783
rect 21284 7698 21312 9279
rect 21376 8430 21404 9522
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21364 8424 21416 8430
rect 21364 8366 21416 8372
rect 21468 7750 21496 8434
rect 21456 7744 21508 7750
rect 21284 7670 21404 7698
rect 21456 7686 21508 7692
rect 21560 7698 21588 9658
rect 21652 9586 21680 11600
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21652 9110 21680 9522
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21640 9104 21692 9110
rect 21640 9046 21692 9052
rect 21744 9042 21772 9318
rect 21732 9036 21784 9042
rect 21732 8978 21784 8984
rect 21744 8537 21772 8978
rect 21928 8634 21956 11600
rect 22204 9654 22232 11600
rect 22192 9648 22244 9654
rect 22192 9590 22244 9596
rect 22204 9110 22232 9590
rect 22282 9480 22338 9489
rect 22282 9415 22338 9424
rect 22192 9104 22244 9110
rect 22192 9046 22244 9052
rect 22008 8900 22060 8906
rect 22008 8842 22060 8848
rect 22020 8809 22048 8842
rect 22006 8800 22062 8809
rect 22006 8735 22062 8744
rect 22098 8664 22154 8673
rect 21916 8628 21968 8634
rect 22098 8599 22154 8608
rect 21916 8570 21968 8576
rect 22008 8560 22060 8566
rect 21730 8528 21786 8537
rect 22008 8502 22060 8508
rect 21730 8463 21786 8472
rect 21732 8424 21784 8430
rect 21730 8392 21732 8401
rect 21824 8424 21876 8430
rect 21784 8392 21786 8401
rect 21876 8384 21956 8412
rect 21824 8366 21876 8372
rect 21730 8327 21786 8336
rect 21560 7670 21772 7698
rect 21192 7568 21266 7596
rect 21008 7534 21076 7562
rect 20824 7358 20852 7534
rect 20824 7330 20892 7358
rect 20864 7276 20892 7330
rect 21048 7276 21076 7534
rect 21238 7344 21266 7568
rect 21376 7562 21404 7670
rect 21594 7608 21646 7614
rect 21376 7534 21450 7562
rect 21594 7550 21646 7556
rect 21744 7562 21772 7670
rect 21928 7585 21956 8384
rect 21914 7576 21970 7585
rect 21422 7344 21450 7534
rect 21606 7344 21634 7550
rect 21744 7534 21818 7562
rect 21790 7344 21818 7534
rect 22020 7546 22048 8502
rect 22112 7596 22140 8599
rect 22112 7568 22186 7596
rect 21914 7511 21970 7520
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21960 7372 22016 7381
rect 22158 7344 22186 7568
rect 22296 7358 22324 9415
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22388 8673 22416 9114
rect 22374 8664 22430 8673
rect 22374 8599 22430 8608
rect 22480 8498 22508 11600
rect 22756 9654 22784 11600
rect 22744 9648 22796 9654
rect 22744 9590 22796 9596
rect 22560 9444 22612 9450
rect 22560 9386 22612 9392
rect 22572 9353 22600 9386
rect 22558 9344 22614 9353
rect 22558 9279 22614 9288
rect 22572 9110 22600 9279
rect 22650 9208 22706 9217
rect 22650 9143 22706 9152
rect 22560 9104 22612 9110
rect 22560 9046 22612 9052
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22480 7596 22508 7822
rect 22664 7596 22692 9143
rect 22756 8634 22784 9590
rect 23032 9586 23060 11600
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 23020 9580 23072 9586
rect 23020 9522 23072 9528
rect 22940 9489 22968 9522
rect 22926 9480 22982 9489
rect 22926 9415 22982 9424
rect 23032 9110 23060 9522
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 23112 8900 23164 8906
rect 23112 8842 23164 8848
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 23020 8424 23072 8430
rect 23018 8392 23020 8401
rect 23072 8392 23074 8401
rect 23018 8327 23074 8336
rect 22834 8256 22890 8265
rect 22834 8191 22890 8200
rect 22848 7596 22876 8191
rect 23124 7596 23152 8842
rect 23308 8537 23336 11600
rect 23584 9654 23612 11600
rect 23572 9648 23624 9654
rect 23572 9590 23624 9596
rect 23480 8968 23532 8974
rect 23480 8910 23532 8916
rect 23388 8832 23440 8838
rect 23388 8774 23440 8780
rect 23294 8528 23350 8537
rect 23294 8463 23350 8472
rect 23204 8084 23256 8090
rect 23204 8026 23256 8032
rect 22480 7568 22554 7596
rect 22664 7568 22738 7596
rect 22848 7568 22922 7596
rect 22296 7330 22364 7358
rect 22526 7344 22554 7568
rect 22710 7344 22738 7568
rect 22894 7344 22922 7568
rect 23078 7568 23152 7596
rect 23216 7596 23244 8026
rect 23400 7596 23428 8774
rect 23492 8090 23520 8910
rect 23584 8838 23612 9590
rect 23860 9466 23888 11600
rect 24136 9738 24164 11600
rect 24308 11212 24360 11218
rect 24308 11154 24360 11160
rect 24216 11008 24268 11014
rect 24216 10950 24268 10956
rect 24044 9710 24164 9738
rect 24044 9586 24072 9710
rect 24032 9580 24084 9586
rect 24032 9522 24084 9528
rect 23860 9438 23980 9466
rect 23756 9376 23808 9382
rect 23756 9318 23808 9324
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23768 9042 23796 9318
rect 23756 9036 23808 9042
rect 23756 8978 23808 8984
rect 23768 8945 23796 8978
rect 23754 8936 23810 8945
rect 23860 8906 23888 9318
rect 23754 8871 23810 8880
rect 23848 8900 23900 8906
rect 23848 8842 23900 8848
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23860 8129 23888 8842
rect 23952 8498 23980 9438
rect 24044 9110 24072 9522
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24032 9104 24084 9110
rect 24032 9046 24084 9052
rect 24030 8800 24086 8809
rect 24030 8735 24086 8744
rect 23940 8492 23992 8498
rect 23940 8434 23992 8440
rect 23952 8294 23980 8434
rect 23940 8288 23992 8294
rect 23940 8230 23992 8236
rect 24044 8242 24072 8735
rect 24136 8430 24164 9454
rect 24124 8424 24176 8430
rect 24122 8392 24124 8401
rect 24176 8392 24178 8401
rect 24122 8327 24178 8336
rect 24044 8214 24164 8242
rect 23846 8120 23902 8129
rect 23480 8084 23532 8090
rect 23846 8055 23902 8064
rect 23480 8026 23532 8032
rect 23938 7984 23994 7993
rect 23938 7919 23994 7928
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23584 7596 23612 7686
rect 23802 7608 23854 7614
rect 23216 7568 23290 7596
rect 23400 7568 23474 7596
rect 23584 7568 23658 7596
rect 23078 7344 23106 7568
rect 23262 7344 23290 7568
rect 23446 7344 23474 7568
rect 23630 7344 23658 7568
rect 23952 7596 23980 7919
rect 23952 7568 24026 7596
rect 23802 7550 23854 7556
rect 23814 7344 23842 7550
rect 23998 7344 24026 7568
rect 24136 7358 24164 8214
rect 24228 7585 24256 10950
rect 24320 10606 24348 11154
rect 24308 10600 24360 10606
rect 24308 10542 24360 10548
rect 24320 10130 24348 10542
rect 24308 10124 24360 10130
rect 24308 10066 24360 10072
rect 24412 8673 24440 11600
rect 24492 10464 24544 10470
rect 24492 10406 24544 10412
rect 24504 9761 24532 10406
rect 24688 10010 24716 11600
rect 24860 10464 24912 10470
rect 24860 10406 24912 10412
rect 24688 9982 24808 10010
rect 24676 9920 24728 9926
rect 24676 9862 24728 9868
rect 24688 9761 24716 9862
rect 24490 9752 24546 9761
rect 24490 9687 24546 9696
rect 24674 9752 24730 9761
rect 24674 9687 24730 9696
rect 24780 9654 24808 9982
rect 24492 9648 24544 9654
rect 24492 9590 24544 9596
rect 24768 9648 24820 9654
rect 24768 9590 24820 9596
rect 24398 8664 24454 8673
rect 24398 8599 24454 8608
rect 24306 8528 24362 8537
rect 24306 8463 24362 8472
rect 24320 8344 24348 8463
rect 24400 8356 24452 8362
rect 24320 8316 24400 8344
rect 24400 8298 24452 8304
rect 24504 8242 24532 9590
rect 24582 9480 24638 9489
rect 24582 9415 24638 9424
rect 24412 8214 24532 8242
rect 24412 7596 24440 8214
rect 24214 7576 24270 7585
rect 24214 7511 24270 7520
rect 24366 7568 24440 7596
rect 24136 7330 24204 7358
rect 24366 7344 24394 7568
rect 24596 7562 24624 9415
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24688 9217 24716 9318
rect 24674 9208 24730 9217
rect 24674 9143 24730 9152
rect 24688 9110 24716 9143
rect 24780 9110 24808 9590
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24768 9104 24820 9110
rect 24768 9046 24820 9052
rect 24676 8968 24728 8974
rect 24676 8910 24728 8916
rect 24688 8362 24716 8910
rect 24676 8356 24728 8362
rect 24676 8298 24728 8304
rect 24688 8129 24716 8298
rect 24674 8120 24730 8129
rect 24674 8055 24730 8064
rect 24676 8016 24728 8022
rect 24676 7958 24728 7964
rect 24688 7596 24716 7958
rect 24688 7568 24756 7596
rect 24872 7585 24900 10406
rect 24964 9674 24992 11600
rect 25240 11098 25268 11600
rect 25516 11354 25544 11600
rect 25504 11348 25556 11354
rect 25504 11290 25556 11296
rect 25240 11070 25728 11098
rect 25228 11008 25280 11014
rect 25228 10950 25280 10956
rect 25136 10464 25188 10470
rect 25136 10406 25188 10412
rect 24964 9646 25084 9674
rect 25056 8974 25084 9646
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25042 8664 25098 8673
rect 25042 8599 25098 8608
rect 25056 8430 25084 8599
rect 24952 8424 25004 8430
rect 24952 8366 25004 8372
rect 25044 8424 25096 8430
rect 25044 8366 25096 8372
rect 24964 7614 24992 8366
rect 25044 8084 25096 8090
rect 25044 8026 25096 8032
rect 24952 7608 25004 7614
rect 24550 7534 24624 7562
rect 24550 7344 24578 7534
rect 21960 7307 22016 7316
rect 22336 7276 22364 7330
rect 24176 7276 24204 7330
rect 24728 7276 24756 7568
rect 24858 7576 24914 7585
rect 24952 7550 25004 7556
rect 24858 7511 24914 7520
rect 25056 7528 25084 8026
rect 25148 7857 25176 10406
rect 25134 7848 25190 7857
rect 25134 7783 25190 7792
rect 25240 7721 25268 10950
rect 25306 10908 25614 10917
rect 25306 10906 25312 10908
rect 25368 10906 25392 10908
rect 25448 10906 25472 10908
rect 25528 10906 25552 10908
rect 25608 10906 25614 10908
rect 25368 10854 25370 10906
rect 25550 10854 25552 10906
rect 25306 10852 25312 10854
rect 25368 10852 25392 10854
rect 25448 10852 25472 10854
rect 25528 10852 25552 10854
rect 25608 10852 25614 10854
rect 25306 10843 25614 10852
rect 25306 9820 25614 9829
rect 25306 9818 25312 9820
rect 25368 9818 25392 9820
rect 25448 9818 25472 9820
rect 25528 9818 25552 9820
rect 25608 9818 25614 9820
rect 25368 9766 25370 9818
rect 25550 9766 25552 9818
rect 25306 9764 25312 9766
rect 25368 9764 25392 9766
rect 25448 9764 25472 9766
rect 25528 9764 25552 9766
rect 25608 9764 25614 9766
rect 25306 9755 25614 9764
rect 25700 9738 25728 11070
rect 25792 10810 25820 11600
rect 26068 11558 26096 11600
rect 25872 11552 25924 11558
rect 25872 11494 25924 11500
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 25780 10804 25832 10810
rect 25780 10746 25832 10752
rect 25884 10266 25912 11494
rect 25946 11452 26254 11461
rect 25946 11450 25952 11452
rect 26008 11450 26032 11452
rect 26088 11450 26112 11452
rect 26168 11450 26192 11452
rect 26248 11450 26254 11452
rect 26008 11398 26010 11450
rect 26190 11398 26192 11450
rect 25946 11396 25952 11398
rect 26008 11396 26032 11398
rect 26088 11396 26112 11398
rect 26168 11396 26192 11398
rect 26248 11396 26254 11398
rect 25946 11387 26254 11396
rect 25964 11212 26016 11218
rect 26240 11212 26292 11218
rect 26016 11172 26240 11200
rect 25964 11154 26016 11160
rect 26240 11154 26292 11160
rect 26252 10452 26280 11154
rect 26344 10742 26372 11600
rect 26424 11008 26476 11014
rect 26424 10950 26476 10956
rect 26332 10736 26384 10742
rect 26332 10678 26384 10684
rect 26252 10424 26372 10452
rect 25946 10364 26254 10373
rect 25946 10362 25952 10364
rect 26008 10362 26032 10364
rect 26088 10362 26112 10364
rect 26168 10362 26192 10364
rect 26248 10362 26254 10364
rect 26008 10310 26010 10362
rect 26190 10310 26192 10362
rect 25946 10308 25952 10310
rect 26008 10308 26032 10310
rect 26088 10308 26112 10310
rect 26168 10308 26192 10310
rect 26248 10308 26254 10310
rect 25946 10299 26254 10308
rect 25872 10260 25924 10266
rect 25872 10202 25924 10208
rect 26344 10130 26372 10424
rect 26332 10124 26384 10130
rect 26332 10066 26384 10072
rect 25700 9710 25820 9738
rect 25412 9444 25464 9450
rect 25412 9386 25464 9392
rect 25424 9081 25452 9386
rect 25410 9072 25466 9081
rect 25410 9007 25466 9016
rect 25594 8800 25650 8809
rect 25594 8735 25650 8744
rect 25412 8628 25464 8634
rect 25412 8570 25464 8576
rect 25226 7712 25282 7721
rect 25226 7647 25282 7656
rect 25424 7596 25452 8570
rect 25504 8424 25556 8430
rect 25504 8366 25556 8372
rect 25516 8265 25544 8366
rect 25502 8256 25558 8265
rect 25502 8191 25558 8200
rect 25608 7596 25636 8735
rect 25792 8634 25820 9710
rect 25964 9172 26016 9178
rect 25964 9114 26016 9120
rect 25870 9072 25926 9081
rect 25870 9007 25872 9016
rect 25924 9007 25926 9016
rect 25872 8978 25924 8984
rect 25780 8628 25832 8634
rect 25780 8570 25832 8576
rect 25870 8528 25926 8537
rect 25870 8463 25872 8472
rect 25924 8463 25926 8472
rect 25872 8434 25924 8440
rect 25826 7608 25878 7614
rect 25424 7568 25492 7596
rect 25608 7568 25676 7596
rect 25274 7540 25326 7546
rect 25056 7500 25124 7528
rect 24898 7304 24954 7313
rect 19378 7239 19434 7248
rect 25096 7276 25124 7500
rect 25274 7482 25326 7488
rect 25286 7344 25314 7482
rect 25464 7276 25492 7568
rect 25648 7276 25676 7568
rect 25976 7596 26004 9114
rect 26240 8832 26292 8838
rect 26240 8774 26292 8780
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 26148 8560 26200 8566
rect 26148 8502 26200 8508
rect 26160 7596 26188 8502
rect 26252 7698 26280 8774
rect 26344 8673 26372 8774
rect 26330 8664 26386 8673
rect 26330 8599 26386 8608
rect 26252 7670 26372 7698
rect 25976 7568 26044 7596
rect 26160 7568 26228 7596
rect 25826 7550 25878 7556
rect 25838 7344 25866 7550
rect 26016 7276 26044 7568
rect 26200 7276 26228 7568
rect 26344 7358 26372 7670
rect 26436 7585 26464 10950
rect 26620 10674 26648 11600
rect 26896 11354 26924 11600
rect 26884 11348 26936 11354
rect 26884 11290 26936 11296
rect 27172 11150 27200 11600
rect 27448 11354 27476 11600
rect 27436 11348 27488 11354
rect 27436 11290 27488 11296
rect 27528 11212 27580 11218
rect 27528 11154 27580 11160
rect 27160 11144 27212 11150
rect 27160 11086 27212 11092
rect 26608 10668 26660 10674
rect 26608 10610 26660 10616
rect 27540 10606 27568 11154
rect 27160 10600 27212 10606
rect 27160 10542 27212 10548
rect 27528 10600 27580 10606
rect 27528 10542 27580 10548
rect 27724 10554 27752 11600
rect 27896 11008 27948 11014
rect 27896 10950 27948 10956
rect 27172 10130 27200 10542
rect 27724 10526 27844 10554
rect 27712 10464 27764 10470
rect 27712 10406 27764 10412
rect 27160 10124 27212 10130
rect 27160 10066 27212 10072
rect 27344 10124 27396 10130
rect 27344 10066 27396 10072
rect 27356 10033 27384 10066
rect 27342 10024 27398 10033
rect 27342 9959 27398 9968
rect 26976 9920 27028 9926
rect 26976 9862 27028 9868
rect 27252 9920 27304 9926
rect 27252 9862 27304 9868
rect 27620 9920 27672 9926
rect 27620 9862 27672 9868
rect 26608 9104 26660 9110
rect 26660 9064 26740 9092
rect 26608 9046 26660 9052
rect 26516 8424 26568 8430
rect 26516 8366 26568 8372
rect 26608 8424 26660 8430
rect 26608 8366 26660 8372
rect 26528 7596 26556 8366
rect 26620 7721 26648 8366
rect 26606 7712 26662 7721
rect 26606 7647 26662 7656
rect 26712 7596 26740 9064
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26792 8832 26844 8838
rect 26792 8774 26844 8780
rect 26804 8401 26832 8774
rect 26790 8392 26846 8401
rect 26790 8327 26846 8336
rect 26896 7596 26924 8842
rect 26988 8673 27016 9862
rect 26974 8664 27030 8673
rect 26974 8599 27030 8608
rect 27068 8424 27120 8430
rect 27068 8366 27120 8372
rect 27080 7596 27108 8366
rect 27264 8362 27292 9862
rect 27632 8537 27660 9862
rect 27618 8528 27674 8537
rect 27618 8463 27674 8472
rect 27252 8356 27304 8362
rect 27252 8298 27304 8304
rect 27526 7984 27582 7993
rect 27526 7919 27582 7928
rect 27540 7596 27568 7919
rect 27724 7857 27752 10406
rect 27816 9178 27844 10526
rect 27804 9172 27856 9178
rect 27804 9114 27856 9120
rect 27908 8809 27936 10950
rect 28000 10266 28028 11600
rect 28172 11008 28224 11014
rect 28172 10950 28224 10956
rect 27988 10260 28040 10266
rect 27988 10202 28040 10208
rect 28080 9988 28132 9994
rect 28080 9930 28132 9936
rect 28092 9518 28120 9930
rect 28080 9512 28132 9518
rect 28080 9454 28132 9460
rect 28092 8974 28120 9454
rect 28080 8968 28132 8974
rect 28184 8945 28212 10950
rect 28276 10062 28304 11600
rect 28552 10266 28580 11600
rect 28632 11348 28684 11354
rect 28632 11290 28684 11296
rect 28644 11218 28672 11290
rect 28632 11212 28684 11218
rect 28684 11172 28764 11200
rect 28632 11154 28684 11160
rect 28736 11014 28764 11172
rect 28632 11008 28684 11014
rect 28632 10950 28684 10956
rect 28724 11008 28776 11014
rect 28724 10950 28776 10956
rect 28540 10260 28592 10266
rect 28540 10202 28592 10208
rect 28264 10056 28316 10062
rect 28262 10024 28264 10033
rect 28316 10024 28318 10033
rect 28262 9959 28318 9968
rect 28356 9376 28408 9382
rect 28356 9318 28408 9324
rect 28080 8910 28132 8916
rect 28170 8936 28226 8945
rect 28170 8871 28226 8880
rect 27894 8800 27950 8809
rect 27894 8735 27950 8744
rect 28368 8537 28396 9318
rect 28354 8528 28410 8537
rect 28354 8463 28410 8472
rect 27894 8120 27950 8129
rect 27894 8055 27950 8064
rect 27710 7848 27766 7857
rect 27710 7783 27766 7792
rect 27710 7712 27766 7721
rect 27710 7647 27766 7656
rect 27724 7596 27752 7647
rect 27908 7596 27936 8055
rect 26422 7576 26478 7585
rect 26528 7568 26596 7596
rect 26712 7568 26786 7596
rect 26896 7568 26964 7596
rect 27080 7568 27148 7596
rect 26422 7511 26478 7520
rect 26344 7330 26412 7358
rect 26384 7276 26412 7330
rect 26568 7276 26596 7568
rect 26758 7344 26786 7568
rect 26936 7276 26964 7568
rect 27120 7276 27148 7568
rect 27494 7568 27568 7596
rect 27678 7568 27752 7596
rect 27862 7568 27936 7596
rect 28402 7608 28454 7614
rect 27298 7540 27350 7546
rect 27298 7482 27350 7488
rect 27310 7344 27338 7482
rect 27494 7344 27522 7568
rect 27678 7344 27706 7568
rect 27862 7344 27890 7568
rect 28644 7585 28672 10950
rect 28828 10810 28856 11600
rect 29104 11150 29132 11600
rect 29380 11354 29408 11600
rect 29368 11348 29420 11354
rect 29368 11290 29420 11296
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 29184 11076 29236 11082
rect 29184 11018 29236 11024
rect 28816 10804 28868 10810
rect 28816 10746 28868 10752
rect 29000 9920 29052 9926
rect 29000 9862 29052 9868
rect 29012 8401 29040 9862
rect 29196 8401 29224 11018
rect 29552 11008 29604 11014
rect 29552 10950 29604 10956
rect 29564 10742 29592 10950
rect 29552 10736 29604 10742
rect 29552 10678 29604 10684
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29564 9926 29592 9998
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 29552 9920 29604 9926
rect 29552 9862 29604 9868
rect 29288 9761 29316 9862
rect 29274 9752 29330 9761
rect 29274 9687 29330 9696
rect 29656 9654 29684 11600
rect 29932 11354 29960 11600
rect 30104 11552 30156 11558
rect 30104 11494 30156 11500
rect 30116 11354 30144 11494
rect 29920 11348 29972 11354
rect 29920 11290 29972 11296
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 29828 11008 29880 11014
rect 29828 10950 29880 10956
rect 29644 9648 29696 9654
rect 29644 9590 29696 9596
rect 28998 8392 29054 8401
rect 28998 8327 29054 8336
rect 29182 8392 29238 8401
rect 29182 8327 29238 8336
rect 29840 8265 29868 10950
rect 30012 10464 30064 10470
rect 30012 10406 30064 10412
rect 30024 10198 30052 10406
rect 30012 10192 30064 10198
rect 30012 10134 30064 10140
rect 30208 10062 30236 11600
rect 30484 11098 30512 11600
rect 30760 11558 30788 11600
rect 30748 11552 30800 11558
rect 30748 11494 30800 11500
rect 30932 11348 30984 11354
rect 31036 11336 31064 11600
rect 30984 11308 31064 11336
rect 31116 11348 31168 11354
rect 30932 11290 30984 11296
rect 31116 11290 31168 11296
rect 30656 11212 30708 11218
rect 30656 11154 30708 11160
rect 30840 11212 30892 11218
rect 31128 11200 31156 11290
rect 30892 11172 31156 11200
rect 30840 11154 30892 11160
rect 30392 11070 30512 11098
rect 30196 10056 30248 10062
rect 30196 9998 30248 10004
rect 30392 9926 30420 11070
rect 30472 11008 30524 11014
rect 30472 10950 30524 10956
rect 30484 10810 30512 10950
rect 30472 10804 30524 10810
rect 30472 10746 30524 10752
rect 30668 10606 30696 11154
rect 31208 10736 31260 10742
rect 31208 10678 31260 10684
rect 30656 10600 30708 10606
rect 30656 10542 30708 10548
rect 30840 10260 30892 10266
rect 30840 10202 30892 10208
rect 30852 10130 30880 10202
rect 30840 10124 30892 10130
rect 30840 10066 30892 10072
rect 31116 10124 31168 10130
rect 31116 10066 31168 10072
rect 31128 9926 31156 10066
rect 30380 9920 30432 9926
rect 30748 9920 30800 9926
rect 30380 9862 30432 9868
rect 30746 9888 30748 9897
rect 31116 9920 31168 9926
rect 30800 9888 30802 9897
rect 31116 9862 31168 9868
rect 30746 9823 30802 9832
rect 29826 8256 29882 8265
rect 29826 8191 29882 8200
rect 30746 8120 30802 8129
rect 29184 8084 29236 8090
rect 30746 8055 30802 8064
rect 29184 8026 29236 8032
rect 28814 7848 28870 7857
rect 28814 7783 28870 7792
rect 28828 7596 28856 7783
rect 29196 7596 29224 8026
rect 30104 8016 30156 8022
rect 30104 7958 30156 7964
rect 29368 7880 29420 7886
rect 29368 7822 29420 7828
rect 29380 7596 29408 7822
rect 29920 7812 29972 7818
rect 29920 7754 29972 7760
rect 29552 7744 29604 7750
rect 29552 7686 29604 7692
rect 29564 7596 29592 7686
rect 29932 7596 29960 7754
rect 30116 7596 30144 7958
rect 30760 7857 30788 8055
rect 30746 7848 30802 7857
rect 31220 7834 31248 10678
rect 31312 9994 31340 11600
rect 31392 11552 31444 11558
rect 31392 11494 31444 11500
rect 31404 10266 31432 11494
rect 31588 11098 31616 11600
rect 31850 11600 31906 12000
rect 32126 11600 32182 12000
rect 32402 11600 32458 12000
rect 32678 11620 32734 12000
rect 32678 11600 32680 11620
rect 31760 11562 31812 11568
rect 31772 11286 31800 11562
rect 31864 11354 31892 11600
rect 32140 11558 32168 11600
rect 32128 11552 32180 11558
rect 32128 11494 32180 11500
rect 32220 11552 32272 11558
rect 32220 11494 32272 11500
rect 31852 11348 31904 11354
rect 31852 11290 31904 11296
rect 31760 11280 31812 11286
rect 31760 11222 31812 11228
rect 32036 11212 32088 11218
rect 32036 11154 32088 11160
rect 31496 11082 31616 11098
rect 31484 11076 31616 11082
rect 31536 11070 31616 11076
rect 31484 11018 31536 11024
rect 31852 11008 31904 11014
rect 31852 10950 31904 10956
rect 31944 11008 31996 11014
rect 31944 10950 31996 10956
rect 31668 10600 31720 10606
rect 31668 10542 31720 10548
rect 31392 10260 31444 10266
rect 31392 10202 31444 10208
rect 31680 10130 31708 10542
rect 31668 10124 31720 10130
rect 31668 10066 31720 10072
rect 31300 9988 31352 9994
rect 31300 9930 31352 9936
rect 31864 8514 31892 10950
rect 31772 8486 31892 8514
rect 31666 7984 31722 7993
rect 31666 7919 31722 7928
rect 31220 7806 31616 7834
rect 30746 7783 30802 7792
rect 31482 7712 31538 7721
rect 31482 7647 31538 7656
rect 28402 7550 28454 7556
rect 28630 7576 28686 7585
rect 28216 7372 28272 7381
rect 28414 7344 28442 7550
rect 28630 7511 28686 7520
rect 28782 7568 28856 7596
rect 29150 7568 29224 7596
rect 29334 7568 29408 7596
rect 29518 7568 29592 7596
rect 29886 7568 29960 7596
rect 30070 7568 30144 7596
rect 30840 7608 30892 7614
rect 28782 7344 28810 7568
rect 28954 7540 29006 7546
rect 28954 7482 29006 7488
rect 28966 7344 28994 7482
rect 29150 7344 29178 7568
rect 29334 7344 29362 7568
rect 29518 7344 29546 7568
rect 29886 7344 29914 7568
rect 30070 7344 30098 7568
rect 30840 7550 30892 7556
rect 30852 7449 30880 7550
rect 30838 7440 30894 7449
rect 30838 7375 30894 7384
rect 28216 7307 28272 7316
rect 29688 7304 29744 7313
rect 24898 7239 24954 7248
rect 29688 7239 29744 7248
rect 14042 7168 14098 7177
rect 14042 7103 14098 7112
rect 28584 7168 28640 7177
rect 14968 7100 15024 7109
rect 14968 7035 15024 7044
rect 15520 7100 15576 7109
rect 15520 7035 15576 7044
rect 17912 7100 17968 7109
rect 17912 7035 17968 7044
rect 18096 7100 18152 7109
rect 18096 7035 18152 7044
rect 28032 7100 28088 7109
rect 28584 7103 28640 7112
rect 28032 7035 28088 7044
rect 30240 7100 30296 7109
rect 30240 7035 30296 7044
rect 31496 6662 31524 7647
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 31484 6656 31536 6662
rect 31484 6598 31536 6604
rect 12990 5400 13046 5409
rect 12990 5335 13046 5344
rect 13004 400 13032 5335
rect 13542 4584 13598 4593
rect 13542 4519 13598 4528
rect 14646 4584 14702 4593
rect 14646 4519 14702 4528
rect 14922 4584 14978 4593
rect 14922 4519 14978 4528
rect 15474 4584 15530 4593
rect 15474 4519 15530 4528
rect 16302 4584 16358 4593
rect 16302 4519 16358 4528
rect 16578 4584 16634 4593
rect 16578 4519 16634 4528
rect 19338 4584 19394 4593
rect 19338 4519 19394 4528
rect 22650 4584 22706 4593
rect 22650 4519 22706 4528
rect 24950 4584 25006 4593
rect 24950 4519 25006 4528
rect 26146 4584 26202 4593
rect 26146 4519 26202 4528
rect 30654 4584 30710 4593
rect 30654 4519 30710 4528
rect 13266 4448 13322 4457
rect 13266 4383 13322 4392
rect 13280 400 13308 4383
rect 13556 400 13584 4519
rect 14370 4448 14426 4457
rect 14370 4383 14426 4392
rect 13818 1184 13874 1193
rect 13818 1119 13874 1128
rect 13832 400 13860 1119
rect 14094 1048 14150 1057
rect 14094 983 14150 992
rect 14108 400 14136 983
rect 14384 400 14412 4383
rect 14660 400 14688 4519
rect 14936 400 14964 4519
rect 15198 4448 15254 4457
rect 15198 4383 15254 4392
rect 15212 400 15240 4383
rect 15488 400 15516 4519
rect 15750 1320 15806 1329
rect 15750 1255 15806 1264
rect 16026 1320 16082 1329
rect 16026 1255 16082 1264
rect 15764 400 15792 1255
rect 16040 400 16068 1255
rect 16316 400 16344 4519
rect 16592 400 16620 4519
rect 17682 4448 17738 4457
rect 17682 4383 17738 4392
rect 18786 4448 18842 4457
rect 18786 4383 18842 4392
rect 17222 4312 17278 4321
rect 17222 4247 17278 4256
rect 16854 2680 16910 2689
rect 16854 2615 16910 2624
rect 16868 400 16896 2615
rect 17130 2544 17186 2553
rect 17130 2479 17186 2488
rect 17144 400 17172 2479
rect 17236 898 17264 4247
rect 17306 2204 17614 2213
rect 17306 2202 17312 2204
rect 17368 2202 17392 2204
rect 17448 2202 17472 2204
rect 17528 2202 17552 2204
rect 17608 2202 17614 2204
rect 17368 2150 17370 2202
rect 17550 2150 17552 2202
rect 17306 2148 17312 2150
rect 17368 2148 17392 2150
rect 17448 2148 17472 2150
rect 17528 2148 17552 2150
rect 17608 2148 17614 2150
rect 17306 2139 17614 2148
rect 17306 1116 17614 1125
rect 17306 1114 17312 1116
rect 17368 1114 17392 1116
rect 17448 1114 17472 1116
rect 17528 1114 17552 1116
rect 17608 1114 17614 1116
rect 17368 1062 17370 1114
rect 17550 1062 17552 1114
rect 17306 1060 17312 1062
rect 17368 1060 17392 1062
rect 17448 1060 17472 1062
rect 17528 1060 17552 1062
rect 17608 1060 17614 1062
rect 17306 1051 17614 1060
rect 17236 870 17448 898
rect 17420 400 17448 870
rect 17696 400 17724 4383
rect 18326 4176 18382 4185
rect 18326 4111 18382 4120
rect 17946 1660 18254 1669
rect 17946 1658 17952 1660
rect 18008 1658 18032 1660
rect 18088 1658 18112 1660
rect 18168 1658 18192 1660
rect 18248 1658 18254 1660
rect 18008 1606 18010 1658
rect 18190 1606 18192 1658
rect 17946 1604 17952 1606
rect 18008 1604 18032 1606
rect 18088 1604 18112 1606
rect 18168 1604 18192 1606
rect 18248 1604 18254 1606
rect 17946 1595 18254 1604
rect 17866 912 17922 921
rect 17866 847 17922 856
rect 17880 456 17908 847
rect 17946 572 18254 581
rect 17946 570 17952 572
rect 18008 570 18032 572
rect 18088 570 18112 572
rect 18168 570 18192 572
rect 18248 570 18254 572
rect 18008 518 18010 570
rect 18190 518 18192 570
rect 17946 516 17952 518
rect 18008 516 18032 518
rect 18088 516 18112 518
rect 18168 516 18192 518
rect 18248 516 18254 518
rect 17946 507 18254 516
rect 18340 456 18368 4111
rect 18510 1320 18566 1329
rect 18510 1255 18566 1264
rect 17880 428 18000 456
rect 17972 400 18000 428
rect 18248 428 18368 456
rect 18248 400 18276 428
rect 18524 400 18552 1255
rect 18800 400 18828 4383
rect 19062 1184 19118 1193
rect 19062 1119 19118 1128
rect 19076 400 19104 1119
rect 19352 400 19380 4519
rect 20442 4448 20498 4457
rect 20442 4383 20498 4392
rect 20166 4176 20222 4185
rect 20166 4111 20222 4120
rect 19890 1048 19946 1057
rect 19890 983 19946 992
rect 19614 776 19670 785
rect 19614 711 19670 720
rect 19628 400 19656 711
rect 19904 400 19932 983
rect 20180 400 20208 4111
rect 20456 400 20484 4383
rect 22374 4312 22430 4321
rect 22374 4247 22430 4256
rect 20994 4176 21050 4185
rect 20994 4111 21050 4120
rect 20718 4040 20774 4049
rect 20718 3975 20774 3984
rect 20732 400 20760 3975
rect 21008 400 21036 4111
rect 21270 3496 21326 3505
rect 21270 3431 21326 3440
rect 21284 400 21312 3431
rect 21548 1352 21600 1358
rect 21548 1294 21600 1300
rect 21822 1320 21878 1329
rect 21560 400 21588 1294
rect 21822 1255 21878 1264
rect 21836 400 21864 1255
rect 22098 1048 22154 1057
rect 22098 983 22154 992
rect 22112 400 22140 983
rect 22388 400 22416 4247
rect 22558 2000 22614 2009
rect 22558 1935 22614 1944
rect 22572 1358 22600 1935
rect 22560 1352 22612 1358
rect 22560 1294 22612 1300
rect 22664 400 22692 4519
rect 24768 2916 24820 2922
rect 24768 2858 24820 2864
rect 24308 2440 24360 2446
rect 24308 2382 24360 2388
rect 23662 1864 23718 1873
rect 23662 1799 23718 1808
rect 23756 1828 23808 1834
rect 23572 1420 23624 1426
rect 23572 1362 23624 1368
rect 23480 1352 23532 1358
rect 22926 1320 22982 1329
rect 22926 1255 22982 1264
rect 23294 1320 23350 1329
rect 23480 1294 23532 1300
rect 23294 1255 23350 1264
rect 22940 400 22968 1255
rect 23204 876 23256 882
rect 23204 818 23256 824
rect 23216 400 23244 818
rect 23308 814 23336 1255
rect 23492 950 23520 1294
rect 23584 1018 23612 1362
rect 23572 1012 23624 1018
rect 23572 954 23624 960
rect 23480 944 23532 950
rect 23480 886 23532 892
rect 23296 808 23348 814
rect 23296 750 23348 756
rect 23492 400 23520 886
rect 23676 814 23704 1799
rect 23756 1770 23808 1776
rect 23768 1222 23796 1770
rect 23756 1216 23808 1222
rect 23756 1158 23808 1164
rect 23664 808 23716 814
rect 23664 750 23716 756
rect 23768 400 23796 1158
rect 24032 740 24084 746
rect 24032 682 24084 688
rect 24044 400 24072 682
rect 24320 400 24348 2382
rect 24584 1964 24636 1970
rect 24584 1906 24636 1912
rect 24596 400 24624 1906
rect 24780 746 24808 2858
rect 24860 2576 24912 2582
rect 24860 2518 24912 2524
rect 24768 740 24820 746
rect 24768 682 24820 688
rect 24872 626 24900 2518
rect 24964 882 24992 4519
rect 25226 4448 25282 4457
rect 25226 4383 25282 4392
rect 25778 4448 25834 4457
rect 25778 4383 25834 4392
rect 25136 2508 25188 2514
rect 25136 2450 25188 2456
rect 25044 1896 25096 1902
rect 25044 1838 25096 1844
rect 25056 1018 25084 1838
rect 25148 1562 25176 2450
rect 25136 1556 25188 1562
rect 25136 1498 25188 1504
rect 25240 1426 25268 4383
rect 25306 2204 25614 2213
rect 25306 2202 25312 2204
rect 25368 2202 25392 2204
rect 25448 2202 25472 2204
rect 25528 2202 25552 2204
rect 25608 2202 25614 2204
rect 25368 2150 25370 2202
rect 25550 2150 25552 2202
rect 25306 2148 25312 2150
rect 25368 2148 25392 2150
rect 25448 2148 25472 2150
rect 25528 2148 25552 2150
rect 25608 2148 25614 2150
rect 25306 2139 25614 2148
rect 25596 1896 25648 1902
rect 25596 1838 25648 1844
rect 25686 1864 25742 1873
rect 25228 1420 25280 1426
rect 25228 1362 25280 1368
rect 25226 1320 25282 1329
rect 25608 1306 25636 1838
rect 25686 1799 25742 1808
rect 25700 1426 25728 1799
rect 25792 1426 25820 4383
rect 25964 2848 26016 2854
rect 25964 2790 26016 2796
rect 25976 2038 26004 2790
rect 26056 2304 26108 2310
rect 26056 2246 26108 2252
rect 25964 2032 26016 2038
rect 25964 1974 26016 1980
rect 26068 1970 26096 2246
rect 26056 1964 26108 1970
rect 26056 1906 26108 1912
rect 26160 1850 26188 4519
rect 28262 4448 28318 4457
rect 28262 4383 28318 4392
rect 29920 4412 29972 4418
rect 27802 4040 27858 4049
rect 27802 3975 27858 3984
rect 26332 2916 26384 2922
rect 26332 2858 26384 2864
rect 25884 1822 26188 1850
rect 25688 1420 25740 1426
rect 25688 1362 25740 1368
rect 25780 1420 25832 1426
rect 25780 1362 25832 1368
rect 25608 1278 25728 1306
rect 25226 1255 25282 1264
rect 25044 1012 25096 1018
rect 25044 954 25096 960
rect 24952 876 25004 882
rect 24952 818 25004 824
rect 25240 814 25268 1255
rect 25306 1116 25614 1125
rect 25306 1114 25312 1116
rect 25368 1114 25392 1116
rect 25448 1114 25472 1116
rect 25528 1114 25552 1116
rect 25608 1114 25614 1116
rect 25368 1062 25370 1114
rect 25550 1062 25552 1114
rect 25306 1060 25312 1062
rect 25368 1060 25392 1062
rect 25448 1060 25472 1062
rect 25528 1060 25552 1062
rect 25608 1060 25614 1062
rect 25306 1051 25614 1060
rect 25700 1018 25728 1278
rect 25780 1284 25832 1290
rect 25780 1226 25832 1232
rect 25688 1012 25740 1018
rect 25688 954 25740 960
rect 25686 912 25742 921
rect 25686 847 25742 856
rect 25228 808 25280 814
rect 25228 750 25280 756
rect 24872 598 25452 626
rect 24872 462 24992 490
rect 24872 400 24900 462
rect 24964 406 24992 462
rect 25148 474 25268 490
rect 25148 468 25280 474
rect 25148 462 25228 468
rect 24952 400 25004 406
rect 25148 400 25176 462
rect 25228 410 25280 416
rect 25424 400 25452 598
rect 25700 400 25728 847
rect 25792 456 25820 1226
rect 25884 814 25912 1822
rect 25946 1660 26254 1669
rect 25946 1658 25952 1660
rect 26008 1658 26032 1660
rect 26088 1658 26112 1660
rect 26168 1658 26192 1660
rect 26248 1658 26254 1660
rect 26008 1606 26010 1658
rect 26190 1606 26192 1658
rect 25946 1604 25952 1606
rect 26008 1604 26032 1606
rect 26088 1604 26112 1606
rect 26168 1604 26192 1606
rect 26248 1604 26254 1606
rect 25946 1595 26254 1604
rect 25964 1352 26016 1358
rect 25964 1294 26016 1300
rect 25976 921 26004 1294
rect 25962 912 26018 921
rect 25962 847 26018 856
rect 25872 808 25924 814
rect 25872 750 25924 756
rect 25872 672 25924 678
rect 25872 614 25924 620
rect 25884 456 25912 614
rect 25946 572 26254 581
rect 25946 570 25952 572
rect 26008 570 26032 572
rect 26088 570 26112 572
rect 26168 570 26192 572
rect 26248 570 26254 572
rect 26008 518 26010 570
rect 26190 518 26192 570
rect 25946 516 25952 518
rect 26008 516 26032 518
rect 26088 516 26112 518
rect 26168 516 26192 518
rect 26248 516 26254 518
rect 25946 507 26254 516
rect 26344 456 26372 2858
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 26424 2032 26476 2038
rect 26424 1974 26476 1980
rect 26436 1494 26464 1974
rect 26792 1896 26844 1902
rect 26792 1838 26844 1844
rect 26804 1562 26832 1838
rect 26792 1556 26844 1562
rect 26792 1498 26844 1504
rect 26424 1488 26476 1494
rect 26896 1442 26924 2382
rect 27068 1760 27120 1766
rect 27068 1702 27120 1708
rect 26424 1430 26476 1436
rect 26804 1414 26924 1442
rect 26516 1284 26568 1290
rect 26516 1226 26568 1232
rect 25792 428 26004 456
rect 25976 400 26004 428
rect 26252 428 26372 456
rect 26252 400 26280 428
rect 26528 400 26556 1226
rect 26804 400 26832 1414
rect 27080 400 27108 1702
rect 27436 1420 27488 1426
rect 27436 1362 27488 1368
rect 27344 876 27396 882
rect 27344 818 27396 824
rect 27356 400 27384 818
rect 27448 406 27476 1362
rect 27436 400 27488 406
rect 27632 400 27660 2586
rect 27712 2508 27764 2514
rect 27712 2450 27764 2456
rect 27724 1018 27752 2450
rect 27712 1012 27764 1018
rect 27712 954 27764 960
rect 27816 814 27844 3975
rect 28080 3052 28132 3058
rect 28080 2994 28132 3000
rect 27988 2848 28040 2854
rect 27988 2790 28040 2796
rect 28000 2582 28028 2790
rect 27988 2576 28040 2582
rect 27988 2518 28040 2524
rect 27896 1828 27948 1834
rect 27896 1770 27948 1776
rect 27804 808 27856 814
rect 27804 750 27856 756
rect 27908 746 27936 1770
rect 28092 1442 28120 2994
rect 28172 2984 28224 2990
rect 28172 2926 28224 2932
rect 28184 2106 28212 2926
rect 28172 2100 28224 2106
rect 28172 2042 28224 2048
rect 28276 1902 28304 4383
rect 29920 4354 29972 4360
rect 28446 4176 28502 4185
rect 28446 4111 28502 4120
rect 28722 4176 28778 4185
rect 28722 4111 28778 4120
rect 28356 3868 28408 3874
rect 28356 3810 28408 3816
rect 28264 1896 28316 1902
rect 28264 1838 28316 1844
rect 27988 1420 28040 1426
rect 28092 1414 28212 1442
rect 27988 1362 28040 1368
rect 28000 1018 28028 1362
rect 28078 1320 28134 1329
rect 28078 1255 28134 1264
rect 27988 1012 28040 1018
rect 27988 954 28040 960
rect 28092 814 28120 1255
rect 28080 808 28132 814
rect 28080 750 28132 756
rect 27896 740 27948 746
rect 27896 682 27948 688
rect 27908 626 27936 682
rect 27816 598 27936 626
rect 27816 474 27844 598
rect 27908 474 28028 490
rect 27804 468 27856 474
rect 27804 410 27856 416
rect 27908 468 28040 474
rect 27908 462 27988 468
rect 27908 400 27936 462
rect 27988 410 28040 416
rect 28184 400 28212 1414
rect 28368 814 28396 3810
rect 28460 2990 28488 4111
rect 28736 2990 28764 4111
rect 29828 3460 29880 3466
rect 29828 3402 29880 3408
rect 29840 3058 29868 3402
rect 29828 3052 29880 3058
rect 29828 2994 29880 3000
rect 28448 2984 28500 2990
rect 28448 2926 28500 2932
rect 28724 2984 28776 2990
rect 28724 2926 28776 2932
rect 29092 2916 29144 2922
rect 29092 2858 29144 2864
rect 28538 2680 28594 2689
rect 28538 2615 28594 2624
rect 28448 2100 28500 2106
rect 28448 2042 28500 2048
rect 28356 808 28408 814
rect 28356 750 28408 756
rect 28460 400 28488 2042
rect 28552 1902 28580 2615
rect 29104 2514 29132 2858
rect 29828 2644 29880 2650
rect 29828 2586 29880 2592
rect 29000 2508 29052 2514
rect 29000 2450 29052 2456
rect 29092 2508 29144 2514
rect 29092 2450 29144 2456
rect 28724 1964 28776 1970
rect 28724 1906 28776 1912
rect 28540 1896 28592 1902
rect 28540 1838 28592 1844
rect 28632 1896 28684 1902
rect 28632 1838 28684 1844
rect 28644 474 28672 1838
rect 28632 468 28684 474
rect 28632 410 28684 416
rect 28736 400 28764 1906
rect 29012 950 29040 2450
rect 29092 2032 29144 2038
rect 29092 1974 29144 1980
rect 29000 944 29052 950
rect 29000 886 29052 892
rect 29104 762 29132 1974
rect 29276 1760 29328 1766
rect 29276 1702 29328 1708
rect 29288 1426 29316 1702
rect 29368 1488 29420 1494
rect 29368 1430 29420 1436
rect 29276 1420 29328 1426
rect 29276 1362 29328 1368
rect 29380 1306 29408 1430
rect 29012 734 29132 762
rect 29288 1278 29408 1306
rect 29012 400 29040 734
rect 29288 400 29316 1278
rect 29552 672 29604 678
rect 29552 614 29604 620
rect 29564 400 29592 614
rect 29840 400 29868 2586
rect 29932 1834 29960 4354
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 30380 3392 30432 3398
rect 30380 3334 30432 3340
rect 30392 2990 30420 3334
rect 30380 2984 30432 2990
rect 30380 2926 30432 2932
rect 30380 2848 30432 2854
rect 30380 2790 30432 2796
rect 30392 1902 30420 2790
rect 30484 2582 30512 3674
rect 30668 2990 30696 4519
rect 31022 4040 31078 4049
rect 31022 3975 31078 3984
rect 30656 2984 30708 2990
rect 30656 2926 30708 2932
rect 30564 2848 30616 2854
rect 30564 2790 30616 2796
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30576 2514 30604 2790
rect 31036 2514 31064 3975
rect 31300 3664 31352 3670
rect 31300 3606 31352 3612
rect 31116 3528 31168 3534
rect 31116 3470 31168 3476
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 31024 2508 31076 2514
rect 31024 2450 31076 2456
rect 30472 2440 30524 2446
rect 30472 2382 30524 2388
rect 30288 1896 30340 1902
rect 30288 1838 30340 1844
rect 30380 1896 30432 1902
rect 30380 1838 30432 1844
rect 29920 1828 29972 1834
rect 29920 1770 29972 1776
rect 30104 1556 30156 1562
rect 30104 1498 30156 1504
rect 30116 400 30144 1498
rect 30300 1018 30328 1838
rect 30378 1320 30434 1329
rect 30378 1255 30434 1264
rect 30288 1012 30340 1018
rect 30288 954 30340 960
rect 30392 814 30420 1255
rect 30380 808 30432 814
rect 30380 750 30432 756
rect 30484 660 30512 2382
rect 31024 2304 31076 2310
rect 31024 2246 31076 2252
rect 30840 1964 30892 1970
rect 30840 1906 30892 1912
rect 30852 1426 30880 1906
rect 31036 1426 31064 2246
rect 30840 1420 30892 1426
rect 30840 1362 30892 1368
rect 31024 1420 31076 1426
rect 31024 1362 31076 1368
rect 30748 1352 30800 1358
rect 30746 1320 30748 1329
rect 30800 1320 30802 1329
rect 30746 1255 30802 1264
rect 30930 1320 30986 1329
rect 30930 1255 30986 1264
rect 30654 1184 30710 1193
rect 30654 1119 30710 1128
rect 30668 814 30696 1119
rect 30840 944 30892 950
rect 30840 886 30892 892
rect 30656 808 30708 814
rect 30656 750 30708 756
rect 30852 660 30880 886
rect 30944 814 30972 1255
rect 30932 808 30984 814
rect 30932 750 30984 756
rect 30392 632 30512 660
rect 30668 632 30880 660
rect 30392 400 30420 632
rect 30668 400 30696 632
rect 31128 626 31156 3470
rect 31312 2854 31340 3606
rect 31484 2916 31536 2922
rect 31484 2858 31536 2864
rect 31300 2848 31352 2854
rect 31300 2790 31352 2796
rect 31312 2650 31340 2790
rect 31300 2644 31352 2650
rect 31300 2586 31352 2592
rect 31392 2644 31444 2650
rect 31392 2586 31444 2592
rect 31404 1834 31432 2586
rect 31496 2514 31524 2858
rect 31588 2582 31616 7806
rect 31680 7721 31708 7919
rect 31666 7712 31722 7721
rect 31666 7647 31722 7656
rect 31772 4978 31800 8486
rect 31852 8356 31904 8362
rect 31852 8298 31904 8304
rect 31680 4950 31800 4978
rect 31680 2990 31708 4950
rect 31864 3874 31892 8298
rect 31956 6361 31984 10950
rect 32048 10674 32076 11154
rect 32232 11150 32260 11494
rect 32220 11144 32272 11150
rect 32220 11086 32272 11092
rect 32220 10804 32272 10810
rect 32220 10746 32272 10752
rect 32036 10668 32088 10674
rect 32036 10610 32088 10616
rect 32128 10192 32180 10198
rect 32128 10134 32180 10140
rect 32140 9674 32168 10134
rect 32048 9646 32168 9674
rect 31942 6352 31998 6361
rect 31942 6287 31998 6296
rect 31944 5092 31996 5098
rect 31944 5034 31996 5040
rect 31852 3868 31904 3874
rect 31852 3810 31904 3816
rect 31668 2984 31720 2990
rect 31852 2984 31904 2990
rect 31668 2926 31720 2932
rect 31772 2944 31852 2972
rect 31576 2576 31628 2582
rect 31576 2518 31628 2524
rect 31484 2508 31536 2514
rect 31484 2450 31536 2456
rect 31668 2440 31720 2446
rect 31668 2382 31720 2388
rect 31484 2372 31536 2378
rect 31484 2314 31536 2320
rect 31392 1828 31444 1834
rect 31392 1770 31444 1776
rect 31208 1284 31260 1290
rect 31208 1226 31260 1232
rect 31220 1018 31248 1226
rect 31208 1012 31260 1018
rect 31208 954 31260 960
rect 30944 598 31156 626
rect 30944 400 30972 598
rect 31220 462 31340 490
rect 31220 400 31248 462
rect 31312 406 31340 462
rect 31300 400 31352 406
rect 31496 400 31524 2314
rect 31680 2038 31708 2382
rect 31668 2032 31720 2038
rect 31668 1974 31720 1980
rect 31772 400 31800 2944
rect 31852 2926 31904 2932
rect 31852 2304 31904 2310
rect 31852 2246 31904 2252
rect 31864 1902 31892 2246
rect 31956 1970 31984 5034
rect 32048 3942 32076 9646
rect 32128 5228 32180 5234
rect 32128 5170 32180 5176
rect 32036 3936 32088 3942
rect 32036 3878 32088 3884
rect 32036 3052 32088 3058
rect 32036 2994 32088 3000
rect 31944 1964 31996 1970
rect 31944 1906 31996 1912
rect 31852 1896 31904 1902
rect 31852 1838 31904 1844
rect 32048 1426 32076 2994
rect 32140 2446 32168 5170
rect 32232 4593 32260 10746
rect 32416 9926 32444 11600
rect 32732 11600 32734 11620
rect 32954 11600 33010 12000
rect 33230 11600 33286 12000
rect 33506 11600 33562 12000
rect 33782 11600 33838 12000
rect 34058 11600 34114 12000
rect 34334 11600 34390 12000
rect 34610 11600 34666 12000
rect 34886 11600 34942 12000
rect 35162 11600 35218 12000
rect 35438 11600 35494 12000
rect 35714 11600 35770 12000
rect 35990 11600 36046 12000
rect 36266 11600 36322 12000
rect 36542 11600 36598 12000
rect 36818 11600 36874 12000
rect 37094 11600 37150 12000
rect 37370 11600 37426 12000
rect 37646 11600 37702 12000
rect 37922 11600 37978 12000
rect 38198 11600 38254 12000
rect 38474 11600 38530 12000
rect 38750 11600 38806 12000
rect 32680 11562 32732 11568
rect 32588 11348 32640 11354
rect 32588 11290 32640 11296
rect 32772 11348 32824 11354
rect 32772 11290 32824 11296
rect 32600 11218 32628 11290
rect 32784 11218 32812 11290
rect 32588 11212 32640 11218
rect 32588 11154 32640 11160
rect 32772 11212 32824 11218
rect 32772 11154 32824 11160
rect 32864 11212 32916 11218
rect 32864 11154 32916 11160
rect 32600 11098 32628 11154
rect 32876 11098 32904 11154
rect 32600 11070 32904 11098
rect 32772 11008 32824 11014
rect 32772 10950 32824 10956
rect 32680 9988 32732 9994
rect 32680 9930 32732 9936
rect 32404 9920 32456 9926
rect 32310 9888 32366 9897
rect 32404 9862 32456 9868
rect 32310 9823 32366 9832
rect 32324 9674 32352 9823
rect 32324 9646 32444 9674
rect 32312 7336 32364 7342
rect 32312 7278 32364 7284
rect 32218 4584 32274 4593
rect 32218 4519 32274 4528
rect 32220 3120 32272 3126
rect 32220 3062 32272 3068
rect 32128 2440 32180 2446
rect 32128 2382 32180 2388
rect 32128 2304 32180 2310
rect 32128 2246 32180 2252
rect 32036 1420 32088 1426
rect 32036 1362 32088 1368
rect 32140 1306 32168 2246
rect 32048 1278 32168 1306
rect 32048 400 32076 1278
rect 32232 1018 32260 3062
rect 32220 1012 32272 1018
rect 32220 954 32272 960
rect 32324 400 32352 7278
rect 32416 3058 32444 9646
rect 32496 6792 32548 6798
rect 32496 6734 32548 6740
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32508 1442 32536 6734
rect 32588 5160 32640 5166
rect 32588 5102 32640 5108
rect 32600 2774 32628 5102
rect 32692 4078 32720 9930
rect 32784 4690 32812 10950
rect 32876 9722 32904 11070
rect 32968 10266 32996 11600
rect 33140 11008 33192 11014
rect 33140 10950 33192 10956
rect 33048 10532 33100 10538
rect 33048 10474 33100 10480
rect 32956 10260 33008 10266
rect 32956 10202 33008 10208
rect 32864 9716 32916 9722
rect 32864 9658 32916 9664
rect 32954 7848 33010 7857
rect 32954 7783 33010 7792
rect 32862 7712 32918 7721
rect 32862 7647 32918 7656
rect 32876 6866 32904 7647
rect 32864 6860 32916 6866
rect 32864 6802 32916 6808
rect 32864 6112 32916 6118
rect 32864 6054 32916 6060
rect 32772 4684 32824 4690
rect 32772 4626 32824 4632
rect 32876 4570 32904 6054
rect 32968 4690 32996 7783
rect 32956 4684 33008 4690
rect 32956 4626 33008 4632
rect 32784 4542 32904 4570
rect 32680 4072 32732 4078
rect 32680 4014 32732 4020
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 32692 3097 32720 3878
rect 32784 3618 32812 4542
rect 32956 4480 33008 4486
rect 32956 4422 33008 4428
rect 32864 4140 32916 4146
rect 32864 4082 32916 4088
rect 32876 3738 32904 4082
rect 32968 4026 32996 4422
rect 33060 4214 33088 10474
rect 33048 4208 33100 4214
rect 33152 4185 33180 10950
rect 33244 10810 33272 11600
rect 33520 11558 33548 11600
rect 33508 11552 33560 11558
rect 33508 11494 33560 11500
rect 33520 11150 33548 11494
rect 33796 11354 33824 11600
rect 34072 11540 34100 11600
rect 33888 11512 34100 11540
rect 33888 11354 33916 11512
rect 33946 11452 34254 11461
rect 33946 11450 33952 11452
rect 34008 11450 34032 11452
rect 34088 11450 34112 11452
rect 34168 11450 34192 11452
rect 34248 11450 34254 11452
rect 34008 11398 34010 11450
rect 34190 11398 34192 11450
rect 33946 11396 33952 11398
rect 34008 11396 34032 11398
rect 34088 11396 34112 11398
rect 34168 11396 34192 11398
rect 34248 11396 34254 11398
rect 33946 11387 34254 11396
rect 34348 11354 34376 11600
rect 33784 11348 33836 11354
rect 33784 11290 33836 11296
rect 33876 11348 33928 11354
rect 33876 11290 33928 11296
rect 34336 11348 34388 11354
rect 34336 11290 34388 11296
rect 33508 11144 33560 11150
rect 33508 11086 33560 11092
rect 33692 11076 33744 11082
rect 33692 11018 33744 11024
rect 33306 10908 33614 10917
rect 33306 10906 33312 10908
rect 33368 10906 33392 10908
rect 33448 10906 33472 10908
rect 33528 10906 33552 10908
rect 33608 10906 33614 10908
rect 33368 10854 33370 10906
rect 33550 10854 33552 10906
rect 33306 10852 33312 10854
rect 33368 10852 33392 10854
rect 33448 10852 33472 10854
rect 33528 10852 33552 10854
rect 33608 10852 33614 10854
rect 33306 10843 33614 10852
rect 33232 10804 33284 10810
rect 33232 10746 33284 10752
rect 33232 10464 33284 10470
rect 33232 10406 33284 10412
rect 33244 4842 33272 10406
rect 33306 9820 33614 9829
rect 33306 9818 33312 9820
rect 33368 9818 33392 9820
rect 33448 9818 33472 9820
rect 33528 9818 33552 9820
rect 33608 9818 33614 9820
rect 33368 9766 33370 9818
rect 33550 9766 33552 9818
rect 33306 9764 33312 9766
rect 33368 9764 33392 9766
rect 33448 9764 33472 9766
rect 33528 9764 33552 9766
rect 33608 9764 33614 9766
rect 33306 9755 33614 9764
rect 33324 9716 33376 9722
rect 33324 9658 33376 9664
rect 33336 7410 33364 9658
rect 33324 7404 33376 7410
rect 33324 7346 33376 7352
rect 33704 5114 33732 11018
rect 33784 11008 33836 11014
rect 33784 10950 33836 10956
rect 33612 5086 33732 5114
rect 33244 4814 33364 4842
rect 33232 4684 33284 4690
rect 33232 4626 33284 4632
rect 33048 4150 33100 4156
rect 33138 4176 33194 4185
rect 33138 4111 33194 4120
rect 33244 4026 33272 4626
rect 32968 3998 33088 4026
rect 32956 3936 33008 3942
rect 32956 3878 33008 3884
rect 32864 3732 32916 3738
rect 32864 3674 32916 3680
rect 32784 3590 32904 3618
rect 32968 3602 32996 3878
rect 32678 3088 32734 3097
rect 32678 3023 32734 3032
rect 32600 2746 32812 2774
rect 32784 2106 32812 2746
rect 32772 2100 32824 2106
rect 32772 2042 32824 2048
rect 32508 1414 32628 1442
rect 32600 400 32628 1414
rect 32784 1358 32812 2042
rect 32772 1352 32824 1358
rect 32772 1294 32824 1300
rect 32876 400 32904 3590
rect 32956 3596 33008 3602
rect 32956 3538 33008 3544
rect 32956 2848 33008 2854
rect 32956 2790 33008 2796
rect 32968 2582 32996 2790
rect 32956 2576 33008 2582
rect 32956 2518 33008 2524
rect 33060 1970 33088 3998
rect 33152 3998 33272 4026
rect 33048 1964 33100 1970
rect 33048 1906 33100 1912
rect 32954 1320 33010 1329
rect 32954 1255 33010 1264
rect 32968 814 32996 1255
rect 32956 808 33008 814
rect 32956 750 33008 756
rect 33152 400 33180 3998
rect 33230 3768 33286 3777
rect 33230 3703 33286 3712
rect 33244 3210 33272 3703
rect 33336 3398 33364 4814
rect 33416 4072 33468 4078
rect 33416 4014 33468 4020
rect 33508 4072 33560 4078
rect 33508 4014 33560 4020
rect 33428 3913 33456 4014
rect 33414 3904 33470 3913
rect 33414 3839 33470 3848
rect 33520 3618 33548 4014
rect 33428 3590 33548 3618
rect 33612 3602 33640 5086
rect 33692 5024 33744 5030
rect 33692 4966 33744 4972
rect 33600 3596 33652 3602
rect 33324 3392 33376 3398
rect 33324 3334 33376 3340
rect 33244 3182 33364 3210
rect 33230 3088 33286 3097
rect 33336 3058 33364 3182
rect 33230 3023 33286 3032
rect 33324 3052 33376 3058
rect 33244 2990 33272 3023
rect 33324 2994 33376 3000
rect 33232 2984 33284 2990
rect 33232 2926 33284 2932
rect 33428 2774 33456 3590
rect 33600 3538 33652 3544
rect 33598 3496 33654 3505
rect 33598 3431 33654 3440
rect 33244 2746 33456 2774
rect 33244 1000 33272 2746
rect 33612 2446 33640 3431
rect 33600 2440 33652 2446
rect 33600 2382 33652 2388
rect 33306 2204 33614 2213
rect 33306 2202 33312 2204
rect 33368 2202 33392 2204
rect 33448 2202 33472 2204
rect 33528 2202 33552 2204
rect 33608 2202 33614 2204
rect 33368 2150 33370 2202
rect 33550 2150 33552 2202
rect 33306 2148 33312 2150
rect 33368 2148 33392 2150
rect 33448 2148 33472 2150
rect 33528 2148 33552 2150
rect 33608 2148 33614 2150
rect 33306 2139 33614 2148
rect 33322 2000 33378 2009
rect 33322 1935 33324 1944
rect 33376 1935 33378 1944
rect 33324 1906 33376 1912
rect 33306 1116 33614 1125
rect 33306 1114 33312 1116
rect 33368 1114 33392 1116
rect 33448 1114 33472 1116
rect 33528 1114 33552 1116
rect 33608 1114 33614 1116
rect 33368 1062 33370 1114
rect 33550 1062 33552 1114
rect 33306 1060 33312 1062
rect 33368 1060 33392 1062
rect 33448 1060 33472 1062
rect 33528 1060 33552 1062
rect 33608 1060 33614 1062
rect 33306 1051 33614 1060
rect 33244 972 33456 1000
rect 33428 400 33456 972
rect 33704 814 33732 4966
rect 33796 4078 33824 10950
rect 33946 10364 34254 10373
rect 33946 10362 33952 10364
rect 34008 10362 34032 10364
rect 34088 10362 34112 10364
rect 34168 10362 34192 10364
rect 34248 10362 34254 10364
rect 34008 10310 34010 10362
rect 34190 10310 34192 10362
rect 33946 10308 33952 10310
rect 34008 10308 34032 10310
rect 34088 10308 34112 10310
rect 34168 10308 34192 10310
rect 34248 10308 34254 10310
rect 33946 10299 34254 10308
rect 33946 9276 34254 9285
rect 33946 9274 33952 9276
rect 34008 9274 34032 9276
rect 34088 9274 34112 9276
rect 34168 9274 34192 9276
rect 34248 9274 34254 9276
rect 34008 9222 34010 9274
rect 34190 9222 34192 9274
rect 33946 9220 33952 9222
rect 34008 9220 34032 9222
rect 34088 9220 34112 9222
rect 34168 9220 34192 9222
rect 34248 9220 34254 9222
rect 33946 9211 34254 9220
rect 33946 8188 34254 8197
rect 33946 8186 33952 8188
rect 34008 8186 34032 8188
rect 34088 8186 34112 8188
rect 34168 8186 34192 8188
rect 34248 8186 34254 8188
rect 34008 8134 34010 8186
rect 34190 8134 34192 8186
rect 33946 8132 33952 8134
rect 34008 8132 34032 8134
rect 34088 8132 34112 8134
rect 34168 8132 34192 8134
rect 34248 8132 34254 8134
rect 33946 8123 34254 8132
rect 33946 7100 34254 7109
rect 33946 7098 33952 7100
rect 34008 7098 34032 7100
rect 34088 7098 34112 7100
rect 34168 7098 34192 7100
rect 34248 7098 34254 7100
rect 34008 7046 34010 7098
rect 34190 7046 34192 7098
rect 33946 7044 33952 7046
rect 34008 7044 34032 7046
rect 34088 7044 34112 7046
rect 34168 7044 34192 7046
rect 34248 7044 34254 7046
rect 33946 7035 34254 7044
rect 34624 6866 34652 11600
rect 34612 6860 34664 6866
rect 34612 6802 34664 6808
rect 34900 6254 34928 11600
rect 34980 8084 35032 8090
rect 34980 8026 35032 8032
rect 34888 6248 34940 6254
rect 34888 6190 34940 6196
rect 33946 6012 34254 6021
rect 33946 6010 33952 6012
rect 34008 6010 34032 6012
rect 34088 6010 34112 6012
rect 34168 6010 34192 6012
rect 34248 6010 34254 6012
rect 34008 5958 34010 6010
rect 34190 5958 34192 6010
rect 33946 5956 33952 5958
rect 34008 5956 34032 5958
rect 34088 5956 34112 5958
rect 34168 5956 34192 5958
rect 34248 5956 34254 5958
rect 33946 5947 34254 5956
rect 33946 4924 34254 4933
rect 33946 4922 33952 4924
rect 34008 4922 34032 4924
rect 34088 4922 34112 4924
rect 34168 4922 34192 4924
rect 34248 4922 34254 4924
rect 34008 4870 34010 4922
rect 34190 4870 34192 4922
rect 33946 4868 33952 4870
rect 34008 4868 34032 4870
rect 34088 4868 34112 4870
rect 34168 4868 34192 4870
rect 34248 4868 34254 4870
rect 33946 4859 34254 4868
rect 34336 4480 34388 4486
rect 34336 4422 34388 4428
rect 34888 4480 34940 4486
rect 34888 4422 34940 4428
rect 33784 4072 33836 4078
rect 33784 4014 33836 4020
rect 33876 4004 33928 4010
rect 33876 3946 33928 3952
rect 33784 3460 33836 3466
rect 33784 3402 33836 3408
rect 33796 3194 33824 3402
rect 33784 3188 33836 3194
rect 33784 3130 33836 3136
rect 33888 2904 33916 3946
rect 33946 3836 34254 3845
rect 33946 3834 33952 3836
rect 34008 3834 34032 3836
rect 34088 3834 34112 3836
rect 34168 3834 34192 3836
rect 34248 3834 34254 3836
rect 34008 3782 34010 3834
rect 34190 3782 34192 3834
rect 33946 3780 33952 3782
rect 34008 3780 34032 3782
rect 34088 3780 34112 3782
rect 34168 3780 34192 3782
rect 34248 3780 34254 3782
rect 33946 3771 34254 3780
rect 34150 3632 34206 3641
rect 34060 3596 34112 3602
rect 34150 3567 34152 3576
rect 34060 3538 34112 3544
rect 34204 3567 34206 3576
rect 34152 3538 34204 3544
rect 34072 3398 34100 3538
rect 34348 3534 34376 4422
rect 34520 4208 34572 4214
rect 34520 4150 34572 4156
rect 34428 4072 34480 4078
rect 34428 4014 34480 4020
rect 34336 3528 34388 3534
rect 34336 3470 34388 3476
rect 34060 3392 34112 3398
rect 34060 3334 34112 3340
rect 33968 3120 34020 3126
rect 33968 3062 34020 3068
rect 33796 2876 33916 2904
rect 33796 1834 33824 2876
rect 33980 2836 34008 3062
rect 33888 2808 34008 2836
rect 34336 2848 34388 2854
rect 33784 1828 33836 1834
rect 33784 1770 33836 1776
rect 33782 1728 33838 1737
rect 33782 1663 33838 1672
rect 33796 882 33824 1663
rect 33784 876 33836 882
rect 33784 818 33836 824
rect 33692 808 33744 814
rect 33888 796 33916 2808
rect 34336 2790 34388 2796
rect 33946 2748 34254 2757
rect 33946 2746 33952 2748
rect 34008 2746 34032 2748
rect 34088 2746 34112 2748
rect 34168 2746 34192 2748
rect 34248 2746 34254 2748
rect 34008 2694 34010 2746
rect 34190 2694 34192 2746
rect 33946 2692 33952 2694
rect 34008 2692 34032 2694
rect 34088 2692 34112 2694
rect 34168 2692 34192 2694
rect 34248 2692 34254 2694
rect 33946 2683 34254 2692
rect 33968 1896 34020 1902
rect 33966 1864 33968 1873
rect 34020 1864 34022 1873
rect 33966 1799 34022 1808
rect 33946 1660 34254 1669
rect 33946 1658 33952 1660
rect 34008 1658 34032 1660
rect 34088 1658 34112 1660
rect 34168 1658 34192 1660
rect 34248 1658 34254 1660
rect 34008 1606 34010 1658
rect 34190 1606 34192 1658
rect 33946 1604 33952 1606
rect 34008 1604 34032 1606
rect 34088 1604 34112 1606
rect 34168 1604 34192 1606
rect 34248 1604 34254 1606
rect 33946 1595 34254 1604
rect 34060 1556 34112 1562
rect 34060 1498 34112 1504
rect 34072 1358 34100 1498
rect 34348 1442 34376 2790
rect 34440 1970 34468 4014
rect 34532 2650 34560 4150
rect 34796 4004 34848 4010
rect 34796 3946 34848 3952
rect 34612 3936 34664 3942
rect 34612 3878 34664 3884
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 34624 3534 34652 3878
rect 34716 3670 34744 3878
rect 34704 3664 34756 3670
rect 34704 3606 34756 3612
rect 34808 3602 34836 3946
rect 34796 3596 34848 3602
rect 34796 3538 34848 3544
rect 34612 3528 34664 3534
rect 34900 3482 34928 4422
rect 34612 3470 34664 3476
rect 34716 3454 34928 3482
rect 34612 3392 34664 3398
rect 34612 3334 34664 3340
rect 34624 2990 34652 3334
rect 34612 2984 34664 2990
rect 34612 2926 34664 2932
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 34716 2514 34744 3454
rect 34888 3052 34940 3058
rect 34888 2994 34940 3000
rect 34900 2961 34928 2994
rect 34992 2990 35020 8026
rect 35070 7304 35126 7313
rect 35070 7239 35126 7248
rect 35084 3097 35112 7239
rect 35176 4690 35204 11600
rect 35256 7880 35308 7886
rect 35256 7822 35308 7828
rect 35164 4684 35216 4690
rect 35164 4626 35216 4632
rect 35164 3936 35216 3942
rect 35164 3878 35216 3884
rect 35176 3505 35204 3878
rect 35162 3496 35218 3505
rect 35268 3466 35296 7822
rect 35452 6338 35480 11600
rect 35728 9738 35756 11600
rect 35728 9710 35940 9738
rect 35624 6792 35676 6798
rect 35624 6734 35676 6740
rect 35360 6310 35480 6338
rect 35360 4146 35388 6310
rect 35636 6254 35664 6734
rect 35624 6248 35676 6254
rect 35624 6190 35676 6196
rect 35912 4978 35940 9710
rect 36004 6440 36032 11600
rect 36084 8016 36136 8022
rect 36084 7958 36136 7964
rect 36096 6934 36124 7958
rect 36176 7744 36228 7750
rect 36176 7686 36228 7692
rect 36084 6928 36136 6934
rect 36084 6870 36136 6876
rect 36004 6412 36124 6440
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 36004 5166 36032 6258
rect 35992 5160 36044 5166
rect 35992 5102 36044 5108
rect 35912 4950 36032 4978
rect 35900 4616 35952 4622
rect 35900 4558 35952 4564
rect 35624 4480 35676 4486
rect 35624 4422 35676 4428
rect 35348 4140 35400 4146
rect 35348 4082 35400 4088
rect 35360 3602 35388 4082
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 35452 3602 35480 3878
rect 35348 3596 35400 3602
rect 35348 3538 35400 3544
rect 35440 3596 35492 3602
rect 35440 3538 35492 3544
rect 35162 3431 35218 3440
rect 35256 3460 35308 3466
rect 35256 3402 35308 3408
rect 35070 3088 35126 3097
rect 35070 3023 35126 3032
rect 34980 2984 35032 2990
rect 34886 2952 34942 2961
rect 34980 2926 35032 2932
rect 34886 2887 34942 2896
rect 35072 2916 35124 2922
rect 35072 2858 35124 2864
rect 34704 2508 34756 2514
rect 34704 2450 34756 2456
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34612 2372 34664 2378
rect 34612 2314 34664 2320
rect 34520 2100 34572 2106
rect 34520 2042 34572 2048
rect 34428 1964 34480 1970
rect 34428 1906 34480 1912
rect 34256 1426 34376 1442
rect 34244 1420 34376 1426
rect 34296 1414 34376 1420
rect 34244 1362 34296 1368
rect 34060 1352 34112 1358
rect 34060 1294 34112 1300
rect 34336 1352 34388 1358
rect 34336 1294 34388 1300
rect 33968 808 34020 814
rect 33888 768 33968 796
rect 33692 750 33744 756
rect 33968 750 34020 756
rect 33704 400 33732 750
rect 33946 572 34254 581
rect 33946 570 33952 572
rect 34008 570 34032 572
rect 34088 570 34112 572
rect 34168 570 34192 572
rect 34248 570 34254 572
rect 34008 518 34010 570
rect 34190 518 34192 570
rect 33946 516 33952 518
rect 34008 516 34032 518
rect 34088 516 34112 518
rect 34168 516 34192 518
rect 34248 516 34254 518
rect 33946 507 34254 516
rect 33876 468 33928 474
rect 34348 456 34376 1294
rect 34440 474 34468 1906
rect 33928 428 34008 456
rect 33876 410 33928 416
rect 33980 400 34008 428
rect 34256 428 34376 456
rect 34428 468 34480 474
rect 34256 400 34284 428
rect 34428 410 34480 416
rect 34532 400 34560 2042
rect 34624 1970 34652 2314
rect 34612 1964 34664 1970
rect 34612 1906 34664 1912
rect 34624 950 34652 1906
rect 34612 944 34664 950
rect 34612 886 34664 892
rect 34808 400 34836 2382
rect 35084 400 35112 2858
rect 35452 2774 35480 3538
rect 35532 3528 35584 3534
rect 35532 3470 35584 3476
rect 35360 2746 35480 2774
rect 35164 2304 35216 2310
rect 35164 2246 35216 2252
rect 35176 2038 35204 2246
rect 35164 2032 35216 2038
rect 35164 1974 35216 1980
rect 35256 740 35308 746
rect 35256 682 35308 688
rect 2778 0 2834 400
rect 3054 0 3110 400
rect 3330 0 3386 400
rect 3606 0 3662 400
rect 3882 0 3938 400
rect 4158 0 4214 400
rect 4434 0 4490 400
rect 4710 0 4766 400
rect 4986 0 5042 400
rect 5262 0 5318 400
rect 5538 0 5594 400
rect 5814 0 5870 400
rect 6090 0 6146 400
rect 6366 0 6422 400
rect 6642 0 6698 400
rect 6918 0 6974 400
rect 7194 0 7250 400
rect 7470 0 7526 400
rect 7746 0 7802 400
rect 8022 0 8078 400
rect 8298 0 8354 400
rect 8574 0 8630 400
rect 8850 0 8906 400
rect 9126 0 9182 400
rect 9402 0 9458 400
rect 9678 0 9734 400
rect 9954 0 10010 400
rect 10230 0 10286 400
rect 10506 0 10562 400
rect 10782 0 10838 400
rect 11058 0 11114 400
rect 11334 0 11390 400
rect 11610 0 11666 400
rect 11886 0 11942 400
rect 12162 0 12218 400
rect 12438 0 12494 400
rect 12714 0 12770 400
rect 12990 0 13046 400
rect 13266 0 13322 400
rect 13542 0 13598 400
rect 13818 0 13874 400
rect 14094 0 14150 400
rect 14370 0 14426 400
rect 14646 0 14702 400
rect 14922 0 14978 400
rect 15198 0 15254 400
rect 15474 0 15530 400
rect 15750 0 15806 400
rect 16026 0 16082 400
rect 16302 0 16358 400
rect 16578 0 16634 400
rect 16854 0 16910 400
rect 17130 0 17186 400
rect 17406 0 17462 400
rect 17682 0 17738 400
rect 17958 0 18014 400
rect 18234 0 18290 400
rect 18510 0 18566 400
rect 18786 0 18842 400
rect 19062 0 19118 400
rect 19338 0 19394 400
rect 19614 0 19670 400
rect 19890 0 19946 400
rect 20166 0 20222 400
rect 20442 0 20498 400
rect 20718 0 20774 400
rect 20994 0 21050 400
rect 21270 0 21326 400
rect 21546 0 21602 400
rect 21822 0 21878 400
rect 22098 0 22154 400
rect 22374 0 22430 400
rect 22650 0 22706 400
rect 22926 0 22982 400
rect 23202 0 23258 400
rect 23478 0 23534 400
rect 23754 0 23810 400
rect 24030 0 24086 400
rect 24306 0 24362 400
rect 24582 0 24638 400
rect 24858 0 24914 400
rect 24952 342 25004 348
rect 25134 0 25190 400
rect 25410 0 25466 400
rect 25686 0 25742 400
rect 25962 0 26018 400
rect 26238 0 26294 400
rect 26514 0 26570 400
rect 26790 0 26846 400
rect 27066 0 27122 400
rect 27342 0 27398 400
rect 27436 342 27488 348
rect 27618 0 27674 400
rect 27894 0 27950 400
rect 28170 0 28226 400
rect 28446 0 28502 400
rect 28722 0 28778 400
rect 28998 0 29054 400
rect 29274 0 29330 400
rect 29550 0 29606 400
rect 29826 0 29882 400
rect 30102 0 30158 400
rect 30378 0 30434 400
rect 30654 0 30710 400
rect 30930 0 30986 400
rect 31206 0 31262 400
rect 31300 342 31352 348
rect 31482 0 31538 400
rect 31758 0 31814 400
rect 32034 0 32090 400
rect 32310 0 32366 400
rect 32586 0 32642 400
rect 32862 0 32918 400
rect 33138 0 33194 400
rect 33414 0 33470 400
rect 33690 0 33746 400
rect 33966 0 34022 400
rect 34242 0 34298 400
rect 34518 0 34574 400
rect 34794 0 34850 400
rect 35070 0 35126 400
rect 35268 338 35296 682
rect 35360 400 35388 2746
rect 35544 1902 35572 3470
rect 35636 2990 35664 4422
rect 35912 4078 35940 4558
rect 35900 4072 35952 4078
rect 35900 4014 35952 4020
rect 35808 4004 35860 4010
rect 35808 3946 35860 3952
rect 35820 3602 35848 3946
rect 35900 3936 35952 3942
rect 35900 3878 35952 3884
rect 35808 3596 35860 3602
rect 35808 3538 35860 3544
rect 35820 3482 35848 3538
rect 35728 3454 35848 3482
rect 35624 2984 35676 2990
rect 35624 2926 35676 2932
rect 35728 2774 35756 3454
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 35820 2990 35848 3334
rect 35808 2984 35860 2990
rect 35808 2926 35860 2932
rect 35636 2746 35756 2774
rect 35532 1896 35584 1902
rect 35532 1838 35584 1844
rect 35636 400 35664 2746
rect 35912 2514 35940 3878
rect 35900 2508 35952 2514
rect 35900 2450 35952 2456
rect 35716 1896 35768 1902
rect 35716 1838 35768 1844
rect 35728 1290 35756 1838
rect 35716 1284 35768 1290
rect 35716 1226 35768 1232
rect 36004 814 36032 4950
rect 36096 4282 36124 6412
rect 36084 4276 36136 4282
rect 36084 4218 36136 4224
rect 36188 3890 36216 7686
rect 36096 3862 36216 3890
rect 36096 3534 36124 3862
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 36176 3460 36228 3466
rect 36176 3402 36228 3408
rect 36084 3120 36136 3126
rect 36084 3062 36136 3068
rect 35992 808 36044 814
rect 35992 750 36044 756
rect 36096 660 36124 3062
rect 35912 632 36124 660
rect 35912 400 35940 632
rect 36188 400 36216 3402
rect 36280 2825 36308 11600
rect 36452 7812 36504 7818
rect 36452 7754 36504 7760
rect 36360 7540 36412 7546
rect 36360 7482 36412 7488
rect 36372 3942 36400 7482
rect 36464 7018 36492 7754
rect 36556 7154 36584 11600
rect 36556 7126 36676 7154
rect 36464 6990 36584 7018
rect 36452 6928 36504 6934
rect 36452 6870 36504 6876
rect 36360 3936 36412 3942
rect 36360 3878 36412 3884
rect 36464 3754 36492 6870
rect 36372 3726 36492 3754
rect 36372 3194 36400 3726
rect 36452 3664 36504 3670
rect 36452 3606 36504 3612
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 36360 3052 36412 3058
rect 36360 2994 36412 3000
rect 36266 2816 36322 2825
rect 36266 2751 36322 2760
rect 36266 2544 36322 2553
rect 36266 2479 36322 2488
rect 36280 1358 36308 2479
rect 36372 1494 36400 2994
rect 36360 1488 36412 1494
rect 36360 1430 36412 1436
rect 36268 1352 36320 1358
rect 36268 1294 36320 1300
rect 36360 1216 36412 1222
rect 36360 1158 36412 1164
rect 36372 1018 36400 1158
rect 36360 1012 36412 1018
rect 36360 954 36412 960
rect 36266 912 36322 921
rect 36266 847 36322 856
rect 36280 814 36308 847
rect 36464 814 36492 3606
rect 36556 3602 36584 6990
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 36544 3188 36596 3194
rect 36544 3130 36596 3136
rect 36556 2582 36584 3130
rect 36544 2576 36596 2582
rect 36544 2518 36596 2524
rect 36542 2136 36598 2145
rect 36542 2071 36598 2080
rect 36268 808 36320 814
rect 36268 750 36320 756
rect 36452 808 36504 814
rect 36452 750 36504 756
rect 36556 660 36584 2071
rect 36648 1970 36676 7126
rect 36728 3936 36780 3942
rect 36728 3878 36780 3884
rect 36740 3466 36768 3878
rect 36728 3460 36780 3466
rect 36728 3402 36780 3408
rect 36832 3369 36860 11600
rect 37004 6112 37056 6118
rect 37004 6054 37056 6060
rect 36912 4276 36964 4282
rect 36912 4218 36964 4224
rect 36818 3360 36874 3369
rect 36818 3295 36874 3304
rect 36924 2904 36952 4218
rect 36740 2876 36952 2904
rect 36740 2258 36768 2876
rect 36910 2816 36966 2825
rect 36910 2751 36966 2760
rect 36818 2680 36874 2689
rect 36818 2615 36874 2624
rect 36832 2378 36860 2615
rect 36820 2372 36872 2378
rect 36820 2314 36872 2320
rect 36740 2230 36860 2258
rect 36728 2100 36780 2106
rect 36728 2042 36780 2048
rect 36636 1964 36688 1970
rect 36636 1906 36688 1912
rect 36634 1864 36690 1873
rect 36634 1799 36690 1808
rect 36648 1426 36676 1799
rect 36740 1494 36768 2042
rect 36728 1488 36780 1494
rect 36728 1430 36780 1436
rect 36832 1426 36860 2230
rect 36924 1494 36952 2751
rect 36912 1488 36964 1494
rect 36912 1430 36964 1436
rect 36636 1420 36688 1426
rect 36636 1362 36688 1368
rect 36820 1420 36872 1426
rect 36820 1362 36872 1368
rect 36728 1216 36780 1222
rect 36728 1158 36780 1164
rect 36820 1216 36872 1222
rect 36820 1158 36872 1164
rect 36740 950 36768 1158
rect 36728 944 36780 950
rect 36728 886 36780 892
rect 36832 762 36860 1158
rect 36464 632 36584 660
rect 36740 734 36860 762
rect 36464 400 36492 632
rect 36740 400 36768 734
rect 37016 400 37044 6054
rect 37108 3738 37136 11600
rect 37280 5024 37332 5030
rect 37280 4966 37332 4972
rect 37096 3732 37148 3738
rect 37096 3674 37148 3680
rect 37108 2972 37136 3674
rect 37292 3482 37320 4966
rect 37384 3602 37412 11600
rect 37660 7206 37688 11600
rect 37648 7200 37700 7206
rect 37648 7142 37700 7148
rect 37936 6458 37964 11600
rect 37924 6452 37976 6458
rect 37924 6394 37976 6400
rect 37924 4140 37976 4146
rect 37924 4082 37976 4088
rect 37740 4004 37792 4010
rect 37740 3946 37792 3952
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 37648 3528 37700 3534
rect 37188 3460 37240 3466
rect 37292 3454 37412 3482
rect 37648 3470 37700 3476
rect 37188 3402 37240 3408
rect 37200 3126 37228 3402
rect 37278 3360 37334 3369
rect 37278 3295 37334 3304
rect 37188 3120 37240 3126
rect 37188 3062 37240 3068
rect 37188 2984 37240 2990
rect 37108 2944 37188 2972
rect 37188 2926 37240 2932
rect 37292 2514 37320 3295
rect 37280 2508 37332 2514
rect 37280 2450 37332 2456
rect 37384 898 37412 3454
rect 37464 3392 37516 3398
rect 37516 3352 37596 3380
rect 37464 3334 37516 3340
rect 37462 3088 37518 3097
rect 37462 3023 37464 3032
rect 37516 3023 37518 3032
rect 37464 2994 37516 3000
rect 37568 2802 37596 3352
rect 37476 2774 37596 2802
rect 37476 2514 37504 2774
rect 37464 2508 37516 2514
rect 37464 2450 37516 2456
rect 37556 2508 37608 2514
rect 37556 2450 37608 2456
rect 37568 2417 37596 2450
rect 37554 2408 37610 2417
rect 37554 2343 37610 2352
rect 37554 2272 37610 2281
rect 37554 2207 37610 2216
rect 37568 1834 37596 2207
rect 37556 1828 37608 1834
rect 37556 1770 37608 1776
rect 37556 1420 37608 1426
rect 37556 1362 37608 1368
rect 37292 870 37412 898
rect 37292 400 37320 870
rect 37464 740 37516 746
rect 37464 682 37516 688
rect 37476 406 37504 682
rect 37464 400 37516 406
rect 37568 400 37596 1362
rect 37660 814 37688 3470
rect 37752 2854 37780 3946
rect 37832 3664 37884 3670
rect 37832 3606 37884 3612
rect 37740 2848 37792 2854
rect 37740 2790 37792 2796
rect 37752 1442 37780 2790
rect 37844 1902 37872 3606
rect 37832 1896 37884 1902
rect 37832 1838 37884 1844
rect 37752 1414 37872 1442
rect 37936 1426 37964 4082
rect 38014 3360 38070 3369
rect 38014 3295 38070 3304
rect 38028 3126 38056 3295
rect 38016 3120 38068 3126
rect 38016 3062 38068 3068
rect 38212 3074 38240 11600
rect 38384 7200 38436 7206
rect 38384 7142 38436 7148
rect 38212 3046 38332 3074
rect 38108 2984 38160 2990
rect 38014 2952 38070 2961
rect 38108 2926 38160 2932
rect 38014 2887 38070 2896
rect 38028 2854 38056 2887
rect 38016 2848 38068 2854
rect 38016 2790 38068 2796
rect 38120 2689 38148 2926
rect 38200 2916 38252 2922
rect 38200 2858 38252 2864
rect 38106 2680 38162 2689
rect 38106 2615 38162 2624
rect 38106 2544 38162 2553
rect 38106 2479 38108 2488
rect 38160 2479 38162 2488
rect 38108 2450 38160 2456
rect 38212 1426 38240 2858
rect 38304 2825 38332 3046
rect 38290 2816 38346 2825
rect 38290 2751 38346 2760
rect 38290 2680 38346 2689
rect 38290 2615 38346 2624
rect 37648 808 37700 814
rect 37648 750 37700 756
rect 37844 400 37872 1414
rect 37924 1420 37976 1426
rect 37924 1362 37976 1368
rect 38200 1420 38252 1426
rect 38200 1362 38252 1368
rect 38304 898 38332 2615
rect 38396 1902 38424 7142
rect 38488 2689 38516 11600
rect 38764 9722 38792 11600
rect 41946 11452 42254 11461
rect 41946 11450 41952 11452
rect 42008 11450 42032 11452
rect 42088 11450 42112 11452
rect 42168 11450 42192 11452
rect 42248 11450 42254 11452
rect 42008 11398 42010 11450
rect 42190 11398 42192 11450
rect 41946 11396 41952 11398
rect 42008 11396 42032 11398
rect 42088 11396 42112 11398
rect 42168 11396 42192 11398
rect 42248 11396 42254 11398
rect 41946 11387 42254 11396
rect 41306 10908 41614 10917
rect 41306 10906 41312 10908
rect 41368 10906 41392 10908
rect 41448 10906 41472 10908
rect 41528 10906 41552 10908
rect 41608 10906 41614 10908
rect 41368 10854 41370 10906
rect 41550 10854 41552 10906
rect 41306 10852 41312 10854
rect 41368 10852 41392 10854
rect 41448 10852 41472 10854
rect 41528 10852 41552 10854
rect 41608 10852 41614 10854
rect 41306 10843 41614 10852
rect 41946 10364 42254 10373
rect 41946 10362 41952 10364
rect 42008 10362 42032 10364
rect 42088 10362 42112 10364
rect 42168 10362 42192 10364
rect 42248 10362 42254 10364
rect 42008 10310 42010 10362
rect 42190 10310 42192 10362
rect 41946 10308 41952 10310
rect 42008 10308 42032 10310
rect 42088 10308 42112 10310
rect 42168 10308 42192 10310
rect 42248 10308 42254 10310
rect 41946 10299 42254 10308
rect 41306 9820 41614 9829
rect 41306 9818 41312 9820
rect 41368 9818 41392 9820
rect 41448 9818 41472 9820
rect 41528 9818 41552 9820
rect 41608 9818 41614 9820
rect 41368 9766 41370 9818
rect 41550 9766 41552 9818
rect 41306 9764 41312 9766
rect 41368 9764 41392 9766
rect 41448 9764 41472 9766
rect 41528 9764 41552 9766
rect 41608 9764 41614 9766
rect 41306 9755 41614 9764
rect 38752 9716 38804 9722
rect 38752 9658 38804 9664
rect 40500 9716 40552 9722
rect 40500 9658 40552 9664
rect 39856 6452 39908 6458
rect 39856 6394 39908 6400
rect 38568 3596 38620 3602
rect 38568 3538 38620 3544
rect 38474 2680 38530 2689
rect 38474 2615 38530 2624
rect 38580 2553 38608 3538
rect 39028 3188 39080 3194
rect 39028 3130 39080 3136
rect 38844 2848 38896 2854
rect 38844 2790 38896 2796
rect 38856 2582 38884 2790
rect 38844 2576 38896 2582
rect 38566 2544 38622 2553
rect 38476 2508 38528 2514
rect 38566 2479 38622 2488
rect 38750 2544 38806 2553
rect 38844 2518 38896 2524
rect 39040 2530 39068 3130
rect 39118 2952 39174 2961
rect 39118 2887 39174 2896
rect 39132 2650 39160 2887
rect 39120 2644 39172 2650
rect 39120 2586 39172 2592
rect 38750 2479 38806 2488
rect 38476 2450 38528 2456
rect 38488 2038 38516 2450
rect 38568 2440 38620 2446
rect 38568 2382 38620 2388
rect 38476 2032 38528 2038
rect 38476 1974 38528 1980
rect 38384 1896 38436 1902
rect 38384 1838 38436 1844
rect 38580 1766 38608 2382
rect 38660 2372 38712 2378
rect 38764 2360 38792 2479
rect 38712 2332 38792 2360
rect 38660 2314 38712 2320
rect 38856 2258 38884 2518
rect 39040 2502 39344 2530
rect 39120 2440 39172 2446
rect 39120 2382 39172 2388
rect 38856 2230 39068 2258
rect 39040 2145 39068 2230
rect 39026 2136 39082 2145
rect 39026 2071 39082 2080
rect 38752 2032 38804 2038
rect 38750 2000 38752 2009
rect 38804 2000 38806 2009
rect 38750 1935 38806 1944
rect 38660 1896 38712 1902
rect 38658 1864 38660 1873
rect 38712 1864 38714 1873
rect 38658 1799 38714 1808
rect 38934 1864 38990 1873
rect 38934 1799 38990 1808
rect 38568 1760 38620 1766
rect 38568 1702 38620 1708
rect 38752 1760 38804 1766
rect 38752 1702 38804 1708
rect 38764 1601 38792 1702
rect 38750 1592 38806 1601
rect 38750 1527 38806 1536
rect 38660 1352 38712 1358
rect 38660 1294 38712 1300
rect 38672 1018 38700 1294
rect 38660 1012 38712 1018
rect 38660 954 38712 960
rect 38304 870 38608 898
rect 38120 474 38240 490
rect 38120 468 38252 474
rect 38120 462 38200 468
rect 38120 400 38148 462
rect 38200 410 38252 416
rect 35256 332 35308 338
rect 35256 274 35308 280
rect 35346 0 35402 400
rect 35622 0 35678 400
rect 35898 0 35954 400
rect 36174 0 36230 400
rect 36450 0 36506 400
rect 36726 0 36782 400
rect 37002 0 37058 400
rect 37278 0 37334 400
rect 37464 342 37516 348
rect 37554 0 37610 400
rect 37830 0 37886 400
rect 38106 0 38162 400
rect 38304 202 38332 870
rect 38580 814 38608 870
rect 38948 814 38976 1799
rect 39132 1426 39160 2382
rect 39212 2304 39264 2310
rect 39212 2246 39264 2252
rect 39224 2009 39252 2246
rect 39210 2000 39266 2009
rect 39210 1935 39266 1944
rect 39316 1902 39344 2502
rect 39394 2408 39450 2417
rect 39394 2343 39450 2352
rect 39580 2372 39632 2378
rect 39408 1902 39436 2343
rect 39580 2314 39632 2320
rect 39592 2106 39620 2314
rect 39672 2304 39724 2310
rect 39670 2272 39672 2281
rect 39764 2304 39816 2310
rect 39724 2272 39726 2281
rect 39764 2246 39816 2252
rect 39670 2207 39726 2216
rect 39580 2100 39632 2106
rect 39580 2042 39632 2048
rect 39488 2032 39540 2038
rect 39488 1974 39540 1980
rect 39304 1896 39356 1902
rect 39304 1838 39356 1844
rect 39396 1896 39448 1902
rect 39396 1838 39448 1844
rect 39212 1760 39264 1766
rect 39212 1702 39264 1708
rect 39224 1562 39252 1702
rect 39302 1592 39358 1601
rect 39212 1556 39264 1562
rect 39302 1527 39358 1536
rect 39212 1498 39264 1504
rect 39120 1420 39172 1426
rect 39120 1362 39172 1368
rect 39316 1306 39344 1527
rect 39224 1278 39344 1306
rect 38568 808 38620 814
rect 38936 808 38988 814
rect 38568 750 38620 756
rect 38658 776 38714 785
rect 38936 750 38988 756
rect 38658 711 38714 720
rect 38396 462 38516 490
rect 38396 400 38424 462
rect 38292 196 38344 202
rect 38292 138 38344 144
rect 38382 0 38438 400
rect 38488 354 38516 462
rect 38672 400 38700 711
rect 39028 672 39080 678
rect 38856 632 39028 660
rect 38856 474 38884 632
rect 39028 614 39080 620
rect 38844 468 38896 474
rect 38844 410 38896 416
rect 38948 462 39068 490
rect 38948 400 38976 462
rect 39040 406 39068 462
rect 39028 400 39080 406
rect 39224 400 39252 1278
rect 39304 1216 39356 1222
rect 39304 1158 39356 1164
rect 39316 814 39344 1158
rect 39304 808 39356 814
rect 39304 750 39356 756
rect 38488 326 38608 354
rect 38580 66 38608 326
rect 38568 60 38620 66
rect 38568 2 38620 8
rect 38658 0 38714 400
rect 38934 0 38990 400
rect 39028 342 39080 348
rect 39210 0 39266 400
rect 39316 134 39344 750
rect 39500 400 39528 1974
rect 39592 1306 39620 2042
rect 39776 2038 39804 2246
rect 39764 2032 39816 2038
rect 39764 1974 39816 1980
rect 39868 1834 39896 6394
rect 40038 2680 40094 2689
rect 40038 2615 40094 2624
rect 39856 1828 39908 1834
rect 39856 1770 39908 1776
rect 39764 1488 39816 1494
rect 39868 1476 39896 1770
rect 40052 1562 40080 2615
rect 40512 2310 40540 9658
rect 41946 9276 42254 9285
rect 41946 9274 41952 9276
rect 42008 9274 42032 9276
rect 42088 9274 42112 9276
rect 42168 9274 42192 9276
rect 42248 9274 42254 9276
rect 42008 9222 42010 9274
rect 42190 9222 42192 9274
rect 41946 9220 41952 9222
rect 42008 9220 42032 9222
rect 42088 9220 42112 9222
rect 42168 9220 42192 9222
rect 42248 9220 42254 9222
rect 41946 9211 42254 9220
rect 41306 8732 41614 8741
rect 41306 8730 41312 8732
rect 41368 8730 41392 8732
rect 41448 8730 41472 8732
rect 41528 8730 41552 8732
rect 41608 8730 41614 8732
rect 41368 8678 41370 8730
rect 41550 8678 41552 8730
rect 41306 8676 41312 8678
rect 41368 8676 41392 8678
rect 41448 8676 41472 8678
rect 41528 8676 41552 8678
rect 41608 8676 41614 8678
rect 41306 8667 41614 8676
rect 41946 8188 42254 8197
rect 41946 8186 41952 8188
rect 42008 8186 42032 8188
rect 42088 8186 42112 8188
rect 42168 8186 42192 8188
rect 42248 8186 42254 8188
rect 42008 8134 42010 8186
rect 42190 8134 42192 8186
rect 41946 8132 41952 8134
rect 42008 8132 42032 8134
rect 42088 8132 42112 8134
rect 42168 8132 42192 8134
rect 42248 8132 42254 8134
rect 41946 8123 42254 8132
rect 41306 7644 41614 7653
rect 41306 7642 41312 7644
rect 41368 7642 41392 7644
rect 41448 7642 41472 7644
rect 41528 7642 41552 7644
rect 41608 7642 41614 7644
rect 41368 7590 41370 7642
rect 41550 7590 41552 7642
rect 41306 7588 41312 7590
rect 41368 7588 41392 7590
rect 41448 7588 41472 7590
rect 41528 7588 41552 7590
rect 41608 7588 41614 7590
rect 41306 7579 41614 7588
rect 41946 7100 42254 7109
rect 41946 7098 41952 7100
rect 42008 7098 42032 7100
rect 42088 7098 42112 7100
rect 42168 7098 42192 7100
rect 42248 7098 42254 7100
rect 42008 7046 42010 7098
rect 42190 7046 42192 7098
rect 41946 7044 41952 7046
rect 42008 7044 42032 7046
rect 42088 7044 42112 7046
rect 42168 7044 42192 7046
rect 42248 7044 42254 7046
rect 41946 7035 42254 7044
rect 41306 6556 41614 6565
rect 41306 6554 41312 6556
rect 41368 6554 41392 6556
rect 41448 6554 41472 6556
rect 41528 6554 41552 6556
rect 41608 6554 41614 6556
rect 41368 6502 41370 6554
rect 41550 6502 41552 6554
rect 41306 6500 41312 6502
rect 41368 6500 41392 6502
rect 41448 6500 41472 6502
rect 41528 6500 41552 6502
rect 41608 6500 41614 6502
rect 41306 6491 41614 6500
rect 41946 6012 42254 6021
rect 41946 6010 41952 6012
rect 42008 6010 42032 6012
rect 42088 6010 42112 6012
rect 42168 6010 42192 6012
rect 42248 6010 42254 6012
rect 42008 5958 42010 6010
rect 42190 5958 42192 6010
rect 41946 5956 41952 5958
rect 42008 5956 42032 5958
rect 42088 5956 42112 5958
rect 42168 5956 42192 5958
rect 42248 5956 42254 5958
rect 41946 5947 42254 5956
rect 41306 5468 41614 5477
rect 41306 5466 41312 5468
rect 41368 5466 41392 5468
rect 41448 5466 41472 5468
rect 41528 5466 41552 5468
rect 41608 5466 41614 5468
rect 41368 5414 41370 5466
rect 41550 5414 41552 5466
rect 41306 5412 41312 5414
rect 41368 5412 41392 5414
rect 41448 5412 41472 5414
rect 41528 5412 41552 5414
rect 41608 5412 41614 5414
rect 41306 5403 41614 5412
rect 41946 4924 42254 4933
rect 41946 4922 41952 4924
rect 42008 4922 42032 4924
rect 42088 4922 42112 4924
rect 42168 4922 42192 4924
rect 42248 4922 42254 4924
rect 42008 4870 42010 4922
rect 42190 4870 42192 4922
rect 41946 4868 41952 4870
rect 42008 4868 42032 4870
rect 42088 4868 42112 4870
rect 42168 4868 42192 4870
rect 42248 4868 42254 4870
rect 41946 4859 42254 4868
rect 41306 4380 41614 4389
rect 41306 4378 41312 4380
rect 41368 4378 41392 4380
rect 41448 4378 41472 4380
rect 41528 4378 41552 4380
rect 41608 4378 41614 4380
rect 41368 4326 41370 4378
rect 41550 4326 41552 4378
rect 41306 4324 41312 4326
rect 41368 4324 41392 4326
rect 41448 4324 41472 4326
rect 41528 4324 41552 4326
rect 41608 4324 41614 4326
rect 41306 4315 41614 4324
rect 41946 3836 42254 3845
rect 41946 3834 41952 3836
rect 42008 3834 42032 3836
rect 42088 3834 42112 3836
rect 42168 3834 42192 3836
rect 42248 3834 42254 3836
rect 42008 3782 42010 3834
rect 42190 3782 42192 3834
rect 41946 3780 41952 3782
rect 42008 3780 42032 3782
rect 42088 3780 42112 3782
rect 42168 3780 42192 3782
rect 42248 3780 42254 3782
rect 41946 3771 42254 3780
rect 41306 3292 41614 3301
rect 41306 3290 41312 3292
rect 41368 3290 41392 3292
rect 41448 3290 41472 3292
rect 41528 3290 41552 3292
rect 41608 3290 41614 3292
rect 41368 3238 41370 3290
rect 41550 3238 41552 3290
rect 41306 3236 41312 3238
rect 41368 3236 41392 3238
rect 41448 3236 41472 3238
rect 41528 3236 41552 3238
rect 41608 3236 41614 3238
rect 41306 3227 41614 3236
rect 41946 2748 42254 2757
rect 41946 2746 41952 2748
rect 42008 2746 42032 2748
rect 42088 2746 42112 2748
rect 42168 2746 42192 2748
rect 42248 2746 42254 2748
rect 42008 2694 42010 2746
rect 42190 2694 42192 2746
rect 41946 2692 41952 2694
rect 42008 2692 42032 2694
rect 42088 2692 42112 2694
rect 42168 2692 42192 2694
rect 42248 2692 42254 2694
rect 41946 2683 42254 2692
rect 40684 2508 40736 2514
rect 40684 2450 40736 2456
rect 40500 2304 40552 2310
rect 40500 2246 40552 2252
rect 40224 2100 40276 2106
rect 40224 2042 40276 2048
rect 40132 1896 40184 1902
rect 40132 1838 40184 1844
rect 40040 1556 40092 1562
rect 40040 1498 40092 1504
rect 39816 1448 39896 1476
rect 39764 1430 39816 1436
rect 40040 1420 40092 1426
rect 40040 1362 40092 1368
rect 39592 1278 39804 1306
rect 39776 400 39804 1278
rect 39948 1216 40000 1222
rect 39948 1158 40000 1164
rect 39960 474 39988 1158
rect 40052 882 40080 1362
rect 40144 1358 40172 1838
rect 40132 1352 40184 1358
rect 40132 1294 40184 1300
rect 40040 876 40092 882
rect 40040 818 40092 824
rect 40236 762 40264 2042
rect 40408 1760 40460 1766
rect 40408 1702 40460 1708
rect 40420 1601 40448 1702
rect 40406 1592 40462 1601
rect 40406 1527 40462 1536
rect 40512 1426 40540 2246
rect 40500 1420 40552 1426
rect 40500 1362 40552 1368
rect 40408 1284 40460 1290
rect 40408 1226 40460 1232
rect 40316 944 40368 950
rect 40316 886 40368 892
rect 40052 734 40264 762
rect 39948 468 40000 474
rect 39948 410 40000 416
rect 40052 400 40080 734
rect 40328 660 40356 886
rect 40420 814 40448 1226
rect 40696 814 40724 2450
rect 41306 2204 41614 2213
rect 41306 2202 41312 2204
rect 41368 2202 41392 2204
rect 41448 2202 41472 2204
rect 41528 2202 41552 2204
rect 41608 2202 41614 2204
rect 41368 2150 41370 2202
rect 41550 2150 41552 2202
rect 41306 2148 41312 2150
rect 41368 2148 41392 2150
rect 41448 2148 41472 2150
rect 41528 2148 41552 2150
rect 41608 2148 41614 2150
rect 41306 2139 41614 2148
rect 40868 1896 40920 1902
rect 40868 1838 40920 1844
rect 40776 1760 40828 1766
rect 40776 1702 40828 1708
rect 40788 950 40816 1702
rect 40776 944 40828 950
rect 40776 886 40828 892
rect 40408 808 40460 814
rect 40500 808 40552 814
rect 40408 750 40460 756
rect 40498 776 40500 785
rect 40684 808 40736 814
rect 40552 776 40554 785
rect 40684 750 40736 756
rect 40498 711 40554 720
rect 40236 632 40356 660
rect 40408 672 40460 678
rect 40406 640 40408 649
rect 40776 672 40828 678
rect 40460 640 40462 649
rect 39304 128 39356 134
rect 39304 70 39356 76
rect 39486 0 39542 400
rect 39762 0 39818 400
rect 40038 0 40094 400
rect 40236 66 40264 632
rect 40776 614 40828 620
rect 40406 575 40462 584
rect 40328 474 40448 490
rect 40328 468 40460 474
rect 40328 462 40408 468
rect 40328 400 40356 462
rect 40408 410 40460 416
rect 40604 462 40724 490
rect 40604 400 40632 462
rect 40224 60 40276 66
rect 40224 2 40276 8
rect 40314 0 40370 400
rect 40590 0 40646 400
rect 40696 270 40724 462
rect 40788 406 40816 614
rect 40776 400 40828 406
rect 40880 400 40908 1838
rect 41946 1660 42254 1669
rect 41946 1658 41952 1660
rect 42008 1658 42032 1660
rect 42088 1658 42112 1660
rect 42168 1658 42192 1660
rect 42248 1658 42254 1660
rect 42008 1606 42010 1658
rect 42190 1606 42192 1658
rect 41946 1604 41952 1606
rect 42008 1604 42032 1606
rect 42088 1604 42112 1606
rect 42168 1604 42192 1606
rect 42248 1604 42254 1606
rect 41946 1595 42254 1604
rect 41144 1488 41196 1494
rect 41144 1430 41196 1436
rect 40960 1284 41012 1290
rect 40960 1226 41012 1232
rect 40776 342 40828 348
rect 40684 264 40736 270
rect 40684 206 40736 212
rect 40866 0 40922 400
rect 40972 202 41000 1226
rect 41052 876 41104 882
rect 41052 818 41104 824
rect 41064 474 41092 818
rect 41052 468 41104 474
rect 41052 410 41104 416
rect 41156 400 41184 1430
rect 41248 1290 41368 1306
rect 41248 1284 41380 1290
rect 41248 1278 41328 1284
rect 41248 1018 41276 1278
rect 41328 1226 41380 1232
rect 41972 1216 42024 1222
rect 41972 1158 42024 1164
rect 41306 1116 41614 1125
rect 41306 1114 41312 1116
rect 41368 1114 41392 1116
rect 41448 1114 41472 1116
rect 41528 1114 41552 1116
rect 41608 1114 41614 1116
rect 41368 1062 41370 1114
rect 41550 1062 41552 1114
rect 41306 1060 41312 1062
rect 41368 1060 41392 1062
rect 41448 1060 41472 1062
rect 41528 1060 41552 1062
rect 41608 1060 41614 1062
rect 41306 1051 41614 1060
rect 41236 1012 41288 1018
rect 41236 954 41288 960
rect 41788 1012 41840 1018
rect 41788 954 41840 960
rect 40960 196 41012 202
rect 40960 138 41012 144
rect 41142 0 41198 400
rect 41248 270 41276 954
rect 41800 921 41828 954
rect 41786 912 41842 921
rect 41984 882 42012 1158
rect 41786 847 41842 856
rect 41972 876 42024 882
rect 41972 818 42024 824
rect 41328 808 41380 814
rect 42340 808 42392 814
rect 41328 750 41380 756
rect 42338 776 42340 785
rect 42392 776 42394 785
rect 41340 649 41368 750
rect 42338 711 42394 720
rect 41512 672 41564 678
rect 41326 640 41382 649
rect 41512 614 41564 620
rect 41788 672 41840 678
rect 41788 614 41840 620
rect 41326 575 41382 584
rect 41524 338 41552 614
rect 41512 332 41564 338
rect 41512 274 41564 280
rect 41800 270 41828 614
rect 41946 572 42254 581
rect 41946 570 41952 572
rect 42008 570 42032 572
rect 42088 570 42112 572
rect 42168 570 42192 572
rect 42248 570 42254 572
rect 42008 518 42010 570
rect 42190 518 42192 570
rect 41946 516 41952 518
rect 42008 516 42032 518
rect 42088 516 42112 518
rect 42168 516 42192 518
rect 42248 516 42254 518
rect 41946 507 42254 516
rect 41236 264 41288 270
rect 41236 206 41288 212
rect 41788 264 41840 270
rect 41788 206 41840 212
<< via2 >>
rect 1952 11450 2008 11452
rect 2032 11450 2088 11452
rect 2112 11450 2168 11452
rect 2192 11450 2248 11452
rect 1952 11398 1998 11450
rect 1998 11398 2008 11450
rect 2032 11398 2062 11450
rect 2062 11398 2074 11450
rect 2074 11398 2088 11450
rect 2112 11398 2126 11450
rect 2126 11398 2138 11450
rect 2138 11398 2168 11450
rect 2192 11398 2202 11450
rect 2202 11398 2248 11450
rect 1952 11396 2008 11398
rect 2032 11396 2088 11398
rect 2112 11396 2168 11398
rect 2192 11396 2248 11398
rect 1312 10906 1368 10908
rect 1392 10906 1448 10908
rect 1472 10906 1528 10908
rect 1552 10906 1608 10908
rect 1312 10854 1358 10906
rect 1358 10854 1368 10906
rect 1392 10854 1422 10906
rect 1422 10854 1434 10906
rect 1434 10854 1448 10906
rect 1472 10854 1486 10906
rect 1486 10854 1498 10906
rect 1498 10854 1528 10906
rect 1552 10854 1562 10906
rect 1562 10854 1608 10906
rect 1312 10852 1368 10854
rect 1392 10852 1448 10854
rect 1472 10852 1528 10854
rect 1552 10852 1608 10854
rect 1952 10362 2008 10364
rect 2032 10362 2088 10364
rect 2112 10362 2168 10364
rect 2192 10362 2248 10364
rect 1952 10310 1998 10362
rect 1998 10310 2008 10362
rect 2032 10310 2062 10362
rect 2062 10310 2074 10362
rect 2074 10310 2088 10362
rect 2112 10310 2126 10362
rect 2126 10310 2138 10362
rect 2138 10310 2168 10362
rect 2192 10310 2202 10362
rect 2202 10310 2248 10362
rect 1952 10308 2008 10310
rect 2032 10308 2088 10310
rect 2112 10308 2168 10310
rect 2192 10308 2248 10310
rect 1312 9818 1368 9820
rect 1392 9818 1448 9820
rect 1472 9818 1528 9820
rect 1552 9818 1608 9820
rect 1312 9766 1358 9818
rect 1358 9766 1368 9818
rect 1392 9766 1422 9818
rect 1422 9766 1434 9818
rect 1434 9766 1448 9818
rect 1472 9766 1486 9818
rect 1486 9766 1498 9818
rect 1498 9766 1528 9818
rect 1552 9766 1562 9818
rect 1562 9766 1608 9818
rect 1312 9764 1368 9766
rect 1392 9764 1448 9766
rect 1472 9764 1528 9766
rect 1552 9764 1608 9766
rect 1952 9274 2008 9276
rect 2032 9274 2088 9276
rect 2112 9274 2168 9276
rect 2192 9274 2248 9276
rect 1952 9222 1998 9274
rect 1998 9222 2008 9274
rect 2032 9222 2062 9274
rect 2062 9222 2074 9274
rect 2074 9222 2088 9274
rect 2112 9222 2126 9274
rect 2126 9222 2138 9274
rect 2138 9222 2168 9274
rect 2192 9222 2202 9274
rect 2202 9222 2248 9274
rect 1952 9220 2008 9222
rect 2032 9220 2088 9222
rect 2112 9220 2168 9222
rect 2192 9220 2248 9222
rect 1312 8730 1368 8732
rect 1392 8730 1448 8732
rect 1472 8730 1528 8732
rect 1552 8730 1608 8732
rect 1312 8678 1358 8730
rect 1358 8678 1368 8730
rect 1392 8678 1422 8730
rect 1422 8678 1434 8730
rect 1434 8678 1448 8730
rect 1472 8678 1486 8730
rect 1486 8678 1498 8730
rect 1498 8678 1528 8730
rect 1552 8678 1562 8730
rect 1562 8678 1608 8730
rect 1312 8676 1368 8678
rect 1392 8676 1448 8678
rect 1472 8676 1528 8678
rect 1552 8676 1608 8678
rect 1952 8186 2008 8188
rect 2032 8186 2088 8188
rect 2112 8186 2168 8188
rect 2192 8186 2248 8188
rect 1952 8134 1998 8186
rect 1998 8134 2008 8186
rect 2032 8134 2062 8186
rect 2062 8134 2074 8186
rect 2074 8134 2088 8186
rect 2112 8134 2126 8186
rect 2126 8134 2138 8186
rect 2138 8134 2168 8186
rect 2192 8134 2202 8186
rect 2202 8134 2248 8186
rect 1952 8132 2008 8134
rect 2032 8132 2088 8134
rect 2112 8132 2168 8134
rect 2192 8132 2248 8134
rect 5170 8200 5226 8256
rect 1312 7642 1368 7644
rect 1392 7642 1448 7644
rect 1472 7642 1528 7644
rect 1552 7642 1608 7644
rect 1312 7590 1358 7642
rect 1358 7590 1368 7642
rect 1392 7590 1422 7642
rect 1422 7590 1434 7642
rect 1434 7590 1448 7642
rect 1472 7590 1486 7642
rect 1486 7590 1498 7642
rect 1498 7590 1528 7642
rect 1552 7590 1562 7642
rect 1562 7590 1608 7642
rect 1312 7588 1368 7590
rect 1392 7588 1448 7590
rect 1472 7588 1528 7590
rect 1552 7588 1608 7590
rect 1952 7098 2008 7100
rect 2032 7098 2088 7100
rect 2112 7098 2168 7100
rect 2192 7098 2248 7100
rect 1952 7046 1998 7098
rect 1998 7046 2008 7098
rect 2032 7046 2062 7098
rect 2062 7046 2074 7098
rect 2074 7046 2088 7098
rect 2112 7046 2126 7098
rect 2126 7046 2138 7098
rect 2138 7046 2168 7098
rect 2192 7046 2202 7098
rect 2202 7046 2248 7098
rect 1952 7044 2008 7046
rect 2032 7044 2088 7046
rect 2112 7044 2168 7046
rect 2192 7044 2248 7046
rect 1312 6554 1368 6556
rect 1392 6554 1448 6556
rect 1472 6554 1528 6556
rect 1552 6554 1608 6556
rect 1312 6502 1358 6554
rect 1358 6502 1368 6554
rect 1392 6502 1422 6554
rect 1422 6502 1434 6554
rect 1434 6502 1448 6554
rect 1472 6502 1486 6554
rect 1486 6502 1498 6554
rect 1498 6502 1528 6554
rect 1552 6502 1562 6554
rect 1562 6502 1608 6554
rect 1312 6500 1368 6502
rect 1392 6500 1448 6502
rect 1472 6500 1528 6502
rect 1552 6500 1608 6502
rect 1952 6010 2008 6012
rect 2032 6010 2088 6012
rect 2112 6010 2168 6012
rect 2192 6010 2248 6012
rect 1952 5958 1998 6010
rect 1998 5958 2008 6010
rect 2032 5958 2062 6010
rect 2062 5958 2074 6010
rect 2074 5958 2088 6010
rect 2112 5958 2126 6010
rect 2126 5958 2138 6010
rect 2138 5958 2168 6010
rect 2192 5958 2202 6010
rect 2202 5958 2248 6010
rect 1952 5956 2008 5958
rect 2032 5956 2088 5958
rect 2112 5956 2168 5958
rect 2192 5956 2248 5958
rect 1312 5466 1368 5468
rect 1392 5466 1448 5468
rect 1472 5466 1528 5468
rect 1552 5466 1608 5468
rect 1312 5414 1358 5466
rect 1358 5414 1368 5466
rect 1392 5414 1422 5466
rect 1422 5414 1434 5466
rect 1434 5414 1448 5466
rect 1472 5414 1486 5466
rect 1486 5414 1498 5466
rect 1498 5414 1528 5466
rect 1552 5414 1562 5466
rect 1562 5414 1608 5466
rect 1312 5412 1368 5414
rect 1392 5412 1448 5414
rect 1472 5412 1528 5414
rect 1552 5412 1608 5414
rect 1952 4922 2008 4924
rect 2032 4922 2088 4924
rect 2112 4922 2168 4924
rect 2192 4922 2248 4924
rect 1952 4870 1998 4922
rect 1998 4870 2008 4922
rect 2032 4870 2062 4922
rect 2062 4870 2074 4922
rect 2074 4870 2088 4922
rect 2112 4870 2126 4922
rect 2126 4870 2138 4922
rect 2138 4870 2168 4922
rect 2192 4870 2202 4922
rect 2202 4870 2248 4922
rect 1952 4868 2008 4870
rect 2032 4868 2088 4870
rect 2112 4868 2168 4870
rect 2192 4868 2248 4870
rect 1312 4378 1368 4380
rect 1392 4378 1448 4380
rect 1472 4378 1528 4380
rect 1552 4378 1608 4380
rect 1312 4326 1358 4378
rect 1358 4326 1368 4378
rect 1392 4326 1422 4378
rect 1422 4326 1434 4378
rect 1434 4326 1448 4378
rect 1472 4326 1486 4378
rect 1486 4326 1498 4378
rect 1498 4326 1528 4378
rect 1552 4326 1562 4378
rect 1562 4326 1608 4378
rect 1312 4324 1368 4326
rect 1392 4324 1448 4326
rect 1472 4324 1528 4326
rect 1552 4324 1608 4326
rect 1952 3834 2008 3836
rect 2032 3834 2088 3836
rect 2112 3834 2168 3836
rect 2192 3834 2248 3836
rect 1952 3782 1998 3834
rect 1998 3782 2008 3834
rect 2032 3782 2062 3834
rect 2062 3782 2074 3834
rect 2074 3782 2088 3834
rect 2112 3782 2126 3834
rect 2126 3782 2138 3834
rect 2138 3782 2168 3834
rect 2192 3782 2202 3834
rect 2202 3782 2248 3834
rect 1952 3780 2008 3782
rect 2032 3780 2088 3782
rect 2112 3780 2168 3782
rect 2192 3780 2248 3782
rect 1312 3290 1368 3292
rect 1392 3290 1448 3292
rect 1472 3290 1528 3292
rect 1552 3290 1608 3292
rect 1312 3238 1358 3290
rect 1358 3238 1368 3290
rect 1392 3238 1422 3290
rect 1422 3238 1434 3290
rect 1434 3238 1448 3290
rect 1472 3238 1486 3290
rect 1486 3238 1498 3290
rect 1498 3238 1528 3290
rect 1552 3238 1562 3290
rect 1562 3238 1608 3290
rect 1312 3236 1368 3238
rect 1392 3236 1448 3238
rect 1472 3236 1528 3238
rect 1552 3236 1608 3238
rect 1952 2746 2008 2748
rect 2032 2746 2088 2748
rect 2112 2746 2168 2748
rect 2192 2746 2248 2748
rect 1952 2694 1998 2746
rect 1998 2694 2008 2746
rect 2032 2694 2062 2746
rect 2062 2694 2074 2746
rect 2074 2694 2088 2746
rect 2112 2694 2126 2746
rect 2126 2694 2138 2746
rect 2138 2694 2168 2746
rect 2192 2694 2202 2746
rect 2202 2694 2248 2746
rect 1952 2692 2008 2694
rect 2032 2692 2088 2694
rect 2112 2692 2168 2694
rect 2192 2692 2248 2694
rect 1312 2202 1368 2204
rect 1392 2202 1448 2204
rect 1472 2202 1528 2204
rect 1552 2202 1608 2204
rect 1312 2150 1358 2202
rect 1358 2150 1368 2202
rect 1392 2150 1422 2202
rect 1422 2150 1434 2202
rect 1434 2150 1448 2202
rect 1472 2150 1486 2202
rect 1486 2150 1498 2202
rect 1498 2150 1528 2202
rect 1552 2150 1562 2202
rect 1562 2150 1608 2202
rect 1312 2148 1368 2150
rect 1392 2148 1448 2150
rect 1472 2148 1528 2150
rect 1552 2148 1608 2150
rect 1952 1658 2008 1660
rect 2032 1658 2088 1660
rect 2112 1658 2168 1660
rect 2192 1658 2248 1660
rect 1952 1606 1998 1658
rect 1998 1606 2008 1658
rect 2032 1606 2062 1658
rect 2062 1606 2074 1658
rect 2074 1606 2088 1658
rect 2112 1606 2126 1658
rect 2126 1606 2138 1658
rect 2138 1606 2168 1658
rect 2192 1606 2202 1658
rect 2202 1606 2248 1658
rect 1952 1604 2008 1606
rect 2032 1604 2088 1606
rect 2112 1604 2168 1606
rect 2192 1604 2248 1606
rect 1312 1114 1368 1116
rect 1392 1114 1448 1116
rect 1472 1114 1528 1116
rect 1552 1114 1608 1116
rect 1312 1062 1358 1114
rect 1358 1062 1368 1114
rect 1392 1062 1422 1114
rect 1422 1062 1434 1114
rect 1434 1062 1448 1114
rect 1472 1062 1486 1114
rect 1486 1062 1498 1114
rect 1498 1062 1528 1114
rect 1552 1062 1562 1114
rect 1562 1062 1608 1114
rect 1312 1060 1368 1062
rect 1392 1060 1448 1062
rect 1472 1060 1528 1062
rect 1552 1060 1608 1062
rect 1952 570 2008 572
rect 2032 570 2088 572
rect 2112 570 2168 572
rect 2192 570 2248 572
rect 1952 518 1998 570
rect 1998 518 2008 570
rect 2032 518 2062 570
rect 2062 518 2074 570
rect 2074 518 2088 570
rect 2112 518 2126 570
rect 2126 518 2138 570
rect 2138 518 2168 570
rect 2192 518 2202 570
rect 2202 518 2248 570
rect 1952 516 2008 518
rect 2032 516 2088 518
rect 2112 516 2168 518
rect 2192 516 2248 518
rect 4894 7928 4950 7984
rect 4986 7404 5042 7440
rect 4986 7384 4988 7404
rect 4988 7384 5040 7404
rect 5040 7384 5042 7404
rect 4894 6740 4896 6760
rect 4896 6740 4948 6760
rect 4948 6740 4950 6760
rect 4894 6704 4950 6740
rect 6826 7828 6828 7848
rect 6828 7828 6880 7848
rect 6880 7828 6882 7848
rect 6826 7792 6882 7828
rect 6274 6160 6330 6216
rect 7378 8472 7434 8528
rect 7102 6296 7158 6352
rect 8114 7248 8170 7304
rect 9312 10906 9368 10908
rect 9392 10906 9448 10908
rect 9472 10906 9528 10908
rect 9552 10906 9608 10908
rect 9312 10854 9358 10906
rect 9358 10854 9368 10906
rect 9392 10854 9422 10906
rect 9422 10854 9434 10906
rect 9434 10854 9448 10906
rect 9472 10854 9486 10906
rect 9486 10854 9498 10906
rect 9498 10854 9528 10906
rect 9552 10854 9562 10906
rect 9562 10854 9608 10906
rect 9312 10852 9368 10854
rect 9392 10852 9448 10854
rect 9472 10852 9528 10854
rect 9552 10852 9608 10854
rect 9312 9818 9368 9820
rect 9392 9818 9448 9820
rect 9472 9818 9528 9820
rect 9552 9818 9608 9820
rect 9312 9766 9358 9818
rect 9358 9766 9368 9818
rect 9392 9766 9422 9818
rect 9422 9766 9434 9818
rect 9434 9766 9448 9818
rect 9472 9766 9486 9818
rect 9486 9766 9498 9818
rect 9498 9766 9528 9818
rect 9552 9766 9562 9818
rect 9562 9766 9608 9818
rect 9312 9764 9368 9766
rect 9392 9764 9448 9766
rect 9472 9764 9528 9766
rect 9552 9764 9608 9766
rect 9952 11450 10008 11452
rect 10032 11450 10088 11452
rect 10112 11450 10168 11452
rect 10192 11450 10248 11452
rect 9952 11398 9998 11450
rect 9998 11398 10008 11450
rect 10032 11398 10062 11450
rect 10062 11398 10074 11450
rect 10074 11398 10088 11450
rect 10112 11398 10126 11450
rect 10126 11398 10138 11450
rect 10138 11398 10168 11450
rect 10192 11398 10202 11450
rect 10202 11398 10248 11450
rect 9952 11396 10008 11398
rect 10032 11396 10088 11398
rect 10112 11396 10168 11398
rect 10192 11396 10248 11398
rect 9952 10362 10008 10364
rect 10032 10362 10088 10364
rect 10112 10362 10168 10364
rect 10192 10362 10248 10364
rect 9952 10310 9998 10362
rect 9998 10310 10008 10362
rect 10032 10310 10062 10362
rect 10062 10310 10074 10362
rect 10074 10310 10088 10362
rect 10112 10310 10126 10362
rect 10126 10310 10138 10362
rect 10138 10310 10168 10362
rect 10192 10310 10202 10362
rect 10202 10310 10248 10362
rect 9952 10308 10008 10310
rect 10032 10308 10088 10310
rect 10112 10308 10168 10310
rect 10192 10308 10248 10310
rect 9952 9274 10008 9276
rect 10032 9274 10088 9276
rect 10112 9274 10168 9276
rect 10192 9274 10248 9276
rect 9952 9222 9998 9274
rect 9998 9222 10008 9274
rect 10032 9222 10062 9274
rect 10062 9222 10074 9274
rect 10074 9222 10088 9274
rect 10112 9222 10126 9274
rect 10126 9222 10138 9274
rect 10138 9222 10168 9274
rect 10192 9222 10202 9274
rect 10202 9222 10248 9274
rect 9952 9220 10008 9222
rect 10032 9220 10088 9222
rect 10112 9220 10168 9222
rect 10192 9220 10248 9222
rect 9770 8744 9826 8800
rect 9312 8730 9368 8732
rect 9392 8730 9448 8732
rect 9472 8730 9528 8732
rect 9552 8730 9608 8732
rect 9312 8678 9358 8730
rect 9358 8678 9368 8730
rect 9392 8678 9422 8730
rect 9422 8678 9434 8730
rect 9434 8678 9448 8730
rect 9472 8678 9486 8730
rect 9486 8678 9498 8730
rect 9498 8678 9528 8730
rect 9552 8678 9562 8730
rect 9562 8678 9608 8730
rect 9312 8676 9368 8678
rect 9392 8676 9448 8678
rect 9472 8676 9528 8678
rect 9552 8676 9608 8678
rect 9678 8064 9734 8120
rect 9952 8186 10008 8188
rect 10032 8186 10088 8188
rect 10112 8186 10168 8188
rect 10192 8186 10248 8188
rect 9952 8134 9998 8186
rect 9998 8134 10008 8186
rect 10032 8134 10062 8186
rect 10062 8134 10074 8186
rect 10074 8134 10088 8186
rect 10112 8134 10126 8186
rect 10126 8134 10138 8186
rect 10138 8134 10168 8186
rect 10192 8134 10202 8186
rect 10202 8134 10248 8186
rect 9952 8132 10008 8134
rect 10032 8132 10088 8134
rect 10112 8132 10168 8134
rect 10192 8132 10248 8134
rect 10690 9016 10746 9072
rect 9312 7642 9368 7644
rect 9392 7642 9448 7644
rect 9472 7642 9528 7644
rect 9552 7642 9608 7644
rect 9312 7590 9358 7642
rect 9358 7590 9368 7642
rect 9392 7590 9422 7642
rect 9422 7590 9434 7642
rect 9434 7590 9448 7642
rect 9472 7590 9486 7642
rect 9486 7590 9498 7642
rect 9498 7590 9528 7642
rect 9552 7590 9562 7642
rect 9562 7590 9608 7642
rect 9312 7588 9368 7590
rect 9392 7588 9448 7590
rect 9472 7588 9528 7590
rect 9552 7588 9608 7590
rect 10138 7520 10194 7576
rect 9952 7098 10008 7100
rect 10032 7098 10088 7100
rect 10112 7098 10168 7100
rect 10192 7098 10248 7100
rect 9952 7046 9998 7098
rect 9998 7046 10008 7098
rect 10032 7046 10062 7098
rect 10062 7046 10074 7098
rect 10074 7046 10088 7098
rect 10112 7046 10126 7098
rect 10126 7046 10138 7098
rect 10138 7046 10168 7098
rect 10192 7046 10202 7098
rect 10202 7046 10248 7098
rect 9952 7044 10008 7046
rect 10032 7044 10088 7046
rect 10112 7044 10168 7046
rect 10192 7044 10248 7046
rect 9494 6860 9550 6896
rect 9494 6840 9496 6860
rect 9496 6840 9548 6860
rect 9548 6840 9550 6860
rect 9312 6554 9368 6556
rect 9392 6554 9448 6556
rect 9472 6554 9528 6556
rect 9552 6554 9608 6556
rect 9312 6502 9358 6554
rect 9358 6502 9368 6554
rect 9392 6502 9422 6554
rect 9422 6502 9434 6554
rect 9434 6502 9448 6554
rect 9472 6502 9486 6554
rect 9486 6502 9498 6554
rect 9498 6502 9528 6554
rect 9552 6502 9562 6554
rect 9562 6502 9608 6554
rect 9312 6500 9368 6502
rect 9392 6500 9448 6502
rect 9472 6500 9528 6502
rect 9552 6500 9608 6502
rect 9770 6432 9826 6488
rect 10138 6568 10194 6624
rect 9952 6010 10008 6012
rect 10032 6010 10088 6012
rect 10112 6010 10168 6012
rect 10192 6010 10248 6012
rect 9952 5958 9998 6010
rect 9998 5958 10008 6010
rect 10032 5958 10062 6010
rect 10062 5958 10074 6010
rect 10074 5958 10088 6010
rect 10112 5958 10126 6010
rect 10126 5958 10138 6010
rect 10138 5958 10168 6010
rect 10192 5958 10202 6010
rect 10202 5958 10248 6010
rect 9952 5956 10008 5958
rect 10032 5956 10088 5958
rect 10112 5956 10168 5958
rect 10192 5956 10248 5958
rect 9312 5466 9368 5468
rect 9392 5466 9448 5468
rect 9472 5466 9528 5468
rect 9552 5466 9608 5468
rect 9312 5414 9358 5466
rect 9358 5414 9368 5466
rect 9392 5414 9422 5466
rect 9422 5414 9434 5466
rect 9434 5414 9448 5466
rect 9472 5414 9486 5466
rect 9486 5414 9498 5466
rect 9498 5414 9528 5466
rect 9552 5414 9562 5466
rect 9562 5414 9608 5466
rect 9312 5412 9368 5414
rect 9392 5412 9448 5414
rect 9472 5412 9528 5414
rect 9552 5412 9608 5414
rect 9312 4378 9368 4380
rect 9392 4378 9448 4380
rect 9472 4378 9528 4380
rect 9552 4378 9608 4380
rect 9312 4326 9358 4378
rect 9358 4326 9368 4378
rect 9392 4326 9422 4378
rect 9422 4326 9434 4378
rect 9434 4326 9448 4378
rect 9472 4326 9486 4378
rect 9486 4326 9498 4378
rect 9498 4326 9528 4378
rect 9552 4326 9562 4378
rect 9562 4326 9608 4378
rect 9312 4324 9368 4326
rect 9392 4324 9448 4326
rect 9472 4324 9528 4326
rect 9552 4324 9608 4326
rect 9678 3984 9734 4040
rect 9312 3290 9368 3292
rect 9392 3290 9448 3292
rect 9472 3290 9528 3292
rect 9552 3290 9608 3292
rect 9312 3238 9358 3290
rect 9358 3238 9368 3290
rect 9392 3238 9422 3290
rect 9422 3238 9434 3290
rect 9434 3238 9448 3290
rect 9472 3238 9486 3290
rect 9486 3238 9498 3290
rect 9498 3238 9528 3290
rect 9552 3238 9562 3290
rect 9562 3238 9608 3290
rect 9312 3236 9368 3238
rect 9392 3236 9448 3238
rect 9472 3236 9528 3238
rect 9552 3236 9608 3238
rect 9312 2202 9368 2204
rect 9392 2202 9448 2204
rect 9472 2202 9528 2204
rect 9552 2202 9608 2204
rect 9312 2150 9358 2202
rect 9358 2150 9368 2202
rect 9392 2150 9422 2202
rect 9422 2150 9434 2202
rect 9434 2150 9448 2202
rect 9472 2150 9486 2202
rect 9486 2150 9498 2202
rect 9498 2150 9528 2202
rect 9552 2150 9562 2202
rect 9562 2150 9608 2202
rect 9312 2148 9368 2150
rect 9392 2148 9448 2150
rect 9472 2148 9528 2150
rect 9552 2148 9608 2150
rect 9312 1114 9368 1116
rect 9392 1114 9448 1116
rect 9472 1114 9528 1116
rect 9552 1114 9608 1116
rect 9312 1062 9358 1114
rect 9358 1062 9368 1114
rect 9392 1062 9422 1114
rect 9422 1062 9434 1114
rect 9434 1062 9448 1114
rect 9472 1062 9486 1114
rect 9486 1062 9498 1114
rect 9498 1062 9528 1114
rect 9552 1062 9562 1114
rect 9562 1062 9608 1114
rect 9312 1060 9368 1062
rect 9392 1060 9448 1062
rect 9472 1060 9528 1062
rect 9552 1060 9608 1062
rect 9952 3834 10008 3836
rect 10032 3834 10088 3836
rect 10112 3834 10168 3836
rect 10192 3834 10248 3836
rect 9952 3782 9998 3834
rect 9998 3782 10008 3834
rect 10032 3782 10062 3834
rect 10062 3782 10074 3834
rect 10074 3782 10088 3834
rect 10112 3782 10126 3834
rect 10126 3782 10138 3834
rect 10138 3782 10168 3834
rect 10192 3782 10202 3834
rect 10202 3782 10248 3834
rect 9952 3780 10008 3782
rect 10032 3780 10088 3782
rect 10112 3780 10168 3782
rect 10192 3780 10248 3782
rect 9952 2746 10008 2748
rect 10032 2746 10088 2748
rect 10112 2746 10168 2748
rect 10192 2746 10248 2748
rect 9952 2694 9998 2746
rect 9998 2694 10008 2746
rect 10032 2694 10062 2746
rect 10062 2694 10074 2746
rect 10074 2694 10088 2746
rect 10112 2694 10126 2746
rect 10126 2694 10138 2746
rect 10138 2694 10168 2746
rect 10192 2694 10202 2746
rect 10202 2694 10248 2746
rect 9952 2692 10008 2694
rect 10032 2692 10088 2694
rect 10112 2692 10168 2694
rect 10192 2692 10248 2694
rect 9952 1658 10008 1660
rect 10032 1658 10088 1660
rect 10112 1658 10168 1660
rect 10192 1658 10248 1660
rect 9952 1606 9998 1658
rect 9998 1606 10008 1658
rect 10032 1606 10062 1658
rect 10062 1606 10074 1658
rect 10074 1606 10088 1658
rect 10112 1606 10126 1658
rect 10126 1606 10138 1658
rect 10138 1606 10168 1658
rect 10192 1606 10202 1658
rect 10202 1606 10248 1658
rect 9952 1604 10008 1606
rect 10032 1604 10088 1606
rect 10112 1604 10168 1606
rect 10192 1604 10248 1606
rect 9952 570 10008 572
rect 10032 570 10088 572
rect 10112 570 10168 572
rect 10192 570 10248 572
rect 9952 518 9998 570
rect 9998 518 10008 570
rect 10032 518 10062 570
rect 10062 518 10074 570
rect 10074 518 10088 570
rect 10112 518 10126 570
rect 10126 518 10138 570
rect 10138 518 10168 570
rect 10192 518 10202 570
rect 10202 518 10248 570
rect 9952 516 10008 518
rect 10032 516 10088 518
rect 10112 516 10168 518
rect 10192 516 10248 518
rect 10414 6976 10470 7032
rect 10690 8356 10746 8392
rect 10690 8336 10692 8356
rect 10692 8336 10744 8356
rect 10744 8336 10746 8356
rect 10690 8200 10746 8256
rect 10690 7520 10746 7576
rect 10874 9152 10930 9208
rect 11334 7520 11390 7576
rect 11518 7928 11574 7984
rect 11610 6976 11666 7032
rect 11886 7248 11942 7304
rect 11886 6976 11942 7032
rect 12254 8064 12310 8120
rect 12254 7248 12310 7304
rect 12622 8608 12678 8664
rect 12438 6976 12494 7032
rect 12438 1264 12494 1320
rect 13174 8336 13230 8392
rect 14002 9560 14058 9616
rect 14094 9460 14096 9480
rect 14096 9460 14148 9480
rect 14148 9460 14150 9480
rect 14094 9424 14150 9460
rect 14002 9016 14058 9072
rect 14370 9152 14426 9208
rect 14738 9016 14794 9072
rect 14922 9016 14978 9072
rect 14646 8880 14702 8936
rect 15106 8608 15162 8664
rect 13450 8356 13506 8392
rect 13450 8336 13452 8356
rect 13452 8336 13504 8356
rect 13504 8336 13506 8356
rect 14554 8200 14610 8256
rect 14738 8200 14794 8256
rect 14186 7792 14242 7848
rect 15658 9288 15714 9344
rect 15382 8200 15438 8256
rect 15014 7792 15070 7848
rect 15290 7656 15346 7712
rect 14416 7316 14472 7372
rect 15658 8472 15714 8528
rect 16026 9288 16082 9344
rect 15842 8880 15898 8936
rect 15934 8472 15990 8528
rect 16210 9460 16212 9480
rect 16212 9460 16264 9480
rect 16264 9460 16266 9480
rect 16210 9424 16266 9460
rect 16486 9172 16542 9208
rect 16486 9152 16488 9172
rect 16488 9152 16540 9172
rect 16540 9152 16542 9172
rect 16670 8744 16726 8800
rect 16578 8608 16634 8664
rect 17038 8880 17094 8936
rect 17312 10906 17368 10908
rect 17392 10906 17448 10908
rect 17472 10906 17528 10908
rect 17552 10906 17608 10908
rect 17312 10854 17358 10906
rect 17358 10854 17368 10906
rect 17392 10854 17422 10906
rect 17422 10854 17434 10906
rect 17434 10854 17448 10906
rect 17472 10854 17486 10906
rect 17486 10854 17498 10906
rect 17498 10854 17528 10906
rect 17552 10854 17562 10906
rect 17562 10854 17608 10906
rect 17312 10852 17368 10854
rect 17392 10852 17448 10854
rect 17472 10852 17528 10854
rect 17552 10852 17608 10854
rect 17952 11450 18008 11452
rect 18032 11450 18088 11452
rect 18112 11450 18168 11452
rect 18192 11450 18248 11452
rect 17952 11398 17998 11450
rect 17998 11398 18008 11450
rect 18032 11398 18062 11450
rect 18062 11398 18074 11450
rect 18074 11398 18088 11450
rect 18112 11398 18126 11450
rect 18126 11398 18138 11450
rect 18138 11398 18168 11450
rect 18192 11398 18202 11450
rect 18202 11398 18248 11450
rect 17952 11396 18008 11398
rect 18032 11396 18088 11398
rect 18112 11396 18168 11398
rect 18192 11396 18248 11398
rect 17952 10362 18008 10364
rect 18032 10362 18088 10364
rect 18112 10362 18168 10364
rect 18192 10362 18248 10364
rect 17952 10310 17998 10362
rect 17998 10310 18008 10362
rect 18032 10310 18062 10362
rect 18062 10310 18074 10362
rect 18074 10310 18088 10362
rect 18112 10310 18126 10362
rect 18126 10310 18138 10362
rect 18138 10310 18168 10362
rect 18192 10310 18202 10362
rect 18202 10310 18248 10362
rect 17952 10308 18008 10310
rect 18032 10308 18088 10310
rect 18112 10308 18168 10310
rect 18192 10308 18248 10310
rect 17312 9818 17368 9820
rect 17392 9818 17448 9820
rect 17472 9818 17528 9820
rect 17552 9818 17608 9820
rect 17312 9766 17358 9818
rect 17358 9766 17368 9818
rect 17392 9766 17422 9818
rect 17422 9766 17434 9818
rect 17434 9766 17448 9818
rect 17472 9766 17486 9818
rect 17486 9766 17498 9818
rect 17498 9766 17528 9818
rect 17552 9766 17562 9818
rect 17562 9766 17608 9818
rect 17312 9764 17368 9766
rect 17392 9764 17448 9766
rect 17472 9764 17528 9766
rect 17552 9764 17608 9766
rect 17498 9460 17500 9480
rect 17500 9460 17552 9480
rect 17552 9460 17554 9480
rect 17498 9424 17554 9460
rect 17222 9152 17278 9208
rect 17314 8880 17370 8936
rect 16486 8372 16488 8392
rect 16488 8372 16540 8392
rect 16540 8372 16542 8392
rect 16486 8336 16542 8372
rect 16210 8200 16266 8256
rect 16302 7676 16358 7712
rect 16302 7656 16304 7676
rect 16304 7656 16356 7676
rect 16356 7656 16358 7676
rect 16762 8064 16818 8120
rect 16670 7928 16726 7984
rect 16578 7656 16634 7712
rect 16992 7520 17048 7576
rect 17866 9560 17922 9616
rect 17682 8608 17738 8664
rect 17682 8356 17738 8392
rect 17682 8336 17684 8356
rect 17684 8336 17736 8356
rect 17736 8336 17738 8356
rect 17498 8200 17554 8256
rect 17774 8064 17830 8120
rect 18142 8472 18198 8528
rect 17866 7928 17922 7984
rect 13858 7248 13914 7304
rect 17866 7520 17922 7576
rect 19246 8880 19302 8936
rect 19430 8880 19486 8936
rect 19430 8472 19486 8528
rect 19522 8336 19578 8392
rect 19982 8880 20038 8936
rect 19062 7928 19118 7984
rect 18970 7792 19026 7848
rect 20442 9016 20498 9072
rect 20534 8880 20590 8936
rect 20442 8372 20444 8392
rect 20444 8372 20496 8392
rect 20496 8372 20498 8392
rect 20442 8336 20498 8372
rect 19292 7384 19348 7440
rect 19378 7248 19434 7304
rect 20718 8372 20720 8392
rect 20720 8372 20772 8392
rect 20772 8372 20774 8392
rect 20718 8336 20774 8372
rect 20718 8064 20774 8120
rect 21270 9288 21326 9344
rect 20902 8744 20958 8800
rect 21178 7792 21234 7848
rect 22282 9424 22338 9480
rect 22006 8744 22062 8800
rect 22098 8608 22154 8664
rect 21730 8472 21786 8528
rect 21730 8372 21732 8392
rect 21732 8372 21784 8392
rect 21784 8372 21786 8392
rect 21730 8336 21786 8372
rect 21914 7520 21970 7576
rect 21960 7316 22016 7372
rect 22374 8608 22430 8664
rect 22558 9288 22614 9344
rect 22650 9152 22706 9208
rect 22926 9424 22982 9480
rect 23018 8372 23020 8392
rect 23020 8372 23072 8392
rect 23072 8372 23074 8392
rect 23018 8336 23074 8372
rect 22834 8200 22890 8256
rect 23294 8472 23350 8528
rect 23754 8880 23810 8936
rect 24030 8744 24086 8800
rect 24122 8372 24124 8392
rect 24124 8372 24176 8392
rect 24176 8372 24178 8392
rect 24122 8336 24178 8372
rect 23846 8064 23902 8120
rect 23938 7928 23994 7984
rect 24490 9696 24546 9752
rect 24674 9696 24730 9752
rect 24398 8608 24454 8664
rect 24306 8472 24362 8528
rect 24582 9424 24638 9480
rect 24214 7520 24270 7576
rect 24674 9152 24730 9208
rect 24674 8064 24730 8120
rect 25042 8608 25098 8664
rect 24858 7520 24914 7576
rect 25134 7792 25190 7848
rect 25312 10906 25368 10908
rect 25392 10906 25448 10908
rect 25472 10906 25528 10908
rect 25552 10906 25608 10908
rect 25312 10854 25358 10906
rect 25358 10854 25368 10906
rect 25392 10854 25422 10906
rect 25422 10854 25434 10906
rect 25434 10854 25448 10906
rect 25472 10854 25486 10906
rect 25486 10854 25498 10906
rect 25498 10854 25528 10906
rect 25552 10854 25562 10906
rect 25562 10854 25608 10906
rect 25312 10852 25368 10854
rect 25392 10852 25448 10854
rect 25472 10852 25528 10854
rect 25552 10852 25608 10854
rect 25312 9818 25368 9820
rect 25392 9818 25448 9820
rect 25472 9818 25528 9820
rect 25552 9818 25608 9820
rect 25312 9766 25358 9818
rect 25358 9766 25368 9818
rect 25392 9766 25422 9818
rect 25422 9766 25434 9818
rect 25434 9766 25448 9818
rect 25472 9766 25486 9818
rect 25486 9766 25498 9818
rect 25498 9766 25528 9818
rect 25552 9766 25562 9818
rect 25562 9766 25608 9818
rect 25312 9764 25368 9766
rect 25392 9764 25448 9766
rect 25472 9764 25528 9766
rect 25552 9764 25608 9766
rect 25952 11450 26008 11452
rect 26032 11450 26088 11452
rect 26112 11450 26168 11452
rect 26192 11450 26248 11452
rect 25952 11398 25998 11450
rect 25998 11398 26008 11450
rect 26032 11398 26062 11450
rect 26062 11398 26074 11450
rect 26074 11398 26088 11450
rect 26112 11398 26126 11450
rect 26126 11398 26138 11450
rect 26138 11398 26168 11450
rect 26192 11398 26202 11450
rect 26202 11398 26248 11450
rect 25952 11396 26008 11398
rect 26032 11396 26088 11398
rect 26112 11396 26168 11398
rect 26192 11396 26248 11398
rect 25952 10362 26008 10364
rect 26032 10362 26088 10364
rect 26112 10362 26168 10364
rect 26192 10362 26248 10364
rect 25952 10310 25998 10362
rect 25998 10310 26008 10362
rect 26032 10310 26062 10362
rect 26062 10310 26074 10362
rect 26074 10310 26088 10362
rect 26112 10310 26126 10362
rect 26126 10310 26138 10362
rect 26138 10310 26168 10362
rect 26192 10310 26202 10362
rect 26202 10310 26248 10362
rect 25952 10308 26008 10310
rect 26032 10308 26088 10310
rect 26112 10308 26168 10310
rect 26192 10308 26248 10310
rect 25410 9016 25466 9072
rect 25594 8744 25650 8800
rect 25226 7656 25282 7712
rect 25502 8200 25558 8256
rect 25870 9036 25926 9072
rect 25870 9016 25872 9036
rect 25872 9016 25924 9036
rect 25924 9016 25926 9036
rect 25870 8492 25926 8528
rect 25870 8472 25872 8492
rect 25872 8472 25924 8492
rect 25924 8472 25926 8492
rect 24898 7248 24954 7304
rect 26330 8608 26386 8664
rect 27342 9968 27398 10024
rect 26606 7656 26662 7712
rect 26790 8336 26846 8392
rect 26974 8608 27030 8664
rect 27618 8472 27674 8528
rect 27526 7928 27582 7984
rect 28262 10004 28264 10024
rect 28264 10004 28316 10024
rect 28316 10004 28318 10024
rect 28262 9968 28318 10004
rect 28170 8880 28226 8936
rect 27894 8744 27950 8800
rect 28354 8472 28410 8528
rect 27894 8064 27950 8120
rect 27710 7792 27766 7848
rect 27710 7656 27766 7712
rect 26422 7520 26478 7576
rect 29274 9696 29330 9752
rect 28998 8336 29054 8392
rect 29182 8336 29238 8392
rect 30746 9868 30748 9888
rect 30748 9868 30800 9888
rect 30800 9868 30802 9888
rect 30746 9832 30802 9868
rect 29826 8200 29882 8256
rect 30746 8064 30802 8120
rect 28814 7792 28870 7848
rect 30746 7792 30802 7848
rect 31666 7928 31722 7984
rect 31482 7656 31538 7712
rect 28216 7316 28272 7372
rect 28630 7520 28686 7576
rect 30838 7384 30894 7440
rect 29688 7248 29744 7304
rect 14042 7112 14098 7168
rect 28584 7112 28640 7168
rect 14968 7044 15024 7100
rect 15520 7044 15576 7100
rect 17912 7044 17968 7100
rect 18096 7044 18152 7100
rect 28032 7044 28088 7100
rect 30240 7044 30296 7100
rect 12990 5344 13046 5400
rect 13542 4528 13598 4584
rect 14646 4528 14702 4584
rect 14922 4528 14978 4584
rect 15474 4528 15530 4584
rect 16302 4528 16358 4584
rect 16578 4528 16634 4584
rect 19338 4528 19394 4584
rect 22650 4528 22706 4584
rect 24950 4528 25006 4584
rect 26146 4528 26202 4584
rect 30654 4528 30710 4584
rect 13266 4392 13322 4448
rect 14370 4392 14426 4448
rect 13818 1128 13874 1184
rect 14094 992 14150 1048
rect 15198 4392 15254 4448
rect 15750 1264 15806 1320
rect 16026 1264 16082 1320
rect 17682 4392 17738 4448
rect 18786 4392 18842 4448
rect 17222 4256 17278 4312
rect 16854 2624 16910 2680
rect 17130 2488 17186 2544
rect 17312 2202 17368 2204
rect 17392 2202 17448 2204
rect 17472 2202 17528 2204
rect 17552 2202 17608 2204
rect 17312 2150 17358 2202
rect 17358 2150 17368 2202
rect 17392 2150 17422 2202
rect 17422 2150 17434 2202
rect 17434 2150 17448 2202
rect 17472 2150 17486 2202
rect 17486 2150 17498 2202
rect 17498 2150 17528 2202
rect 17552 2150 17562 2202
rect 17562 2150 17608 2202
rect 17312 2148 17368 2150
rect 17392 2148 17448 2150
rect 17472 2148 17528 2150
rect 17552 2148 17608 2150
rect 17312 1114 17368 1116
rect 17392 1114 17448 1116
rect 17472 1114 17528 1116
rect 17552 1114 17608 1116
rect 17312 1062 17358 1114
rect 17358 1062 17368 1114
rect 17392 1062 17422 1114
rect 17422 1062 17434 1114
rect 17434 1062 17448 1114
rect 17472 1062 17486 1114
rect 17486 1062 17498 1114
rect 17498 1062 17528 1114
rect 17552 1062 17562 1114
rect 17562 1062 17608 1114
rect 17312 1060 17368 1062
rect 17392 1060 17448 1062
rect 17472 1060 17528 1062
rect 17552 1060 17608 1062
rect 18326 4120 18382 4176
rect 17952 1658 18008 1660
rect 18032 1658 18088 1660
rect 18112 1658 18168 1660
rect 18192 1658 18248 1660
rect 17952 1606 17998 1658
rect 17998 1606 18008 1658
rect 18032 1606 18062 1658
rect 18062 1606 18074 1658
rect 18074 1606 18088 1658
rect 18112 1606 18126 1658
rect 18126 1606 18138 1658
rect 18138 1606 18168 1658
rect 18192 1606 18202 1658
rect 18202 1606 18248 1658
rect 17952 1604 18008 1606
rect 18032 1604 18088 1606
rect 18112 1604 18168 1606
rect 18192 1604 18248 1606
rect 17866 856 17922 912
rect 17952 570 18008 572
rect 18032 570 18088 572
rect 18112 570 18168 572
rect 18192 570 18248 572
rect 17952 518 17998 570
rect 17998 518 18008 570
rect 18032 518 18062 570
rect 18062 518 18074 570
rect 18074 518 18088 570
rect 18112 518 18126 570
rect 18126 518 18138 570
rect 18138 518 18168 570
rect 18192 518 18202 570
rect 18202 518 18248 570
rect 17952 516 18008 518
rect 18032 516 18088 518
rect 18112 516 18168 518
rect 18192 516 18248 518
rect 18510 1264 18566 1320
rect 19062 1128 19118 1184
rect 20442 4392 20498 4448
rect 20166 4120 20222 4176
rect 19890 992 19946 1048
rect 19614 720 19670 776
rect 22374 4256 22430 4312
rect 20994 4120 21050 4176
rect 20718 3984 20774 4040
rect 21270 3440 21326 3496
rect 21822 1264 21878 1320
rect 22098 992 22154 1048
rect 22558 1944 22614 2000
rect 23662 1808 23718 1864
rect 22926 1264 22982 1320
rect 23294 1264 23350 1320
rect 25226 4392 25282 4448
rect 25778 4392 25834 4448
rect 25312 2202 25368 2204
rect 25392 2202 25448 2204
rect 25472 2202 25528 2204
rect 25552 2202 25608 2204
rect 25312 2150 25358 2202
rect 25358 2150 25368 2202
rect 25392 2150 25422 2202
rect 25422 2150 25434 2202
rect 25434 2150 25448 2202
rect 25472 2150 25486 2202
rect 25486 2150 25498 2202
rect 25498 2150 25528 2202
rect 25552 2150 25562 2202
rect 25562 2150 25608 2202
rect 25312 2148 25368 2150
rect 25392 2148 25448 2150
rect 25472 2148 25528 2150
rect 25552 2148 25608 2150
rect 25226 1264 25282 1320
rect 25686 1808 25742 1864
rect 28262 4392 28318 4448
rect 27802 3984 27858 4040
rect 25312 1114 25368 1116
rect 25392 1114 25448 1116
rect 25472 1114 25528 1116
rect 25552 1114 25608 1116
rect 25312 1062 25358 1114
rect 25358 1062 25368 1114
rect 25392 1062 25422 1114
rect 25422 1062 25434 1114
rect 25434 1062 25448 1114
rect 25472 1062 25486 1114
rect 25486 1062 25498 1114
rect 25498 1062 25528 1114
rect 25552 1062 25562 1114
rect 25562 1062 25608 1114
rect 25312 1060 25368 1062
rect 25392 1060 25448 1062
rect 25472 1060 25528 1062
rect 25552 1060 25608 1062
rect 25686 856 25742 912
rect 25952 1658 26008 1660
rect 26032 1658 26088 1660
rect 26112 1658 26168 1660
rect 26192 1658 26248 1660
rect 25952 1606 25998 1658
rect 25998 1606 26008 1658
rect 26032 1606 26062 1658
rect 26062 1606 26074 1658
rect 26074 1606 26088 1658
rect 26112 1606 26126 1658
rect 26126 1606 26138 1658
rect 26138 1606 26168 1658
rect 26192 1606 26202 1658
rect 26202 1606 26248 1658
rect 25952 1604 26008 1606
rect 26032 1604 26088 1606
rect 26112 1604 26168 1606
rect 26192 1604 26248 1606
rect 25962 856 26018 912
rect 25952 570 26008 572
rect 26032 570 26088 572
rect 26112 570 26168 572
rect 26192 570 26248 572
rect 25952 518 25998 570
rect 25998 518 26008 570
rect 26032 518 26062 570
rect 26062 518 26074 570
rect 26074 518 26088 570
rect 26112 518 26126 570
rect 26126 518 26138 570
rect 26138 518 26168 570
rect 26192 518 26202 570
rect 26202 518 26248 570
rect 25952 516 26008 518
rect 26032 516 26088 518
rect 26112 516 26168 518
rect 26192 516 26248 518
rect 28446 4120 28502 4176
rect 28722 4120 28778 4176
rect 28078 1264 28134 1320
rect 28538 2624 28594 2680
rect 31022 3984 31078 4040
rect 30378 1264 30434 1320
rect 30746 1300 30748 1320
rect 30748 1300 30800 1320
rect 30800 1300 30802 1320
rect 30746 1264 30802 1300
rect 30930 1264 30986 1320
rect 30654 1128 30710 1184
rect 31666 7656 31722 7712
rect 31942 6296 31998 6352
rect 32310 9832 32366 9888
rect 32218 4528 32274 4584
rect 32954 7792 33010 7848
rect 32862 7656 32918 7712
rect 33952 11450 34008 11452
rect 34032 11450 34088 11452
rect 34112 11450 34168 11452
rect 34192 11450 34248 11452
rect 33952 11398 33998 11450
rect 33998 11398 34008 11450
rect 34032 11398 34062 11450
rect 34062 11398 34074 11450
rect 34074 11398 34088 11450
rect 34112 11398 34126 11450
rect 34126 11398 34138 11450
rect 34138 11398 34168 11450
rect 34192 11398 34202 11450
rect 34202 11398 34248 11450
rect 33952 11396 34008 11398
rect 34032 11396 34088 11398
rect 34112 11396 34168 11398
rect 34192 11396 34248 11398
rect 33312 10906 33368 10908
rect 33392 10906 33448 10908
rect 33472 10906 33528 10908
rect 33552 10906 33608 10908
rect 33312 10854 33358 10906
rect 33358 10854 33368 10906
rect 33392 10854 33422 10906
rect 33422 10854 33434 10906
rect 33434 10854 33448 10906
rect 33472 10854 33486 10906
rect 33486 10854 33498 10906
rect 33498 10854 33528 10906
rect 33552 10854 33562 10906
rect 33562 10854 33608 10906
rect 33312 10852 33368 10854
rect 33392 10852 33448 10854
rect 33472 10852 33528 10854
rect 33552 10852 33608 10854
rect 33312 9818 33368 9820
rect 33392 9818 33448 9820
rect 33472 9818 33528 9820
rect 33552 9818 33608 9820
rect 33312 9766 33358 9818
rect 33358 9766 33368 9818
rect 33392 9766 33422 9818
rect 33422 9766 33434 9818
rect 33434 9766 33448 9818
rect 33472 9766 33486 9818
rect 33486 9766 33498 9818
rect 33498 9766 33528 9818
rect 33552 9766 33562 9818
rect 33562 9766 33608 9818
rect 33312 9764 33368 9766
rect 33392 9764 33448 9766
rect 33472 9764 33528 9766
rect 33552 9764 33608 9766
rect 33138 4120 33194 4176
rect 32678 3032 32734 3088
rect 32954 1264 33010 1320
rect 33230 3712 33286 3768
rect 33414 3848 33470 3904
rect 33230 3032 33286 3088
rect 33598 3440 33654 3496
rect 33312 2202 33368 2204
rect 33392 2202 33448 2204
rect 33472 2202 33528 2204
rect 33552 2202 33608 2204
rect 33312 2150 33358 2202
rect 33358 2150 33368 2202
rect 33392 2150 33422 2202
rect 33422 2150 33434 2202
rect 33434 2150 33448 2202
rect 33472 2150 33486 2202
rect 33486 2150 33498 2202
rect 33498 2150 33528 2202
rect 33552 2150 33562 2202
rect 33562 2150 33608 2202
rect 33312 2148 33368 2150
rect 33392 2148 33448 2150
rect 33472 2148 33528 2150
rect 33552 2148 33608 2150
rect 33322 1964 33378 2000
rect 33322 1944 33324 1964
rect 33324 1944 33376 1964
rect 33376 1944 33378 1964
rect 33312 1114 33368 1116
rect 33392 1114 33448 1116
rect 33472 1114 33528 1116
rect 33552 1114 33608 1116
rect 33312 1062 33358 1114
rect 33358 1062 33368 1114
rect 33392 1062 33422 1114
rect 33422 1062 33434 1114
rect 33434 1062 33448 1114
rect 33472 1062 33486 1114
rect 33486 1062 33498 1114
rect 33498 1062 33528 1114
rect 33552 1062 33562 1114
rect 33562 1062 33608 1114
rect 33312 1060 33368 1062
rect 33392 1060 33448 1062
rect 33472 1060 33528 1062
rect 33552 1060 33608 1062
rect 33952 10362 34008 10364
rect 34032 10362 34088 10364
rect 34112 10362 34168 10364
rect 34192 10362 34248 10364
rect 33952 10310 33998 10362
rect 33998 10310 34008 10362
rect 34032 10310 34062 10362
rect 34062 10310 34074 10362
rect 34074 10310 34088 10362
rect 34112 10310 34126 10362
rect 34126 10310 34138 10362
rect 34138 10310 34168 10362
rect 34192 10310 34202 10362
rect 34202 10310 34248 10362
rect 33952 10308 34008 10310
rect 34032 10308 34088 10310
rect 34112 10308 34168 10310
rect 34192 10308 34248 10310
rect 33952 9274 34008 9276
rect 34032 9274 34088 9276
rect 34112 9274 34168 9276
rect 34192 9274 34248 9276
rect 33952 9222 33998 9274
rect 33998 9222 34008 9274
rect 34032 9222 34062 9274
rect 34062 9222 34074 9274
rect 34074 9222 34088 9274
rect 34112 9222 34126 9274
rect 34126 9222 34138 9274
rect 34138 9222 34168 9274
rect 34192 9222 34202 9274
rect 34202 9222 34248 9274
rect 33952 9220 34008 9222
rect 34032 9220 34088 9222
rect 34112 9220 34168 9222
rect 34192 9220 34248 9222
rect 33952 8186 34008 8188
rect 34032 8186 34088 8188
rect 34112 8186 34168 8188
rect 34192 8186 34248 8188
rect 33952 8134 33998 8186
rect 33998 8134 34008 8186
rect 34032 8134 34062 8186
rect 34062 8134 34074 8186
rect 34074 8134 34088 8186
rect 34112 8134 34126 8186
rect 34126 8134 34138 8186
rect 34138 8134 34168 8186
rect 34192 8134 34202 8186
rect 34202 8134 34248 8186
rect 33952 8132 34008 8134
rect 34032 8132 34088 8134
rect 34112 8132 34168 8134
rect 34192 8132 34248 8134
rect 33952 7098 34008 7100
rect 34032 7098 34088 7100
rect 34112 7098 34168 7100
rect 34192 7098 34248 7100
rect 33952 7046 33998 7098
rect 33998 7046 34008 7098
rect 34032 7046 34062 7098
rect 34062 7046 34074 7098
rect 34074 7046 34088 7098
rect 34112 7046 34126 7098
rect 34126 7046 34138 7098
rect 34138 7046 34168 7098
rect 34192 7046 34202 7098
rect 34202 7046 34248 7098
rect 33952 7044 34008 7046
rect 34032 7044 34088 7046
rect 34112 7044 34168 7046
rect 34192 7044 34248 7046
rect 33952 6010 34008 6012
rect 34032 6010 34088 6012
rect 34112 6010 34168 6012
rect 34192 6010 34248 6012
rect 33952 5958 33998 6010
rect 33998 5958 34008 6010
rect 34032 5958 34062 6010
rect 34062 5958 34074 6010
rect 34074 5958 34088 6010
rect 34112 5958 34126 6010
rect 34126 5958 34138 6010
rect 34138 5958 34168 6010
rect 34192 5958 34202 6010
rect 34202 5958 34248 6010
rect 33952 5956 34008 5958
rect 34032 5956 34088 5958
rect 34112 5956 34168 5958
rect 34192 5956 34248 5958
rect 33952 4922 34008 4924
rect 34032 4922 34088 4924
rect 34112 4922 34168 4924
rect 34192 4922 34248 4924
rect 33952 4870 33998 4922
rect 33998 4870 34008 4922
rect 34032 4870 34062 4922
rect 34062 4870 34074 4922
rect 34074 4870 34088 4922
rect 34112 4870 34126 4922
rect 34126 4870 34138 4922
rect 34138 4870 34168 4922
rect 34192 4870 34202 4922
rect 34202 4870 34248 4922
rect 33952 4868 34008 4870
rect 34032 4868 34088 4870
rect 34112 4868 34168 4870
rect 34192 4868 34248 4870
rect 33952 3834 34008 3836
rect 34032 3834 34088 3836
rect 34112 3834 34168 3836
rect 34192 3834 34248 3836
rect 33952 3782 33998 3834
rect 33998 3782 34008 3834
rect 34032 3782 34062 3834
rect 34062 3782 34074 3834
rect 34074 3782 34088 3834
rect 34112 3782 34126 3834
rect 34126 3782 34138 3834
rect 34138 3782 34168 3834
rect 34192 3782 34202 3834
rect 34202 3782 34248 3834
rect 33952 3780 34008 3782
rect 34032 3780 34088 3782
rect 34112 3780 34168 3782
rect 34192 3780 34248 3782
rect 34150 3596 34206 3632
rect 34150 3576 34152 3596
rect 34152 3576 34204 3596
rect 34204 3576 34206 3596
rect 33782 1672 33838 1728
rect 33952 2746 34008 2748
rect 34032 2746 34088 2748
rect 34112 2746 34168 2748
rect 34192 2746 34248 2748
rect 33952 2694 33998 2746
rect 33998 2694 34008 2746
rect 34032 2694 34062 2746
rect 34062 2694 34074 2746
rect 34074 2694 34088 2746
rect 34112 2694 34126 2746
rect 34126 2694 34138 2746
rect 34138 2694 34168 2746
rect 34192 2694 34202 2746
rect 34202 2694 34248 2746
rect 33952 2692 34008 2694
rect 34032 2692 34088 2694
rect 34112 2692 34168 2694
rect 34192 2692 34248 2694
rect 33966 1844 33968 1864
rect 33968 1844 34020 1864
rect 34020 1844 34022 1864
rect 33966 1808 34022 1844
rect 33952 1658 34008 1660
rect 34032 1658 34088 1660
rect 34112 1658 34168 1660
rect 34192 1658 34248 1660
rect 33952 1606 33998 1658
rect 33998 1606 34008 1658
rect 34032 1606 34062 1658
rect 34062 1606 34074 1658
rect 34074 1606 34088 1658
rect 34112 1606 34126 1658
rect 34126 1606 34138 1658
rect 34138 1606 34168 1658
rect 34192 1606 34202 1658
rect 34202 1606 34248 1658
rect 33952 1604 34008 1606
rect 34032 1604 34088 1606
rect 34112 1604 34168 1606
rect 34192 1604 34248 1606
rect 35070 7248 35126 7304
rect 35162 3440 35218 3496
rect 35070 3032 35126 3088
rect 34886 2896 34942 2952
rect 33952 570 34008 572
rect 34032 570 34088 572
rect 34112 570 34168 572
rect 34192 570 34248 572
rect 33952 518 33998 570
rect 33998 518 34008 570
rect 34032 518 34062 570
rect 34062 518 34074 570
rect 34074 518 34088 570
rect 34112 518 34126 570
rect 34126 518 34138 570
rect 34138 518 34168 570
rect 34192 518 34202 570
rect 34202 518 34248 570
rect 33952 516 34008 518
rect 34032 516 34088 518
rect 34112 516 34168 518
rect 34192 516 34248 518
rect 36266 2760 36322 2816
rect 36266 2488 36322 2544
rect 36266 856 36322 912
rect 36542 2080 36598 2136
rect 36818 3304 36874 3360
rect 36910 2760 36966 2816
rect 36818 2624 36874 2680
rect 36634 1808 36690 1864
rect 37278 3304 37334 3360
rect 37462 3052 37518 3088
rect 37462 3032 37464 3052
rect 37464 3032 37516 3052
rect 37516 3032 37518 3052
rect 37554 2352 37610 2408
rect 37554 2216 37610 2272
rect 38014 3304 38070 3360
rect 38014 2896 38070 2952
rect 38106 2624 38162 2680
rect 38106 2508 38162 2544
rect 38106 2488 38108 2508
rect 38108 2488 38160 2508
rect 38160 2488 38162 2508
rect 38290 2760 38346 2816
rect 38290 2624 38346 2680
rect 41952 11450 42008 11452
rect 42032 11450 42088 11452
rect 42112 11450 42168 11452
rect 42192 11450 42248 11452
rect 41952 11398 41998 11450
rect 41998 11398 42008 11450
rect 42032 11398 42062 11450
rect 42062 11398 42074 11450
rect 42074 11398 42088 11450
rect 42112 11398 42126 11450
rect 42126 11398 42138 11450
rect 42138 11398 42168 11450
rect 42192 11398 42202 11450
rect 42202 11398 42248 11450
rect 41952 11396 42008 11398
rect 42032 11396 42088 11398
rect 42112 11396 42168 11398
rect 42192 11396 42248 11398
rect 41312 10906 41368 10908
rect 41392 10906 41448 10908
rect 41472 10906 41528 10908
rect 41552 10906 41608 10908
rect 41312 10854 41358 10906
rect 41358 10854 41368 10906
rect 41392 10854 41422 10906
rect 41422 10854 41434 10906
rect 41434 10854 41448 10906
rect 41472 10854 41486 10906
rect 41486 10854 41498 10906
rect 41498 10854 41528 10906
rect 41552 10854 41562 10906
rect 41562 10854 41608 10906
rect 41312 10852 41368 10854
rect 41392 10852 41448 10854
rect 41472 10852 41528 10854
rect 41552 10852 41608 10854
rect 41952 10362 42008 10364
rect 42032 10362 42088 10364
rect 42112 10362 42168 10364
rect 42192 10362 42248 10364
rect 41952 10310 41998 10362
rect 41998 10310 42008 10362
rect 42032 10310 42062 10362
rect 42062 10310 42074 10362
rect 42074 10310 42088 10362
rect 42112 10310 42126 10362
rect 42126 10310 42138 10362
rect 42138 10310 42168 10362
rect 42192 10310 42202 10362
rect 42202 10310 42248 10362
rect 41952 10308 42008 10310
rect 42032 10308 42088 10310
rect 42112 10308 42168 10310
rect 42192 10308 42248 10310
rect 41312 9818 41368 9820
rect 41392 9818 41448 9820
rect 41472 9818 41528 9820
rect 41552 9818 41608 9820
rect 41312 9766 41358 9818
rect 41358 9766 41368 9818
rect 41392 9766 41422 9818
rect 41422 9766 41434 9818
rect 41434 9766 41448 9818
rect 41472 9766 41486 9818
rect 41486 9766 41498 9818
rect 41498 9766 41528 9818
rect 41552 9766 41562 9818
rect 41562 9766 41608 9818
rect 41312 9764 41368 9766
rect 41392 9764 41448 9766
rect 41472 9764 41528 9766
rect 41552 9764 41608 9766
rect 38474 2624 38530 2680
rect 38566 2488 38622 2544
rect 38750 2488 38806 2544
rect 39118 2896 39174 2952
rect 39026 2080 39082 2136
rect 38750 1980 38752 2000
rect 38752 1980 38804 2000
rect 38804 1980 38806 2000
rect 38750 1944 38806 1980
rect 38658 1844 38660 1864
rect 38660 1844 38712 1864
rect 38712 1844 38714 1864
rect 38658 1808 38714 1844
rect 38934 1808 38990 1864
rect 38750 1536 38806 1592
rect 39210 1944 39266 2000
rect 39394 2352 39450 2408
rect 39670 2252 39672 2272
rect 39672 2252 39724 2272
rect 39724 2252 39726 2272
rect 39670 2216 39726 2252
rect 39302 1536 39358 1592
rect 38658 720 38714 776
rect 40038 2624 40094 2680
rect 41952 9274 42008 9276
rect 42032 9274 42088 9276
rect 42112 9274 42168 9276
rect 42192 9274 42248 9276
rect 41952 9222 41998 9274
rect 41998 9222 42008 9274
rect 42032 9222 42062 9274
rect 42062 9222 42074 9274
rect 42074 9222 42088 9274
rect 42112 9222 42126 9274
rect 42126 9222 42138 9274
rect 42138 9222 42168 9274
rect 42192 9222 42202 9274
rect 42202 9222 42248 9274
rect 41952 9220 42008 9222
rect 42032 9220 42088 9222
rect 42112 9220 42168 9222
rect 42192 9220 42248 9222
rect 41312 8730 41368 8732
rect 41392 8730 41448 8732
rect 41472 8730 41528 8732
rect 41552 8730 41608 8732
rect 41312 8678 41358 8730
rect 41358 8678 41368 8730
rect 41392 8678 41422 8730
rect 41422 8678 41434 8730
rect 41434 8678 41448 8730
rect 41472 8678 41486 8730
rect 41486 8678 41498 8730
rect 41498 8678 41528 8730
rect 41552 8678 41562 8730
rect 41562 8678 41608 8730
rect 41312 8676 41368 8678
rect 41392 8676 41448 8678
rect 41472 8676 41528 8678
rect 41552 8676 41608 8678
rect 41952 8186 42008 8188
rect 42032 8186 42088 8188
rect 42112 8186 42168 8188
rect 42192 8186 42248 8188
rect 41952 8134 41998 8186
rect 41998 8134 42008 8186
rect 42032 8134 42062 8186
rect 42062 8134 42074 8186
rect 42074 8134 42088 8186
rect 42112 8134 42126 8186
rect 42126 8134 42138 8186
rect 42138 8134 42168 8186
rect 42192 8134 42202 8186
rect 42202 8134 42248 8186
rect 41952 8132 42008 8134
rect 42032 8132 42088 8134
rect 42112 8132 42168 8134
rect 42192 8132 42248 8134
rect 41312 7642 41368 7644
rect 41392 7642 41448 7644
rect 41472 7642 41528 7644
rect 41552 7642 41608 7644
rect 41312 7590 41358 7642
rect 41358 7590 41368 7642
rect 41392 7590 41422 7642
rect 41422 7590 41434 7642
rect 41434 7590 41448 7642
rect 41472 7590 41486 7642
rect 41486 7590 41498 7642
rect 41498 7590 41528 7642
rect 41552 7590 41562 7642
rect 41562 7590 41608 7642
rect 41312 7588 41368 7590
rect 41392 7588 41448 7590
rect 41472 7588 41528 7590
rect 41552 7588 41608 7590
rect 41952 7098 42008 7100
rect 42032 7098 42088 7100
rect 42112 7098 42168 7100
rect 42192 7098 42248 7100
rect 41952 7046 41998 7098
rect 41998 7046 42008 7098
rect 42032 7046 42062 7098
rect 42062 7046 42074 7098
rect 42074 7046 42088 7098
rect 42112 7046 42126 7098
rect 42126 7046 42138 7098
rect 42138 7046 42168 7098
rect 42192 7046 42202 7098
rect 42202 7046 42248 7098
rect 41952 7044 42008 7046
rect 42032 7044 42088 7046
rect 42112 7044 42168 7046
rect 42192 7044 42248 7046
rect 41312 6554 41368 6556
rect 41392 6554 41448 6556
rect 41472 6554 41528 6556
rect 41552 6554 41608 6556
rect 41312 6502 41358 6554
rect 41358 6502 41368 6554
rect 41392 6502 41422 6554
rect 41422 6502 41434 6554
rect 41434 6502 41448 6554
rect 41472 6502 41486 6554
rect 41486 6502 41498 6554
rect 41498 6502 41528 6554
rect 41552 6502 41562 6554
rect 41562 6502 41608 6554
rect 41312 6500 41368 6502
rect 41392 6500 41448 6502
rect 41472 6500 41528 6502
rect 41552 6500 41608 6502
rect 41952 6010 42008 6012
rect 42032 6010 42088 6012
rect 42112 6010 42168 6012
rect 42192 6010 42248 6012
rect 41952 5958 41998 6010
rect 41998 5958 42008 6010
rect 42032 5958 42062 6010
rect 42062 5958 42074 6010
rect 42074 5958 42088 6010
rect 42112 5958 42126 6010
rect 42126 5958 42138 6010
rect 42138 5958 42168 6010
rect 42192 5958 42202 6010
rect 42202 5958 42248 6010
rect 41952 5956 42008 5958
rect 42032 5956 42088 5958
rect 42112 5956 42168 5958
rect 42192 5956 42248 5958
rect 41312 5466 41368 5468
rect 41392 5466 41448 5468
rect 41472 5466 41528 5468
rect 41552 5466 41608 5468
rect 41312 5414 41358 5466
rect 41358 5414 41368 5466
rect 41392 5414 41422 5466
rect 41422 5414 41434 5466
rect 41434 5414 41448 5466
rect 41472 5414 41486 5466
rect 41486 5414 41498 5466
rect 41498 5414 41528 5466
rect 41552 5414 41562 5466
rect 41562 5414 41608 5466
rect 41312 5412 41368 5414
rect 41392 5412 41448 5414
rect 41472 5412 41528 5414
rect 41552 5412 41608 5414
rect 41952 4922 42008 4924
rect 42032 4922 42088 4924
rect 42112 4922 42168 4924
rect 42192 4922 42248 4924
rect 41952 4870 41998 4922
rect 41998 4870 42008 4922
rect 42032 4870 42062 4922
rect 42062 4870 42074 4922
rect 42074 4870 42088 4922
rect 42112 4870 42126 4922
rect 42126 4870 42138 4922
rect 42138 4870 42168 4922
rect 42192 4870 42202 4922
rect 42202 4870 42248 4922
rect 41952 4868 42008 4870
rect 42032 4868 42088 4870
rect 42112 4868 42168 4870
rect 42192 4868 42248 4870
rect 41312 4378 41368 4380
rect 41392 4378 41448 4380
rect 41472 4378 41528 4380
rect 41552 4378 41608 4380
rect 41312 4326 41358 4378
rect 41358 4326 41368 4378
rect 41392 4326 41422 4378
rect 41422 4326 41434 4378
rect 41434 4326 41448 4378
rect 41472 4326 41486 4378
rect 41486 4326 41498 4378
rect 41498 4326 41528 4378
rect 41552 4326 41562 4378
rect 41562 4326 41608 4378
rect 41312 4324 41368 4326
rect 41392 4324 41448 4326
rect 41472 4324 41528 4326
rect 41552 4324 41608 4326
rect 41952 3834 42008 3836
rect 42032 3834 42088 3836
rect 42112 3834 42168 3836
rect 42192 3834 42248 3836
rect 41952 3782 41998 3834
rect 41998 3782 42008 3834
rect 42032 3782 42062 3834
rect 42062 3782 42074 3834
rect 42074 3782 42088 3834
rect 42112 3782 42126 3834
rect 42126 3782 42138 3834
rect 42138 3782 42168 3834
rect 42192 3782 42202 3834
rect 42202 3782 42248 3834
rect 41952 3780 42008 3782
rect 42032 3780 42088 3782
rect 42112 3780 42168 3782
rect 42192 3780 42248 3782
rect 41312 3290 41368 3292
rect 41392 3290 41448 3292
rect 41472 3290 41528 3292
rect 41552 3290 41608 3292
rect 41312 3238 41358 3290
rect 41358 3238 41368 3290
rect 41392 3238 41422 3290
rect 41422 3238 41434 3290
rect 41434 3238 41448 3290
rect 41472 3238 41486 3290
rect 41486 3238 41498 3290
rect 41498 3238 41528 3290
rect 41552 3238 41562 3290
rect 41562 3238 41608 3290
rect 41312 3236 41368 3238
rect 41392 3236 41448 3238
rect 41472 3236 41528 3238
rect 41552 3236 41608 3238
rect 41952 2746 42008 2748
rect 42032 2746 42088 2748
rect 42112 2746 42168 2748
rect 42192 2746 42248 2748
rect 41952 2694 41998 2746
rect 41998 2694 42008 2746
rect 42032 2694 42062 2746
rect 42062 2694 42074 2746
rect 42074 2694 42088 2746
rect 42112 2694 42126 2746
rect 42126 2694 42138 2746
rect 42138 2694 42168 2746
rect 42192 2694 42202 2746
rect 42202 2694 42248 2746
rect 41952 2692 42008 2694
rect 42032 2692 42088 2694
rect 42112 2692 42168 2694
rect 42192 2692 42248 2694
rect 40406 1536 40462 1592
rect 41312 2202 41368 2204
rect 41392 2202 41448 2204
rect 41472 2202 41528 2204
rect 41552 2202 41608 2204
rect 41312 2150 41358 2202
rect 41358 2150 41368 2202
rect 41392 2150 41422 2202
rect 41422 2150 41434 2202
rect 41434 2150 41448 2202
rect 41472 2150 41486 2202
rect 41486 2150 41498 2202
rect 41498 2150 41528 2202
rect 41552 2150 41562 2202
rect 41562 2150 41608 2202
rect 41312 2148 41368 2150
rect 41392 2148 41448 2150
rect 41472 2148 41528 2150
rect 41552 2148 41608 2150
rect 40498 756 40500 776
rect 40500 756 40552 776
rect 40552 756 40554 776
rect 40498 720 40554 756
rect 40406 620 40408 640
rect 40408 620 40460 640
rect 40460 620 40462 640
rect 40406 584 40462 620
rect 41952 1658 42008 1660
rect 42032 1658 42088 1660
rect 42112 1658 42168 1660
rect 42192 1658 42248 1660
rect 41952 1606 41998 1658
rect 41998 1606 42008 1658
rect 42032 1606 42062 1658
rect 42062 1606 42074 1658
rect 42074 1606 42088 1658
rect 42112 1606 42126 1658
rect 42126 1606 42138 1658
rect 42138 1606 42168 1658
rect 42192 1606 42202 1658
rect 42202 1606 42248 1658
rect 41952 1604 42008 1606
rect 42032 1604 42088 1606
rect 42112 1604 42168 1606
rect 42192 1604 42248 1606
rect 41312 1114 41368 1116
rect 41392 1114 41448 1116
rect 41472 1114 41528 1116
rect 41552 1114 41608 1116
rect 41312 1062 41358 1114
rect 41358 1062 41368 1114
rect 41392 1062 41422 1114
rect 41422 1062 41434 1114
rect 41434 1062 41448 1114
rect 41472 1062 41486 1114
rect 41486 1062 41498 1114
rect 41498 1062 41528 1114
rect 41552 1062 41562 1114
rect 41562 1062 41608 1114
rect 41312 1060 41368 1062
rect 41392 1060 41448 1062
rect 41472 1060 41528 1062
rect 41552 1060 41608 1062
rect 41786 856 41842 912
rect 42338 756 42340 776
rect 42340 756 42392 776
rect 42392 756 42394 776
rect 42338 720 42394 756
rect 41326 584 41382 640
rect 41952 570 42008 572
rect 42032 570 42088 572
rect 42112 570 42168 572
rect 42192 570 42248 572
rect 41952 518 41998 570
rect 41998 518 42008 570
rect 42032 518 42062 570
rect 42062 518 42074 570
rect 42074 518 42088 570
rect 42112 518 42126 570
rect 42126 518 42138 570
rect 42138 518 42168 570
rect 42192 518 42202 570
rect 42202 518 42248 570
rect 41952 516 42008 518
rect 42032 516 42088 518
rect 42112 516 42168 518
rect 42192 516 42248 518
<< metal3 >>
rect 1942 11456 2258 11457
rect 1942 11392 1948 11456
rect 2012 11392 2028 11456
rect 2092 11392 2108 11456
rect 2172 11392 2188 11456
rect 2252 11392 2258 11456
rect 1942 11391 2258 11392
rect 9942 11456 10258 11457
rect 9942 11392 9948 11456
rect 10012 11392 10028 11456
rect 10092 11392 10108 11456
rect 10172 11392 10188 11456
rect 10252 11392 10258 11456
rect 9942 11391 10258 11392
rect 17942 11456 18258 11457
rect 17942 11392 17948 11456
rect 18012 11392 18028 11456
rect 18092 11392 18108 11456
rect 18172 11392 18188 11456
rect 18252 11392 18258 11456
rect 17942 11391 18258 11392
rect 25942 11456 26258 11457
rect 25942 11392 25948 11456
rect 26012 11392 26028 11456
rect 26092 11392 26108 11456
rect 26172 11392 26188 11456
rect 26252 11392 26258 11456
rect 25942 11391 26258 11392
rect 33942 11456 34258 11457
rect 33942 11392 33948 11456
rect 34012 11392 34028 11456
rect 34092 11392 34108 11456
rect 34172 11392 34188 11456
rect 34252 11392 34258 11456
rect 33942 11391 34258 11392
rect 41942 11456 42258 11457
rect 41942 11392 41948 11456
rect 42012 11392 42028 11456
rect 42092 11392 42108 11456
rect 42172 11392 42188 11456
rect 42252 11392 42258 11456
rect 41942 11391 42258 11392
rect 1302 10912 1618 10913
rect 1302 10848 1308 10912
rect 1372 10848 1388 10912
rect 1452 10848 1468 10912
rect 1532 10848 1548 10912
rect 1612 10848 1618 10912
rect 1302 10847 1618 10848
rect 9302 10912 9618 10913
rect 9302 10848 9308 10912
rect 9372 10848 9388 10912
rect 9452 10848 9468 10912
rect 9532 10848 9548 10912
rect 9612 10848 9618 10912
rect 9302 10847 9618 10848
rect 17302 10912 17618 10913
rect 17302 10848 17308 10912
rect 17372 10848 17388 10912
rect 17452 10848 17468 10912
rect 17532 10848 17548 10912
rect 17612 10848 17618 10912
rect 17302 10847 17618 10848
rect 25302 10912 25618 10913
rect 25302 10848 25308 10912
rect 25372 10848 25388 10912
rect 25452 10848 25468 10912
rect 25532 10848 25548 10912
rect 25612 10848 25618 10912
rect 25302 10847 25618 10848
rect 33302 10912 33618 10913
rect 33302 10848 33308 10912
rect 33372 10848 33388 10912
rect 33452 10848 33468 10912
rect 33532 10848 33548 10912
rect 33612 10848 33618 10912
rect 33302 10847 33618 10848
rect 41302 10912 41618 10913
rect 41302 10848 41308 10912
rect 41372 10848 41388 10912
rect 41452 10848 41468 10912
rect 41532 10848 41548 10912
rect 41612 10848 41618 10912
rect 41302 10847 41618 10848
rect 1942 10368 2258 10369
rect 1942 10304 1948 10368
rect 2012 10304 2028 10368
rect 2092 10304 2108 10368
rect 2172 10304 2188 10368
rect 2252 10304 2258 10368
rect 1942 10303 2258 10304
rect 9942 10368 10258 10369
rect 9942 10304 9948 10368
rect 10012 10304 10028 10368
rect 10092 10304 10108 10368
rect 10172 10304 10188 10368
rect 10252 10304 10258 10368
rect 9942 10303 10258 10304
rect 17942 10368 18258 10369
rect 17942 10304 17948 10368
rect 18012 10304 18028 10368
rect 18092 10304 18108 10368
rect 18172 10304 18188 10368
rect 18252 10304 18258 10368
rect 17942 10303 18258 10304
rect 25942 10368 26258 10369
rect 25942 10304 25948 10368
rect 26012 10304 26028 10368
rect 26092 10304 26108 10368
rect 26172 10304 26188 10368
rect 26252 10304 26258 10368
rect 25942 10303 26258 10304
rect 33942 10368 34258 10369
rect 33942 10304 33948 10368
rect 34012 10304 34028 10368
rect 34092 10304 34108 10368
rect 34172 10304 34188 10368
rect 34252 10304 34258 10368
rect 33942 10303 34258 10304
rect 41942 10368 42258 10369
rect 41942 10304 41948 10368
rect 42012 10304 42028 10368
rect 42092 10304 42108 10368
rect 42172 10304 42188 10368
rect 42252 10304 42258 10368
rect 41942 10303 42258 10304
rect 27337 10026 27403 10029
rect 28257 10026 28323 10029
rect 27337 10024 28323 10026
rect 27337 9968 27342 10024
rect 27398 9968 28262 10024
rect 28318 9968 28323 10024
rect 27337 9966 28323 9968
rect 27337 9963 27403 9966
rect 28257 9963 28323 9966
rect 30741 9890 30807 9893
rect 32305 9890 32371 9893
rect 30741 9888 32371 9890
rect 30741 9832 30746 9888
rect 30802 9832 32310 9888
rect 32366 9832 32371 9888
rect 30741 9830 32371 9832
rect 30741 9827 30807 9830
rect 32305 9827 32371 9830
rect 1302 9824 1618 9825
rect 1302 9760 1308 9824
rect 1372 9760 1388 9824
rect 1452 9760 1468 9824
rect 1532 9760 1548 9824
rect 1612 9760 1618 9824
rect 1302 9759 1618 9760
rect 9302 9824 9618 9825
rect 9302 9760 9308 9824
rect 9372 9760 9388 9824
rect 9452 9760 9468 9824
rect 9532 9760 9548 9824
rect 9612 9760 9618 9824
rect 9302 9759 9618 9760
rect 17302 9824 17618 9825
rect 17302 9760 17308 9824
rect 17372 9760 17388 9824
rect 17452 9760 17468 9824
rect 17532 9760 17548 9824
rect 17612 9760 17618 9824
rect 17302 9759 17618 9760
rect 25302 9824 25618 9825
rect 25302 9760 25308 9824
rect 25372 9760 25388 9824
rect 25452 9760 25468 9824
rect 25532 9760 25548 9824
rect 25612 9760 25618 9824
rect 25302 9759 25618 9760
rect 33302 9824 33618 9825
rect 33302 9760 33308 9824
rect 33372 9760 33388 9824
rect 33452 9760 33468 9824
rect 33532 9760 33548 9824
rect 33612 9760 33618 9824
rect 33302 9759 33618 9760
rect 41302 9824 41618 9825
rect 41302 9760 41308 9824
rect 41372 9760 41388 9824
rect 41452 9760 41468 9824
rect 41532 9760 41548 9824
rect 41612 9760 41618 9824
rect 41302 9759 41618 9760
rect 24485 9756 24551 9757
rect 24669 9756 24735 9757
rect 24485 9754 24532 9756
rect 24440 9752 24532 9754
rect 24440 9696 24490 9752
rect 24440 9694 24532 9696
rect 24485 9692 24532 9694
rect 24596 9692 24602 9756
rect 24669 9752 24716 9756
rect 24780 9754 24786 9756
rect 29269 9754 29335 9757
rect 32990 9754 32996 9756
rect 24669 9696 24674 9752
rect 24669 9692 24716 9696
rect 24780 9694 24826 9754
rect 29269 9752 32996 9754
rect 29269 9696 29274 9752
rect 29330 9696 32996 9752
rect 29269 9694 32996 9696
rect 24780 9692 24786 9694
rect 24485 9691 24551 9692
rect 24669 9691 24735 9692
rect 29269 9691 29335 9694
rect 32990 9692 32996 9694
rect 33060 9692 33066 9756
rect 13997 9618 14063 9621
rect 17861 9618 17927 9621
rect 13997 9616 17927 9618
rect 13997 9560 14002 9616
rect 14058 9560 17866 9616
rect 17922 9560 17927 9616
rect 13997 9558 17927 9560
rect 13997 9555 14063 9558
rect 17861 9555 17927 9558
rect 14089 9484 14155 9485
rect 14038 9420 14044 9484
rect 14108 9482 14155 9484
rect 14108 9480 14200 9482
rect 14150 9424 14200 9480
rect 14108 9422 14200 9424
rect 14108 9420 14155 9422
rect 14590 9420 14596 9484
rect 14660 9482 14666 9484
rect 16205 9482 16271 9485
rect 14660 9480 16271 9482
rect 14660 9424 16210 9480
rect 16266 9424 16271 9480
rect 14660 9422 16271 9424
rect 14660 9420 14666 9422
rect 14089 9419 14155 9420
rect 16205 9419 16271 9422
rect 17493 9482 17559 9485
rect 22277 9482 22343 9485
rect 17493 9480 22343 9482
rect 17493 9424 17498 9480
rect 17554 9424 22282 9480
rect 22338 9424 22343 9480
rect 17493 9422 22343 9424
rect 17493 9419 17559 9422
rect 22277 9419 22343 9422
rect 22921 9482 22987 9485
rect 24577 9482 24643 9485
rect 22921 9480 24643 9482
rect 22921 9424 22926 9480
rect 22982 9424 24582 9480
rect 24638 9424 24643 9480
rect 22921 9422 24643 9424
rect 22921 9419 22987 9422
rect 24577 9419 24643 9422
rect 15653 9346 15719 9349
rect 14230 9344 15719 9346
rect 14230 9288 15658 9344
rect 15714 9288 15719 9344
rect 14230 9286 15719 9288
rect 1942 9280 2258 9281
rect 1942 9216 1948 9280
rect 2012 9216 2028 9280
rect 2092 9216 2108 9280
rect 2172 9216 2188 9280
rect 2252 9216 2258 9280
rect 1942 9215 2258 9216
rect 9942 9280 10258 9281
rect 9942 9216 9948 9280
rect 10012 9216 10028 9280
rect 10092 9216 10108 9280
rect 10172 9216 10188 9280
rect 10252 9216 10258 9280
rect 9942 9215 10258 9216
rect 10869 9210 10935 9213
rect 14230 9210 14290 9286
rect 15653 9283 15719 9286
rect 16021 9346 16087 9349
rect 21265 9346 21331 9349
rect 16021 9344 21331 9346
rect 16021 9288 16026 9344
rect 16082 9288 21270 9344
rect 21326 9288 21331 9344
rect 16021 9286 21331 9288
rect 16021 9283 16087 9286
rect 21265 9283 21331 9286
rect 22318 9284 22324 9348
rect 22388 9346 22394 9348
rect 22553 9346 22619 9349
rect 22388 9344 22619 9346
rect 22388 9288 22558 9344
rect 22614 9288 22619 9344
rect 22388 9286 22619 9288
rect 22388 9284 22394 9286
rect 22553 9283 22619 9286
rect 33942 9280 34258 9281
rect 33942 9216 33948 9280
rect 34012 9216 34028 9280
rect 34092 9216 34108 9280
rect 34172 9216 34188 9280
rect 34252 9216 34258 9280
rect 33942 9215 34258 9216
rect 41942 9280 42258 9281
rect 41942 9216 41948 9280
rect 42012 9216 42028 9280
rect 42092 9216 42108 9280
rect 42172 9216 42188 9280
rect 42252 9216 42258 9280
rect 41942 9215 42258 9216
rect 10869 9208 14290 9210
rect 10869 9152 10874 9208
rect 10930 9152 14290 9208
rect 10869 9150 14290 9152
rect 14365 9210 14431 9213
rect 16481 9210 16547 9213
rect 14365 9208 16547 9210
rect 14365 9152 14370 9208
rect 14426 9152 16486 9208
rect 16542 9152 16547 9208
rect 14365 9150 16547 9152
rect 10869 9147 10935 9150
rect 14365 9147 14431 9150
rect 16481 9147 16547 9150
rect 17217 9210 17283 9213
rect 22645 9210 22711 9213
rect 17217 9208 22711 9210
rect 17217 9152 17222 9208
rect 17278 9152 22650 9208
rect 22706 9152 22711 9208
rect 17217 9150 22711 9152
rect 17217 9147 17283 9150
rect 22645 9147 22711 9150
rect 23238 9148 23244 9212
rect 23308 9210 23314 9212
rect 24669 9210 24735 9213
rect 23308 9208 24735 9210
rect 23308 9152 24674 9208
rect 24730 9152 24735 9208
rect 23308 9150 24735 9152
rect 23308 9148 23314 9150
rect 24669 9147 24735 9150
rect 10685 9074 10751 9077
rect 13997 9074 14063 9077
rect 10685 9072 14063 9074
rect 10685 9016 10690 9072
rect 10746 9016 14002 9072
rect 14058 9016 14063 9072
rect 10685 9014 14063 9016
rect 10685 9011 10751 9014
rect 13997 9011 14063 9014
rect 14406 9012 14412 9076
rect 14476 9074 14482 9076
rect 14733 9074 14799 9077
rect 14476 9072 14799 9074
rect 14476 9016 14738 9072
rect 14794 9016 14799 9072
rect 14476 9014 14799 9016
rect 14476 9012 14482 9014
rect 14733 9011 14799 9014
rect 14917 9074 14983 9077
rect 20437 9074 20503 9077
rect 14917 9072 20503 9074
rect 14917 9016 14922 9072
rect 14978 9016 20442 9072
rect 20498 9016 20503 9072
rect 14917 9014 20503 9016
rect 14917 9011 14983 9014
rect 20437 9011 20503 9014
rect 22502 9012 22508 9076
rect 22572 9074 22578 9076
rect 25405 9074 25471 9077
rect 25865 9074 25931 9077
rect 22572 9072 25931 9074
rect 22572 9016 25410 9072
rect 25466 9016 25870 9072
rect 25926 9016 25931 9072
rect 22572 9014 25931 9016
rect 22572 9012 22578 9014
rect 25405 9011 25471 9014
rect 25865 9011 25931 9014
rect 13670 8876 13676 8940
rect 13740 8938 13746 8940
rect 14641 8938 14707 8941
rect 13740 8936 14707 8938
rect 13740 8880 14646 8936
rect 14702 8880 14707 8936
rect 13740 8878 14707 8880
rect 13740 8876 13746 8878
rect 14641 8875 14707 8878
rect 15837 8938 15903 8941
rect 16062 8938 16068 8940
rect 15837 8936 16068 8938
rect 15837 8880 15842 8936
rect 15898 8880 16068 8936
rect 15837 8878 16068 8880
rect 15837 8875 15903 8878
rect 16062 8876 16068 8878
rect 16132 8876 16138 8940
rect 16430 8876 16436 8940
rect 16500 8938 16506 8940
rect 17033 8938 17099 8941
rect 17309 8938 17375 8941
rect 16500 8936 17375 8938
rect 16500 8880 17038 8936
rect 17094 8880 17314 8936
rect 17370 8880 17375 8936
rect 16500 8878 17375 8880
rect 16500 8876 16506 8878
rect 17033 8875 17099 8878
rect 17309 8875 17375 8878
rect 19006 8876 19012 8940
rect 19076 8938 19082 8940
rect 19241 8938 19307 8941
rect 19076 8936 19307 8938
rect 19076 8880 19246 8936
rect 19302 8880 19307 8936
rect 19076 8878 19307 8880
rect 19076 8876 19082 8878
rect 19241 8875 19307 8878
rect 19425 8938 19491 8941
rect 19977 8940 20043 8941
rect 19742 8938 19748 8940
rect 19425 8936 19748 8938
rect 19425 8880 19430 8936
rect 19486 8880 19748 8936
rect 19425 8878 19748 8880
rect 19425 8875 19491 8878
rect 19742 8876 19748 8878
rect 19812 8876 19818 8940
rect 19926 8876 19932 8940
rect 19996 8938 20043 8940
rect 19996 8936 20088 8938
rect 20038 8880 20088 8936
rect 19996 8878 20088 8880
rect 19996 8876 20043 8878
rect 20294 8876 20300 8940
rect 20364 8938 20370 8940
rect 20529 8938 20595 8941
rect 20364 8936 20595 8938
rect 20364 8880 20534 8936
rect 20590 8880 20595 8936
rect 20364 8878 20595 8880
rect 20364 8876 20370 8878
rect 19977 8875 20043 8876
rect 20529 8875 20595 8878
rect 23606 8876 23612 8940
rect 23676 8938 23682 8940
rect 23749 8938 23815 8941
rect 23676 8936 23815 8938
rect 23676 8880 23754 8936
rect 23810 8880 23815 8936
rect 23676 8878 23815 8880
rect 23676 8876 23682 8878
rect 23749 8875 23815 8878
rect 28165 8938 28231 8941
rect 30782 8938 30788 8940
rect 28165 8936 30788 8938
rect 28165 8880 28170 8936
rect 28226 8880 30788 8936
rect 28165 8878 30788 8880
rect 28165 8875 28231 8878
rect 30782 8876 30788 8878
rect 30852 8876 30858 8940
rect 9765 8802 9831 8805
rect 10542 8802 10548 8804
rect 9765 8800 10548 8802
rect 9765 8744 9770 8800
rect 9826 8744 10548 8800
rect 9765 8742 10548 8744
rect 9765 8739 9831 8742
rect 10542 8740 10548 8742
rect 10612 8740 10618 8804
rect 15694 8740 15700 8804
rect 15764 8802 15770 8804
rect 16665 8802 16731 8805
rect 20897 8802 20963 8805
rect 15764 8800 16731 8802
rect 15764 8744 16670 8800
rect 16726 8744 16731 8800
rect 15764 8742 16731 8744
rect 15764 8740 15770 8742
rect 16665 8739 16731 8742
rect 16852 8800 20963 8802
rect 16852 8744 20902 8800
rect 20958 8744 20963 8800
rect 16852 8742 20963 8744
rect 1302 8736 1618 8737
rect 1302 8672 1308 8736
rect 1372 8672 1388 8736
rect 1452 8672 1468 8736
rect 1532 8672 1548 8736
rect 1612 8672 1618 8736
rect 1302 8671 1618 8672
rect 9302 8736 9618 8737
rect 9302 8672 9308 8736
rect 9372 8672 9388 8736
rect 9452 8672 9468 8736
rect 9532 8672 9548 8736
rect 9612 8672 9618 8736
rect 9302 8671 9618 8672
rect 9806 8604 9812 8668
rect 9876 8666 9882 8668
rect 10358 8666 10364 8668
rect 9876 8606 10364 8666
rect 9876 8604 9882 8606
rect 10358 8604 10364 8606
rect 10428 8604 10434 8668
rect 12617 8666 12683 8669
rect 15101 8666 15167 8669
rect 12617 8664 15167 8666
rect 12617 8608 12622 8664
rect 12678 8608 15106 8664
rect 15162 8608 15167 8664
rect 12617 8606 15167 8608
rect 12617 8603 12683 8606
rect 15101 8603 15167 8606
rect 15510 8604 15516 8668
rect 15580 8666 15586 8668
rect 16573 8666 16639 8669
rect 15580 8664 16639 8666
rect 15580 8608 16578 8664
rect 16634 8608 16639 8664
rect 15580 8606 16639 8608
rect 15580 8604 15586 8606
rect 16573 8603 16639 8606
rect 7373 8530 7439 8533
rect 15653 8530 15719 8533
rect 7373 8528 15719 8530
rect 7373 8472 7378 8528
rect 7434 8472 15658 8528
rect 15714 8472 15719 8528
rect 7373 8470 15719 8472
rect 7373 8467 7439 8470
rect 15653 8467 15719 8470
rect 15929 8530 15995 8533
rect 16852 8530 16912 8742
rect 20897 8739 20963 8742
rect 22001 8802 22067 8805
rect 24025 8802 24091 8805
rect 25589 8802 25655 8805
rect 22001 8800 24091 8802
rect 22001 8744 22006 8800
rect 22062 8744 24030 8800
rect 24086 8744 24091 8800
rect 22001 8742 24091 8744
rect 22001 8739 22067 8742
rect 24025 8739 24091 8742
rect 24212 8800 25655 8802
rect 24212 8744 25594 8800
rect 25650 8744 25655 8800
rect 24212 8742 25655 8744
rect 17677 8666 17743 8669
rect 22093 8666 22159 8669
rect 17677 8664 22159 8666
rect 17677 8608 17682 8664
rect 17738 8608 22098 8664
rect 22154 8608 22159 8664
rect 17677 8606 22159 8608
rect 17677 8603 17743 8606
rect 22093 8603 22159 8606
rect 22369 8666 22435 8669
rect 24212 8666 24272 8742
rect 25589 8739 25655 8742
rect 27889 8802 27955 8805
rect 30414 8802 30420 8804
rect 27889 8800 30420 8802
rect 27889 8744 27894 8800
rect 27950 8744 30420 8800
rect 27889 8742 30420 8744
rect 27889 8739 27955 8742
rect 30414 8740 30420 8742
rect 30484 8740 30490 8804
rect 41302 8736 41618 8737
rect 41302 8672 41308 8736
rect 41372 8672 41388 8736
rect 41452 8672 41468 8736
rect 41532 8672 41548 8736
rect 41612 8672 41618 8736
rect 41302 8671 41618 8672
rect 22369 8664 24272 8666
rect 22369 8608 22374 8664
rect 22430 8608 24272 8664
rect 22369 8606 24272 8608
rect 24393 8666 24459 8669
rect 25037 8666 25103 8669
rect 26325 8666 26391 8669
rect 24393 8664 26391 8666
rect 24393 8608 24398 8664
rect 24454 8608 25042 8664
rect 25098 8608 26330 8664
rect 26386 8608 26391 8664
rect 24393 8606 26391 8608
rect 22369 8603 22435 8606
rect 24393 8603 24459 8606
rect 25037 8603 25103 8606
rect 26325 8603 26391 8606
rect 26969 8666 27035 8669
rect 28390 8666 28396 8668
rect 26969 8664 28396 8666
rect 26969 8608 26974 8664
rect 27030 8608 28396 8664
rect 26969 8606 28396 8608
rect 26969 8603 27035 8606
rect 28390 8604 28396 8606
rect 28460 8604 28466 8668
rect 15929 8528 16912 8530
rect 15929 8472 15934 8528
rect 15990 8472 16912 8528
rect 15929 8470 16912 8472
rect 15929 8467 15995 8470
rect 16982 8468 16988 8532
rect 17052 8530 17058 8532
rect 18137 8530 18203 8533
rect 17052 8528 18203 8530
rect 17052 8472 18142 8528
rect 18198 8472 18203 8528
rect 17052 8470 18203 8472
rect 17052 8468 17058 8470
rect 18137 8467 18203 8470
rect 19425 8530 19491 8533
rect 20846 8530 20852 8532
rect 19425 8528 20852 8530
rect 19425 8472 19430 8528
rect 19486 8472 20852 8528
rect 19425 8470 20852 8472
rect 19425 8467 19491 8470
rect 20846 8468 20852 8470
rect 20916 8468 20922 8532
rect 21398 8468 21404 8532
rect 21468 8530 21474 8532
rect 21725 8530 21791 8533
rect 21468 8528 21791 8530
rect 21468 8472 21730 8528
rect 21786 8472 21791 8528
rect 21468 8470 21791 8472
rect 21468 8468 21474 8470
rect 21725 8467 21791 8470
rect 23289 8530 23355 8533
rect 24301 8530 24367 8533
rect 25865 8530 25931 8533
rect 23289 8528 25931 8530
rect 23289 8472 23294 8528
rect 23350 8472 24306 8528
rect 24362 8472 25870 8528
rect 25926 8472 25931 8528
rect 23289 8470 25931 8472
rect 23289 8467 23355 8470
rect 24301 8467 24367 8470
rect 25865 8467 25931 8470
rect 27613 8530 27679 8533
rect 27838 8530 27844 8532
rect 27613 8528 27844 8530
rect 27613 8472 27618 8528
rect 27674 8472 27844 8528
rect 27613 8470 27844 8472
rect 27613 8467 27679 8470
rect 27838 8468 27844 8470
rect 27908 8468 27914 8532
rect 28349 8530 28415 8533
rect 30966 8530 30972 8532
rect 28349 8528 30972 8530
rect 28349 8472 28354 8528
rect 28410 8472 30972 8528
rect 28349 8470 30972 8472
rect 28349 8467 28415 8470
rect 30966 8468 30972 8470
rect 31036 8468 31042 8532
rect 10685 8394 10751 8397
rect 13169 8394 13235 8397
rect 9814 8334 10426 8394
rect 5165 8258 5231 8261
rect 9814 8258 9874 8334
rect 5165 8256 9874 8258
rect 5165 8200 5170 8256
rect 5226 8200 9874 8256
rect 5165 8198 9874 8200
rect 5165 8195 5231 8198
rect 1942 8192 2258 8193
rect 1942 8128 1948 8192
rect 2012 8128 2028 8192
rect 2092 8128 2108 8192
rect 2172 8128 2188 8192
rect 2252 8128 2258 8192
rect 1942 8127 2258 8128
rect 9942 8192 10258 8193
rect 9942 8128 9948 8192
rect 10012 8128 10028 8192
rect 10092 8128 10108 8192
rect 10172 8128 10188 8192
rect 10252 8128 10258 8192
rect 9942 8127 10258 8128
rect 9673 8122 9739 8125
rect 9806 8122 9812 8124
rect 9673 8120 9812 8122
rect 9673 8064 9678 8120
rect 9734 8064 9812 8120
rect 9673 8062 9812 8064
rect 9673 8059 9739 8062
rect 9806 8060 9812 8062
rect 9876 8060 9882 8124
rect 10366 8122 10426 8334
rect 10685 8392 13235 8394
rect 10685 8336 10690 8392
rect 10746 8336 13174 8392
rect 13230 8336 13235 8392
rect 10685 8334 13235 8336
rect 10685 8331 10751 8334
rect 13169 8331 13235 8334
rect 13302 8332 13308 8396
rect 13372 8394 13378 8396
rect 13445 8394 13511 8397
rect 13372 8392 13511 8394
rect 13372 8336 13450 8392
rect 13506 8336 13511 8392
rect 13372 8334 13511 8336
rect 13372 8332 13378 8334
rect 13445 8331 13511 8334
rect 16062 8332 16068 8396
rect 16132 8394 16138 8396
rect 16481 8394 16547 8397
rect 16132 8392 16547 8394
rect 16132 8336 16486 8392
rect 16542 8336 16547 8392
rect 16132 8334 16547 8336
rect 16132 8332 16138 8334
rect 16481 8331 16547 8334
rect 16798 8332 16804 8396
rect 16868 8394 16874 8396
rect 17677 8394 17743 8397
rect 16868 8392 17743 8394
rect 16868 8336 17682 8392
rect 17738 8336 17743 8392
rect 16868 8334 17743 8336
rect 16868 8332 16874 8334
rect 17677 8331 17743 8334
rect 19517 8394 19583 8397
rect 20110 8394 20116 8396
rect 19517 8392 20116 8394
rect 19517 8336 19522 8392
rect 19578 8336 20116 8392
rect 19517 8334 20116 8336
rect 19517 8331 19583 8334
rect 20110 8332 20116 8334
rect 20180 8394 20186 8396
rect 20437 8394 20503 8397
rect 20713 8396 20779 8397
rect 20180 8392 20503 8394
rect 20180 8336 20442 8392
rect 20498 8336 20503 8392
rect 20180 8334 20503 8336
rect 20180 8332 20186 8334
rect 20437 8331 20503 8334
rect 20662 8332 20668 8396
rect 20732 8394 20779 8396
rect 20732 8392 20824 8394
rect 20774 8336 20824 8392
rect 20732 8334 20824 8336
rect 20732 8332 20779 8334
rect 21582 8332 21588 8396
rect 21652 8394 21658 8396
rect 21725 8394 21791 8397
rect 21652 8392 21791 8394
rect 21652 8336 21730 8392
rect 21786 8336 21791 8392
rect 21652 8334 21791 8336
rect 21652 8332 21658 8334
rect 20713 8331 20779 8332
rect 21725 8331 21791 8334
rect 22870 8332 22876 8396
rect 22940 8394 22946 8396
rect 23013 8394 23079 8397
rect 22940 8392 23079 8394
rect 22940 8336 23018 8392
rect 23074 8336 23079 8392
rect 22940 8334 23079 8336
rect 22940 8332 22946 8334
rect 23013 8331 23079 8334
rect 23790 8332 23796 8396
rect 23860 8394 23866 8396
rect 24117 8394 24183 8397
rect 23860 8392 24183 8394
rect 23860 8336 24122 8392
rect 24178 8336 24183 8392
rect 23860 8334 24183 8336
rect 23860 8332 23866 8334
rect 24117 8331 24183 8334
rect 26785 8394 26851 8397
rect 28993 8396 29059 8397
rect 29177 8396 29243 8397
rect 27654 8394 27660 8396
rect 26785 8392 27660 8394
rect 26785 8336 26790 8392
rect 26846 8336 27660 8392
rect 26785 8334 27660 8336
rect 26785 8331 26851 8334
rect 27654 8332 27660 8334
rect 27724 8332 27730 8396
rect 28942 8394 28948 8396
rect 28902 8334 28948 8394
rect 29012 8392 29059 8396
rect 29054 8336 29059 8392
rect 28942 8332 28948 8334
rect 29012 8332 29059 8336
rect 29126 8332 29132 8396
rect 29196 8394 29243 8396
rect 29196 8392 29288 8394
rect 29238 8336 29288 8392
rect 29196 8334 29288 8336
rect 29196 8332 29243 8334
rect 28993 8331 29059 8332
rect 29177 8331 29243 8332
rect 10685 8258 10751 8261
rect 14549 8258 14615 8261
rect 10685 8256 14615 8258
rect 10685 8200 10690 8256
rect 10746 8200 14554 8256
rect 14610 8200 14615 8256
rect 10685 8198 14615 8200
rect 10685 8195 10751 8198
rect 14549 8195 14615 8198
rect 14733 8260 14799 8261
rect 15377 8260 15443 8261
rect 14733 8256 14780 8260
rect 14844 8258 14850 8260
rect 14733 8200 14738 8256
rect 14733 8196 14780 8200
rect 14844 8198 14890 8258
rect 14844 8196 14850 8198
rect 15326 8196 15332 8260
rect 15396 8258 15443 8260
rect 15396 8256 15488 8258
rect 15438 8200 15488 8256
rect 15396 8198 15488 8200
rect 15396 8196 15443 8198
rect 15878 8196 15884 8260
rect 15948 8258 15954 8260
rect 16205 8258 16271 8261
rect 15948 8256 16271 8258
rect 15948 8200 16210 8256
rect 16266 8200 16271 8256
rect 15948 8198 16271 8200
rect 15948 8196 15954 8198
rect 14733 8195 14799 8196
rect 15377 8195 15443 8196
rect 16205 8195 16271 8198
rect 17166 8196 17172 8260
rect 17236 8258 17242 8260
rect 17493 8258 17559 8261
rect 22829 8258 22895 8261
rect 17236 8256 17559 8258
rect 17236 8200 17498 8256
rect 17554 8200 17559 8256
rect 17236 8198 17559 8200
rect 17236 8196 17242 8198
rect 17493 8195 17559 8198
rect 19934 8256 22895 8258
rect 19934 8200 22834 8256
rect 22890 8200 22895 8256
rect 19934 8198 22895 8200
rect 12249 8122 12315 8125
rect 10366 8120 12315 8122
rect 10366 8064 12254 8120
rect 12310 8064 12315 8120
rect 10366 8062 12315 8064
rect 12249 8059 12315 8062
rect 12382 8060 12388 8124
rect 12452 8122 12458 8124
rect 16757 8122 16823 8125
rect 12452 8120 16823 8122
rect 12452 8064 16762 8120
rect 16818 8064 16823 8120
rect 12452 8062 16823 8064
rect 12452 8060 12458 8062
rect 16757 8059 16823 8062
rect 17769 8122 17835 8125
rect 19934 8122 19994 8198
rect 22829 8195 22895 8198
rect 23422 8196 23428 8260
rect 23492 8258 23498 8260
rect 25497 8258 25563 8261
rect 23492 8256 25563 8258
rect 23492 8200 25502 8256
rect 25558 8200 25563 8256
rect 23492 8198 25563 8200
rect 23492 8196 23498 8198
rect 25497 8195 25563 8198
rect 29821 8258 29887 8261
rect 30046 8258 30052 8260
rect 29821 8256 30052 8258
rect 29821 8200 29826 8256
rect 29882 8200 30052 8256
rect 29821 8198 30052 8200
rect 29821 8195 29887 8198
rect 30046 8196 30052 8198
rect 30116 8196 30122 8260
rect 33942 8192 34258 8193
rect 33942 8128 33948 8192
rect 34012 8128 34028 8192
rect 34092 8128 34108 8192
rect 34172 8128 34188 8192
rect 34252 8128 34258 8192
rect 33942 8127 34258 8128
rect 41942 8192 42258 8193
rect 41942 8128 41948 8192
rect 42012 8128 42028 8192
rect 42092 8128 42108 8192
rect 42172 8128 42188 8192
rect 42252 8128 42258 8192
rect 41942 8127 42258 8128
rect 17769 8120 19994 8122
rect 17769 8064 17774 8120
rect 17830 8064 19994 8120
rect 17769 8062 19994 8064
rect 20713 8122 20779 8125
rect 21030 8122 21036 8124
rect 20713 8120 21036 8122
rect 20713 8064 20718 8120
rect 20774 8064 21036 8120
rect 20713 8062 21036 8064
rect 17769 8059 17835 8062
rect 20713 8059 20779 8062
rect 21030 8060 21036 8062
rect 21100 8060 21106 8124
rect 21950 8060 21956 8124
rect 22020 8122 22026 8124
rect 23841 8122 23907 8125
rect 22020 8120 23907 8122
rect 22020 8064 23846 8120
rect 23902 8064 23907 8120
rect 22020 8062 23907 8064
rect 22020 8060 22026 8062
rect 23841 8059 23907 8062
rect 23974 8060 23980 8124
rect 24044 8122 24050 8124
rect 24669 8122 24735 8125
rect 24044 8120 24735 8122
rect 24044 8064 24674 8120
rect 24730 8064 24735 8120
rect 24044 8062 24735 8064
rect 24044 8060 24050 8062
rect 24669 8059 24735 8062
rect 27889 8122 27955 8125
rect 30741 8122 30807 8125
rect 27889 8120 30807 8122
rect 27889 8064 27894 8120
rect 27950 8064 30746 8120
rect 30802 8064 30807 8120
rect 27889 8062 30807 8064
rect 27889 8059 27955 8062
rect 30741 8059 30807 8062
rect 4889 7986 4955 7989
rect 11513 7986 11579 7989
rect 4889 7984 10058 7986
rect 4889 7928 4894 7984
rect 4950 7928 10058 7984
rect 4889 7926 10058 7928
rect 4889 7923 4955 7926
rect 6821 7850 6887 7853
rect 9998 7850 10058 7926
rect 11513 7984 15762 7986
rect 11513 7928 11518 7984
rect 11574 7928 15762 7984
rect 11513 7926 15762 7928
rect 11513 7923 11579 7926
rect 14181 7850 14247 7853
rect 6821 7848 9874 7850
rect 6821 7792 6826 7848
rect 6882 7792 9874 7848
rect 6821 7790 9874 7792
rect 9998 7848 14247 7850
rect 9998 7792 14186 7848
rect 14242 7792 14247 7848
rect 9998 7790 14247 7792
rect 6821 7787 6887 7790
rect 9814 7714 9874 7790
rect 14181 7787 14247 7790
rect 15009 7850 15075 7853
rect 15702 7850 15762 7926
rect 16246 7924 16252 7988
rect 16316 7986 16322 7988
rect 16665 7986 16731 7989
rect 16316 7984 16731 7986
rect 16316 7928 16670 7984
rect 16726 7928 16731 7984
rect 16316 7926 16731 7928
rect 16316 7924 16322 7926
rect 16665 7923 16731 7926
rect 17718 7924 17724 7988
rect 17788 7986 17794 7988
rect 17861 7986 17927 7989
rect 17788 7984 17927 7986
rect 17788 7928 17866 7984
rect 17922 7928 17927 7984
rect 17788 7926 17927 7928
rect 17788 7924 17794 7926
rect 17861 7923 17927 7926
rect 19057 7986 19123 7989
rect 23933 7986 23999 7989
rect 19057 7984 23999 7986
rect 19057 7928 19062 7984
rect 19118 7928 23938 7984
rect 23994 7928 23999 7984
rect 19057 7926 23999 7928
rect 19057 7923 19123 7926
rect 23933 7923 23999 7926
rect 27521 7986 27587 7989
rect 31661 7986 31727 7989
rect 27521 7984 31727 7986
rect 27521 7928 27526 7984
rect 27582 7928 31666 7984
rect 31722 7928 31727 7984
rect 27521 7926 31727 7928
rect 27521 7923 27587 7926
rect 31661 7923 31727 7926
rect 18965 7850 19031 7853
rect 21173 7850 21239 7853
rect 25129 7852 25195 7853
rect 15009 7848 15578 7850
rect 15009 7792 15014 7848
rect 15070 7792 15578 7848
rect 15009 7790 15578 7792
rect 15702 7848 19031 7850
rect 15702 7792 18970 7848
rect 19026 7792 19031 7848
rect 15702 7790 19031 7792
rect 15009 7787 15075 7790
rect 15285 7714 15351 7717
rect 9814 7712 15351 7714
rect 9814 7656 15290 7712
rect 15346 7656 15351 7712
rect 9814 7654 15351 7656
rect 15518 7714 15578 7790
rect 18965 7787 19031 7790
rect 19290 7848 21239 7850
rect 19290 7792 21178 7848
rect 21234 7792 21239 7848
rect 19290 7790 21239 7792
rect 16297 7714 16363 7717
rect 15518 7712 16363 7714
rect 15518 7656 16302 7712
rect 16358 7656 16363 7712
rect 15518 7654 16363 7656
rect 15285 7651 15351 7654
rect 16297 7651 16363 7654
rect 16573 7714 16639 7717
rect 19290 7714 19350 7790
rect 21173 7787 21239 7790
rect 25078 7788 25084 7852
rect 25148 7850 25195 7852
rect 27705 7850 27771 7853
rect 28206 7850 28212 7852
rect 25148 7848 25240 7850
rect 25190 7792 25240 7848
rect 25148 7790 25240 7792
rect 27705 7848 28212 7850
rect 27705 7792 27710 7848
rect 27766 7792 28212 7848
rect 27705 7790 28212 7792
rect 25148 7788 25195 7790
rect 25129 7787 25195 7788
rect 27705 7787 27771 7790
rect 28206 7788 28212 7790
rect 28276 7788 28282 7852
rect 28809 7850 28875 7853
rect 30598 7850 30604 7852
rect 28809 7848 30604 7850
rect 28809 7792 28814 7848
rect 28870 7792 30604 7848
rect 28809 7790 30604 7792
rect 28809 7787 28875 7790
rect 30598 7788 30604 7790
rect 30668 7788 30674 7852
rect 30741 7850 30807 7853
rect 32949 7850 33015 7853
rect 30741 7848 33015 7850
rect 30741 7792 30746 7848
rect 30802 7792 32954 7848
rect 33010 7792 33015 7848
rect 30741 7790 33015 7792
rect 30741 7787 30807 7790
rect 32949 7787 33015 7790
rect 16573 7712 19350 7714
rect 16573 7656 16578 7712
rect 16634 7656 19350 7712
rect 16573 7654 19350 7656
rect 16573 7651 16639 7654
rect 24342 7652 24348 7716
rect 24412 7714 24418 7716
rect 25221 7714 25287 7717
rect 26601 7714 26667 7717
rect 24412 7712 25287 7714
rect 24412 7656 25226 7712
rect 25282 7656 25287 7712
rect 24412 7654 25287 7656
rect 24412 7652 24418 7654
rect 25221 7651 25287 7654
rect 26558 7712 26667 7714
rect 26558 7656 26606 7712
rect 26662 7656 26667 7712
rect 26558 7651 26667 7656
rect 27705 7714 27771 7717
rect 31477 7714 31543 7717
rect 27705 7712 31543 7714
rect 27705 7656 27710 7712
rect 27766 7656 31482 7712
rect 31538 7656 31543 7712
rect 27705 7654 31543 7656
rect 27705 7651 27771 7654
rect 31477 7651 31543 7654
rect 31661 7714 31727 7717
rect 32857 7714 32923 7717
rect 31661 7712 32923 7714
rect 31661 7656 31666 7712
rect 31722 7656 32862 7712
rect 32918 7656 32923 7712
rect 31661 7654 32923 7656
rect 31661 7651 31727 7654
rect 32857 7651 32923 7654
rect 1302 7648 1618 7649
rect 1302 7584 1308 7648
rect 1372 7584 1388 7648
rect 1452 7584 1468 7648
rect 1532 7584 1548 7648
rect 1612 7584 1618 7648
rect 1302 7583 1618 7584
rect 9302 7648 9618 7649
rect 9302 7584 9308 7648
rect 9372 7584 9388 7648
rect 9452 7584 9468 7648
rect 9532 7584 9548 7648
rect 9612 7584 9618 7648
rect 9302 7583 9618 7584
rect 10133 7578 10199 7581
rect 10685 7578 10751 7581
rect 10133 7576 10751 7578
rect 10133 7520 10138 7576
rect 10194 7520 10690 7576
rect 10746 7520 10751 7576
rect 10133 7518 10751 7520
rect 10133 7515 10199 7518
rect 10685 7515 10751 7518
rect 11329 7578 11395 7581
rect 16987 7578 17053 7581
rect 11329 7576 17053 7578
rect 11329 7520 11334 7576
rect 11390 7520 16992 7576
rect 17048 7520 17053 7576
rect 11329 7518 17053 7520
rect 11329 7515 11395 7518
rect 16987 7515 17053 7518
rect 17861 7578 17927 7581
rect 21909 7578 21975 7581
rect 24209 7580 24275 7581
rect 24158 7578 24164 7580
rect 17861 7576 19488 7578
rect 17861 7520 17866 7576
rect 17922 7520 19488 7576
rect 17861 7518 19488 7520
rect 17861 7515 17927 7518
rect 4981 7442 5047 7445
rect 4981 7440 14106 7442
rect 4981 7384 4986 7440
rect 5042 7384 14106 7440
rect 4981 7382 14106 7384
rect 4981 7379 5047 7382
rect 14046 7374 14106 7382
rect 16614 7380 16620 7444
rect 16684 7442 16690 7444
rect 19287 7442 19353 7445
rect 16684 7440 19353 7442
rect 16684 7384 19292 7440
rect 19348 7384 19353 7440
rect 16684 7382 19353 7384
rect 19428 7442 19488 7518
rect 21909 7576 22984 7578
rect 21909 7520 21914 7576
rect 21970 7520 22984 7576
rect 21909 7518 22984 7520
rect 24118 7518 24164 7578
rect 24228 7576 24275 7580
rect 24853 7580 24919 7581
rect 26417 7580 26483 7581
rect 24853 7578 24900 7580
rect 24270 7520 24275 7576
rect 21909 7515 21975 7518
rect 19428 7382 21466 7442
rect 16684 7380 16690 7382
rect 19287 7379 19353 7382
rect 14411 7374 14477 7377
rect 14046 7372 14477 7374
rect 14046 7316 14416 7372
rect 14472 7316 14477 7372
rect 14046 7314 14477 7316
rect 21406 7374 21466 7382
rect 21955 7374 22021 7377
rect 21406 7372 22021 7374
rect 21406 7316 21960 7372
rect 22016 7316 22021 7372
rect 21406 7314 22021 7316
rect 14411 7311 14477 7314
rect 21955 7311 22021 7314
rect 8109 7306 8175 7309
rect 11881 7306 11947 7309
rect 8109 7304 11947 7306
rect 8109 7248 8114 7304
rect 8170 7248 11886 7304
rect 11942 7248 11947 7304
rect 8109 7246 11947 7248
rect 8109 7243 8175 7246
rect 11881 7243 11947 7246
rect 12249 7306 12315 7309
rect 13853 7306 13919 7309
rect 19373 7306 19439 7309
rect 12249 7304 13919 7306
rect 12249 7248 12254 7304
rect 12310 7248 13858 7304
rect 13914 7248 13919 7304
rect 12249 7246 13919 7248
rect 12249 7243 12315 7246
rect 13853 7243 13919 7246
rect 14736 7304 19439 7306
rect 14736 7248 19378 7304
rect 19434 7248 19439 7304
rect 14736 7246 19439 7248
rect 22924 7306 22984 7518
rect 24158 7516 24164 7518
rect 24228 7516 24275 7520
rect 24808 7576 24900 7578
rect 24808 7520 24858 7576
rect 24808 7518 24900 7520
rect 24209 7515 24275 7516
rect 24853 7516 24900 7518
rect 24964 7516 24970 7580
rect 26366 7578 26372 7580
rect 26326 7518 26372 7578
rect 26436 7576 26483 7580
rect 26478 7520 26483 7576
rect 26366 7516 26372 7518
rect 26436 7516 26483 7520
rect 24853 7515 24919 7516
rect 26417 7515 26483 7516
rect 23054 7380 23060 7444
rect 23124 7442 23130 7444
rect 26558 7442 26618 7651
rect 41302 7648 41618 7649
rect 41302 7584 41308 7648
rect 41372 7584 41388 7648
rect 41452 7584 41468 7648
rect 41532 7584 41548 7648
rect 41612 7584 41618 7648
rect 41302 7583 41618 7584
rect 28625 7580 28691 7581
rect 28574 7578 28580 7580
rect 28534 7518 28580 7578
rect 28644 7576 28691 7580
rect 31886 7578 31892 7580
rect 28686 7520 28691 7576
rect 28574 7516 28580 7518
rect 28644 7516 28691 7520
rect 28625 7515 28691 7516
rect 28766 7518 31892 7578
rect 23124 7382 26618 7442
rect 23124 7380 23130 7382
rect 28211 7374 28277 7377
rect 28766 7374 28826 7518
rect 31886 7516 31892 7518
rect 31956 7516 31962 7580
rect 30833 7442 30899 7445
rect 31150 7442 31156 7444
rect 30833 7440 31156 7442
rect 30833 7384 30838 7440
rect 30894 7384 31156 7440
rect 30833 7382 31156 7384
rect 30833 7379 30899 7382
rect 31150 7380 31156 7382
rect 31220 7380 31226 7444
rect 28211 7372 28826 7374
rect 28211 7316 28216 7372
rect 28272 7316 28826 7372
rect 28211 7314 28826 7316
rect 28211 7311 28277 7314
rect 24893 7306 24959 7309
rect 22924 7304 24959 7306
rect 22924 7248 24898 7304
rect 24954 7248 24959 7304
rect 22924 7246 24959 7248
rect 11094 7108 11100 7172
rect 11164 7170 11170 7172
rect 14037 7170 14103 7173
rect 11164 7168 14103 7170
rect 11164 7112 14042 7168
rect 14098 7112 14103 7168
rect 11164 7110 14103 7112
rect 11164 7108 11170 7110
rect 14037 7107 14103 7110
rect 1942 7104 2258 7105
rect 1942 7040 1948 7104
rect 2012 7040 2028 7104
rect 2092 7040 2108 7104
rect 2172 7040 2188 7104
rect 2252 7040 2258 7104
rect 1942 7039 2258 7040
rect 9942 7104 10258 7105
rect 9942 7040 9948 7104
rect 10012 7040 10028 7104
rect 10092 7040 10108 7104
rect 10172 7040 10188 7104
rect 10252 7040 10258 7104
rect 9942 7039 10258 7040
rect 10409 7034 10475 7037
rect 11605 7034 11671 7037
rect 10409 7032 11671 7034
rect 10409 6976 10414 7032
rect 10470 6976 11610 7032
rect 11666 6976 11671 7032
rect 10409 6974 11671 6976
rect 10409 6971 10475 6974
rect 11605 6971 11671 6974
rect 11881 7034 11947 7037
rect 12198 7034 12204 7036
rect 11881 7032 12204 7034
rect 11881 6976 11886 7032
rect 11942 6976 12204 7032
rect 11881 6974 12204 6976
rect 11881 6971 11947 6974
rect 12198 6972 12204 6974
rect 12268 6972 12274 7036
rect 12433 7034 12499 7037
rect 14736 7034 14796 7246
rect 19373 7243 19439 7246
rect 24893 7243 24959 7246
rect 29683 7306 29749 7309
rect 35065 7306 35131 7309
rect 29683 7304 35131 7306
rect 29683 7248 29688 7304
rect 29744 7248 35070 7304
rect 35126 7248 35131 7304
rect 29683 7246 35131 7248
rect 29683 7243 29749 7246
rect 35065 7243 35131 7246
rect 28579 7170 28645 7173
rect 29678 7170 29684 7172
rect 28579 7168 29684 7170
rect 28579 7112 28584 7168
rect 28640 7112 29684 7168
rect 28579 7110 29684 7112
rect 28579 7107 28645 7110
rect 29678 7108 29684 7110
rect 29748 7108 29754 7172
rect 14963 7104 15029 7105
rect 14958 7102 14964 7104
rect 14876 7042 14964 7102
rect 14958 7040 14964 7042
rect 15028 7040 15034 7104
rect 15142 7040 15148 7104
rect 15212 7102 15218 7104
rect 15515 7102 15581 7105
rect 17907 7102 17973 7105
rect 15212 7100 15581 7102
rect 15212 7044 15520 7100
rect 15576 7044 15581 7100
rect 15212 7042 15581 7044
rect 15212 7040 15218 7042
rect 14963 7039 15029 7040
rect 15515 7039 15581 7042
rect 17358 7100 17973 7102
rect 17358 7044 17912 7100
rect 17968 7044 17973 7100
rect 17358 7042 17973 7044
rect 17358 7034 17418 7042
rect 17907 7039 17973 7042
rect 18091 7100 18157 7105
rect 28027 7104 28093 7105
rect 30235 7104 30301 7105
rect 33942 7104 34258 7105
rect 28022 7102 28028 7104
rect 18091 7044 18096 7100
rect 18152 7044 18157 7100
rect 18091 7039 18157 7044
rect 27940 7042 28028 7102
rect 28022 7040 28028 7042
rect 28092 7040 28098 7104
rect 30230 7102 30236 7104
rect 30148 7042 30236 7102
rect 30230 7040 30236 7042
rect 30300 7040 30306 7104
rect 33942 7040 33948 7104
rect 34012 7040 34028 7104
rect 34092 7040 34108 7104
rect 34172 7040 34188 7104
rect 34252 7040 34258 7104
rect 28027 7039 28093 7040
rect 30235 7039 30301 7040
rect 33942 7039 34258 7040
rect 41942 7104 42258 7105
rect 41942 7040 41948 7104
rect 42012 7040 42028 7104
rect 42092 7040 42108 7104
rect 42172 7040 42188 7104
rect 42252 7040 42258 7104
rect 41942 7039 42258 7040
rect 12433 7032 14796 7034
rect 12433 6976 12438 7032
rect 12494 6976 14796 7032
rect 12433 6974 14796 6976
rect 15702 6974 17418 7034
rect 12433 6971 12499 6974
rect 9489 6898 9555 6901
rect 15702 6898 15762 6974
rect 9489 6896 15762 6898
rect 9489 6840 9494 6896
rect 9550 6840 15762 6896
rect 9489 6838 15762 6840
rect 9489 6835 9555 6838
rect 4889 6762 4955 6765
rect 11094 6762 11100 6764
rect 4889 6760 11100 6762
rect 4889 6704 4894 6760
rect 4950 6704 11100 6760
rect 4889 6702 11100 6704
rect 4889 6699 4955 6702
rect 11094 6700 11100 6702
rect 11164 6700 11170 6764
rect 10133 6626 10199 6629
rect 18094 6626 18154 7039
rect 10133 6624 18154 6626
rect 10133 6568 10138 6624
rect 10194 6568 18154 6624
rect 10133 6566 18154 6568
rect 10133 6563 10199 6566
rect 1302 6560 1618 6561
rect 1302 6496 1308 6560
rect 1372 6496 1388 6560
rect 1452 6496 1468 6560
rect 1532 6496 1548 6560
rect 1612 6496 1618 6560
rect 1302 6495 1618 6496
rect 9302 6560 9618 6561
rect 9302 6496 9308 6560
rect 9372 6496 9388 6560
rect 9452 6496 9468 6560
rect 9532 6496 9548 6560
rect 9612 6496 9618 6560
rect 9302 6495 9618 6496
rect 41302 6560 41618 6561
rect 41302 6496 41308 6560
rect 41372 6496 41388 6560
rect 41452 6496 41468 6560
rect 41532 6496 41548 6560
rect 41612 6496 41618 6560
rect 41302 6495 41618 6496
rect 9765 6490 9831 6493
rect 10542 6490 10548 6492
rect 9765 6488 10548 6490
rect 9765 6432 9770 6488
rect 9826 6432 10548 6488
rect 9765 6430 10548 6432
rect 9765 6427 9831 6430
rect 10542 6428 10548 6430
rect 10612 6428 10618 6492
rect 7097 6354 7163 6357
rect 15142 6354 15148 6356
rect 7097 6352 15148 6354
rect 7097 6296 7102 6352
rect 7158 6296 15148 6352
rect 7097 6294 15148 6296
rect 7097 6291 7163 6294
rect 15142 6292 15148 6294
rect 15212 6292 15218 6356
rect 31937 6354 32003 6357
rect 32622 6354 32628 6356
rect 31937 6352 32628 6354
rect 31937 6296 31942 6352
rect 31998 6296 32628 6352
rect 31937 6294 32628 6296
rect 31937 6291 32003 6294
rect 32622 6292 32628 6294
rect 32692 6292 32698 6356
rect 6269 6218 6335 6221
rect 14958 6218 14964 6220
rect 6269 6216 14964 6218
rect 6269 6160 6274 6216
rect 6330 6160 14964 6216
rect 6269 6158 14964 6160
rect 6269 6155 6335 6158
rect 14958 6156 14964 6158
rect 15028 6156 15034 6220
rect 1942 6016 2258 6017
rect 1942 5952 1948 6016
rect 2012 5952 2028 6016
rect 2092 5952 2108 6016
rect 2172 5952 2188 6016
rect 2252 5952 2258 6016
rect 1942 5951 2258 5952
rect 9942 6016 10258 6017
rect 9942 5952 9948 6016
rect 10012 5952 10028 6016
rect 10092 5952 10108 6016
rect 10172 5952 10188 6016
rect 10252 5952 10258 6016
rect 9942 5951 10258 5952
rect 33942 6016 34258 6017
rect 33942 5952 33948 6016
rect 34012 5952 34028 6016
rect 34092 5952 34108 6016
rect 34172 5952 34188 6016
rect 34252 5952 34258 6016
rect 33942 5951 34258 5952
rect 41942 6016 42258 6017
rect 41942 5952 41948 6016
rect 42012 5952 42028 6016
rect 42092 5952 42108 6016
rect 42172 5952 42188 6016
rect 42252 5952 42258 6016
rect 41942 5951 42258 5952
rect 19220 5832 19540 5840
rect 19220 5768 19228 5832
rect 19292 5768 19308 5832
rect 19372 5768 19388 5832
rect 19452 5768 19468 5832
rect 19532 5768 19540 5832
rect 19220 5752 19540 5768
rect 19220 5688 19228 5752
rect 19292 5688 19308 5752
rect 19372 5688 19388 5752
rect 19452 5688 19468 5752
rect 19532 5688 19540 5752
rect 19220 5672 19540 5688
rect 19220 5608 19228 5672
rect 19292 5608 19308 5672
rect 19372 5608 19388 5672
rect 19452 5608 19468 5672
rect 19532 5608 19540 5672
rect 19220 5592 19540 5608
rect 19220 5528 19228 5592
rect 19292 5528 19308 5592
rect 19372 5528 19388 5592
rect 19452 5528 19468 5592
rect 19532 5528 19540 5592
rect 19220 5520 19540 5528
rect 27220 5832 27540 5840
rect 27220 5768 27228 5832
rect 27292 5768 27308 5832
rect 27372 5768 27388 5832
rect 27452 5768 27468 5832
rect 27532 5768 27540 5832
rect 27220 5752 27540 5768
rect 27220 5688 27228 5752
rect 27292 5688 27308 5752
rect 27372 5688 27388 5752
rect 27452 5688 27468 5752
rect 27532 5688 27540 5752
rect 27220 5672 27540 5688
rect 27220 5608 27228 5672
rect 27292 5608 27308 5672
rect 27372 5608 27388 5672
rect 27452 5608 27468 5672
rect 27532 5608 27540 5672
rect 27220 5592 27540 5608
rect 27220 5528 27228 5592
rect 27292 5528 27308 5592
rect 27372 5528 27388 5592
rect 27452 5528 27468 5592
rect 27532 5528 27540 5592
rect 27220 5520 27540 5528
rect 1302 5472 1618 5473
rect 1302 5408 1308 5472
rect 1372 5408 1388 5472
rect 1452 5408 1468 5472
rect 1532 5408 1548 5472
rect 1612 5408 1618 5472
rect 1302 5407 1618 5408
rect 9302 5472 9618 5473
rect 9302 5408 9308 5472
rect 9372 5408 9388 5472
rect 9452 5408 9468 5472
rect 9532 5408 9548 5472
rect 9612 5408 9618 5472
rect 9302 5407 9618 5408
rect 41302 5472 41618 5473
rect 41302 5408 41308 5472
rect 41372 5408 41388 5472
rect 41452 5408 41468 5472
rect 41532 5408 41548 5472
rect 41612 5408 41618 5472
rect 41302 5407 41618 5408
rect 12985 5402 13051 5405
rect 13302 5402 13308 5404
rect 12985 5400 13308 5402
rect 12985 5344 12990 5400
rect 13046 5344 13308 5400
rect 12985 5342 13308 5344
rect 12985 5339 13051 5342
rect 13302 5340 13308 5342
rect 13372 5340 13378 5404
rect 18580 5192 18900 5200
rect 18580 5128 18588 5192
rect 18652 5128 18668 5192
rect 18732 5128 18748 5192
rect 18812 5128 18828 5192
rect 18892 5128 18900 5192
rect 18580 5112 18900 5128
rect 18580 5048 18588 5112
rect 18652 5048 18668 5112
rect 18732 5048 18748 5112
rect 18812 5048 18828 5112
rect 18892 5048 18900 5112
rect 18580 5032 18900 5048
rect 18580 4968 18588 5032
rect 18652 4968 18668 5032
rect 18732 4968 18748 5032
rect 18812 4968 18828 5032
rect 18892 4968 18900 5032
rect 18580 4952 18900 4968
rect 1942 4928 2258 4929
rect 1942 4864 1948 4928
rect 2012 4864 2028 4928
rect 2092 4864 2108 4928
rect 2172 4864 2188 4928
rect 2252 4864 2258 4928
rect 18580 4888 18588 4952
rect 18652 4888 18668 4952
rect 18732 4888 18748 4952
rect 18812 4888 18828 4952
rect 18892 4888 18900 4952
rect 18580 4880 18900 4888
rect 26580 5192 26900 5200
rect 26580 5128 26588 5192
rect 26652 5128 26668 5192
rect 26732 5128 26748 5192
rect 26812 5128 26828 5192
rect 26892 5128 26900 5192
rect 26580 5112 26900 5128
rect 26580 5048 26588 5112
rect 26652 5048 26668 5112
rect 26732 5048 26748 5112
rect 26812 5048 26828 5112
rect 26892 5048 26900 5112
rect 26580 5032 26900 5048
rect 26580 4968 26588 5032
rect 26652 4968 26668 5032
rect 26732 4968 26748 5032
rect 26812 4968 26828 5032
rect 26892 4968 26900 5032
rect 26580 4952 26900 4968
rect 26580 4888 26588 4952
rect 26652 4888 26668 4952
rect 26732 4888 26748 4952
rect 26812 4888 26828 4952
rect 26892 4888 26900 4952
rect 26580 4880 26900 4888
rect 33942 4928 34258 4929
rect 1942 4863 2258 4864
rect 33942 4864 33948 4928
rect 34012 4864 34028 4928
rect 34092 4864 34108 4928
rect 34172 4864 34188 4928
rect 34252 4864 34258 4928
rect 33942 4863 34258 4864
rect 41942 4928 42258 4929
rect 41942 4864 41948 4928
rect 42012 4864 42028 4928
rect 42092 4864 42108 4928
rect 42172 4864 42188 4928
rect 42252 4864 42258 4928
rect 41942 4863 42258 4864
rect 15694 4722 15700 4724
rect 15334 4662 15700 4722
rect 13537 4586 13603 4589
rect 14406 4586 14412 4588
rect 13537 4584 14412 4586
rect 13537 4528 13542 4584
rect 13598 4528 14412 4584
rect 13537 4526 14412 4528
rect 13537 4523 13603 4526
rect 14406 4524 14412 4526
rect 14476 4524 14482 4588
rect 14641 4586 14707 4589
rect 14774 4586 14780 4588
rect 14641 4584 14780 4586
rect 14641 4528 14646 4584
rect 14702 4528 14780 4584
rect 14641 4526 14780 4528
rect 14641 4523 14707 4526
rect 14774 4524 14780 4526
rect 14844 4524 14850 4588
rect 14917 4586 14983 4589
rect 15334 4586 15394 4662
rect 15694 4660 15700 4662
rect 15764 4660 15770 4724
rect 14917 4584 15394 4586
rect 14917 4528 14922 4584
rect 14978 4528 15394 4584
rect 14917 4526 15394 4528
rect 15469 4586 15535 4589
rect 15878 4586 15884 4588
rect 15469 4584 15884 4586
rect 15469 4528 15474 4584
rect 15530 4528 15884 4584
rect 15469 4526 15884 4528
rect 14917 4523 14983 4526
rect 15469 4523 15535 4526
rect 15878 4524 15884 4526
rect 15948 4524 15954 4588
rect 16297 4586 16363 4589
rect 16430 4586 16436 4588
rect 16297 4584 16436 4586
rect 16297 4528 16302 4584
rect 16358 4528 16436 4584
rect 16297 4526 16436 4528
rect 16297 4523 16363 4526
rect 16430 4524 16436 4526
rect 16500 4524 16506 4588
rect 16573 4586 16639 4589
rect 17166 4586 17172 4588
rect 16573 4584 17172 4586
rect 16573 4528 16578 4584
rect 16634 4528 17172 4584
rect 16573 4526 17172 4528
rect 16573 4523 16639 4526
rect 17166 4524 17172 4526
rect 17236 4524 17242 4588
rect 19333 4586 19399 4589
rect 19926 4586 19932 4588
rect 19333 4584 19932 4586
rect 19333 4528 19338 4584
rect 19394 4528 19932 4584
rect 19333 4526 19932 4528
rect 19333 4523 19399 4526
rect 19926 4524 19932 4526
rect 19996 4524 20002 4588
rect 21030 4586 21036 4588
rect 20302 4526 21036 4586
rect 13261 4450 13327 4453
rect 13670 4450 13676 4452
rect 13261 4448 13676 4450
rect 13261 4392 13266 4448
rect 13322 4392 13676 4448
rect 13261 4390 13676 4392
rect 13261 4387 13327 4390
rect 13670 4388 13676 4390
rect 13740 4388 13746 4452
rect 14365 4450 14431 4453
rect 14590 4450 14596 4452
rect 14365 4448 14596 4450
rect 14365 4392 14370 4448
rect 14426 4392 14596 4448
rect 14365 4390 14596 4392
rect 14365 4387 14431 4390
rect 14590 4388 14596 4390
rect 14660 4388 14666 4452
rect 15193 4450 15259 4453
rect 16246 4450 16252 4452
rect 15193 4448 16252 4450
rect 15193 4392 15198 4448
rect 15254 4392 16252 4448
rect 15193 4390 16252 4392
rect 15193 4387 15259 4390
rect 16246 4388 16252 4390
rect 16316 4388 16322 4452
rect 16614 4388 16620 4452
rect 16684 4450 16690 4452
rect 17677 4450 17743 4453
rect 16684 4448 17743 4450
rect 16684 4392 17682 4448
rect 17738 4392 17743 4448
rect 16684 4390 17743 4392
rect 16684 4388 16690 4390
rect 17677 4387 17743 4390
rect 18781 4450 18847 4453
rect 20302 4450 20362 4526
rect 21030 4524 21036 4526
rect 21100 4524 21106 4588
rect 22502 4524 22508 4588
rect 22572 4586 22578 4588
rect 22645 4586 22711 4589
rect 24945 4588 25011 4589
rect 22572 4584 22711 4586
rect 22572 4528 22650 4584
rect 22706 4528 22711 4584
rect 22572 4526 22711 4528
rect 22572 4524 22578 4526
rect 22645 4523 22711 4526
rect 24894 4524 24900 4588
rect 24964 4586 25011 4588
rect 26141 4586 26207 4589
rect 29126 4586 29132 4588
rect 24964 4584 25056 4586
rect 25006 4528 25056 4584
rect 24964 4526 25056 4528
rect 26141 4584 29132 4586
rect 26141 4528 26146 4584
rect 26202 4528 29132 4584
rect 26141 4526 29132 4528
rect 24964 4524 25011 4526
rect 24945 4523 25011 4524
rect 26141 4523 26207 4526
rect 29126 4524 29132 4526
rect 29196 4524 29202 4588
rect 30649 4586 30715 4589
rect 32213 4586 32279 4589
rect 30649 4584 32279 4586
rect 30649 4528 30654 4584
rect 30710 4528 32218 4584
rect 32274 4528 32279 4584
rect 30649 4526 32279 4528
rect 30649 4523 30715 4526
rect 32213 4523 32279 4526
rect 18781 4448 20362 4450
rect 18781 4392 18786 4448
rect 18842 4392 20362 4448
rect 18781 4390 20362 4392
rect 20437 4450 20503 4453
rect 22870 4450 22876 4452
rect 20437 4448 22876 4450
rect 20437 4392 20442 4448
rect 20498 4392 22876 4448
rect 20437 4390 22876 4392
rect 18781 4387 18847 4390
rect 20437 4387 20503 4390
rect 22870 4388 22876 4390
rect 22940 4388 22946 4452
rect 24342 4388 24348 4452
rect 24412 4450 24418 4452
rect 24894 4450 24900 4452
rect 24412 4390 24900 4450
rect 24412 4388 24418 4390
rect 24894 4388 24900 4390
rect 24964 4388 24970 4452
rect 25078 4388 25084 4452
rect 25148 4450 25154 4452
rect 25221 4450 25287 4453
rect 25148 4448 25287 4450
rect 25148 4392 25226 4448
rect 25282 4392 25287 4448
rect 25148 4390 25287 4392
rect 25148 4388 25154 4390
rect 25221 4387 25287 4390
rect 25773 4450 25839 4453
rect 26366 4450 26372 4452
rect 25773 4448 26372 4450
rect 25773 4392 25778 4448
rect 25834 4392 26372 4448
rect 25773 4390 26372 4392
rect 25773 4387 25839 4390
rect 26366 4388 26372 4390
rect 26436 4388 26442 4452
rect 27838 4388 27844 4452
rect 27908 4450 27914 4452
rect 28257 4450 28323 4453
rect 27908 4448 28323 4450
rect 27908 4392 28262 4448
rect 28318 4392 28323 4448
rect 27908 4390 28323 4392
rect 27908 4388 27914 4390
rect 28257 4387 28323 4390
rect 1302 4384 1618 4385
rect 1302 4320 1308 4384
rect 1372 4320 1388 4384
rect 1452 4320 1468 4384
rect 1532 4320 1548 4384
rect 1612 4320 1618 4384
rect 1302 4319 1618 4320
rect 9302 4384 9618 4385
rect 9302 4320 9308 4384
rect 9372 4320 9388 4384
rect 9452 4320 9468 4384
rect 9532 4320 9548 4384
rect 9612 4320 9618 4384
rect 9302 4319 9618 4320
rect 41302 4384 41618 4385
rect 41302 4320 41308 4384
rect 41372 4320 41388 4384
rect 41452 4320 41468 4384
rect 41532 4320 41548 4384
rect 41612 4320 41618 4384
rect 41302 4319 41618 4320
rect 17217 4314 17283 4317
rect 20846 4314 20852 4316
rect 17217 4312 20852 4314
rect 17217 4256 17222 4312
rect 17278 4256 20852 4312
rect 17217 4254 20852 4256
rect 17217 4251 17283 4254
rect 20846 4252 20852 4254
rect 20916 4252 20922 4316
rect 22369 4314 22435 4317
rect 23238 4314 23244 4316
rect 22369 4312 23244 4314
rect 22369 4256 22374 4312
rect 22430 4256 23244 4312
rect 22369 4254 23244 4256
rect 22369 4251 22435 4254
rect 23238 4252 23244 4254
rect 23308 4252 23314 4316
rect 18321 4178 18387 4181
rect 19006 4178 19012 4180
rect 18321 4176 19012 4178
rect 18321 4120 18326 4176
rect 18382 4120 19012 4176
rect 18321 4118 19012 4120
rect 18321 4115 18387 4118
rect 19006 4116 19012 4118
rect 19076 4116 19082 4180
rect 20161 4178 20227 4181
rect 20662 4178 20668 4180
rect 20161 4176 20668 4178
rect 20161 4120 20166 4176
rect 20222 4120 20668 4176
rect 20161 4118 20668 4120
rect 20161 4115 20227 4118
rect 20662 4116 20668 4118
rect 20732 4116 20738 4180
rect 20989 4178 21055 4181
rect 23974 4178 23980 4180
rect 20989 4176 23980 4178
rect 20989 4120 20994 4176
rect 21050 4120 23980 4176
rect 20989 4118 23980 4120
rect 20989 4115 21055 4118
rect 23974 4116 23980 4118
rect 24044 4116 24050 4180
rect 28441 4178 28507 4181
rect 28574 4178 28580 4180
rect 28441 4176 28580 4178
rect 28441 4120 28446 4176
rect 28502 4120 28580 4176
rect 28441 4118 28580 4120
rect 28441 4115 28507 4118
rect 28574 4116 28580 4118
rect 28644 4116 28650 4180
rect 28717 4178 28783 4181
rect 28942 4178 28948 4180
rect 28717 4176 28948 4178
rect 28717 4120 28722 4176
rect 28778 4120 28948 4176
rect 28717 4118 28948 4120
rect 28717 4115 28783 4118
rect 28942 4116 28948 4118
rect 29012 4116 29018 4180
rect 33133 4178 33199 4181
rect 33133 4176 33610 4178
rect 33133 4120 33138 4176
rect 33194 4120 33610 4176
rect 33133 4118 33610 4120
rect 33133 4115 33199 4118
rect 9673 4042 9739 4045
rect 10358 4042 10364 4044
rect 9673 4040 10364 4042
rect 9673 3984 9678 4040
rect 9734 3984 10364 4040
rect 9673 3982 10364 3984
rect 9673 3979 9739 3982
rect 10358 3980 10364 3982
rect 10428 3980 10434 4044
rect 20713 4042 20779 4045
rect 22318 4042 22324 4044
rect 20713 4040 22324 4042
rect 20713 3984 20718 4040
rect 20774 3984 22324 4040
rect 20713 3982 22324 3984
rect 20713 3979 20779 3982
rect 22318 3980 22324 3982
rect 22388 3980 22394 4044
rect 27654 3980 27660 4044
rect 27724 4042 27730 4044
rect 27797 4042 27863 4045
rect 27724 4040 27863 4042
rect 27724 3984 27802 4040
rect 27858 3984 27863 4040
rect 27724 3982 27863 3984
rect 27724 3980 27730 3982
rect 27797 3979 27863 3982
rect 30046 3980 30052 4044
rect 30116 4042 30122 4044
rect 31017 4042 31083 4045
rect 30116 4040 31083 4042
rect 30116 3984 31022 4040
rect 31078 3984 31083 4040
rect 30116 3982 31083 3984
rect 30116 3980 30122 3982
rect 31017 3979 31083 3982
rect 28022 3844 28028 3908
rect 28092 3906 28098 3908
rect 33409 3906 33475 3909
rect 28092 3904 33475 3906
rect 28092 3848 33414 3904
rect 33470 3848 33475 3904
rect 28092 3846 33475 3848
rect 28092 3844 28098 3846
rect 33409 3843 33475 3846
rect 1942 3840 2258 3841
rect 1942 3776 1948 3840
rect 2012 3776 2028 3840
rect 2092 3776 2108 3840
rect 2172 3776 2188 3840
rect 2252 3776 2258 3840
rect 1942 3775 2258 3776
rect 9942 3840 10258 3841
rect 9942 3776 9948 3840
rect 10012 3776 10028 3840
rect 10092 3776 10108 3840
rect 10172 3776 10188 3840
rect 10252 3776 10258 3840
rect 9942 3775 10258 3776
rect 32622 3708 32628 3772
rect 32692 3770 32698 3772
rect 33225 3770 33291 3773
rect 32692 3768 33291 3770
rect 32692 3712 33230 3768
rect 33286 3712 33291 3768
rect 32692 3710 33291 3712
rect 32692 3708 32698 3710
rect 33225 3707 33291 3710
rect 33550 3634 33610 4118
rect 33942 3840 34258 3841
rect 33942 3776 33948 3840
rect 34012 3776 34028 3840
rect 34092 3776 34108 3840
rect 34172 3776 34188 3840
rect 34252 3776 34258 3840
rect 33942 3775 34258 3776
rect 41942 3840 42258 3841
rect 41942 3776 41948 3840
rect 42012 3776 42028 3840
rect 42092 3776 42108 3840
rect 42172 3776 42188 3840
rect 42252 3776 42258 3840
rect 41942 3775 42258 3776
rect 34145 3634 34211 3637
rect 33550 3632 34211 3634
rect 33550 3576 34150 3632
rect 34206 3576 34211 3632
rect 33550 3574 34211 3576
rect 34145 3571 34211 3574
rect 21265 3498 21331 3501
rect 23606 3498 23612 3500
rect 21265 3496 23612 3498
rect 21265 3440 21270 3496
rect 21326 3440 23612 3496
rect 21265 3438 23612 3440
rect 21265 3435 21331 3438
rect 23606 3436 23612 3438
rect 23676 3436 23682 3500
rect 33593 3498 33659 3501
rect 35157 3498 35223 3501
rect 33593 3496 35223 3498
rect 33593 3440 33598 3496
rect 33654 3440 35162 3496
rect 35218 3440 35223 3496
rect 33593 3438 35223 3440
rect 33593 3435 33659 3438
rect 35157 3435 35223 3438
rect 36813 3362 36879 3365
rect 37273 3362 37339 3365
rect 38009 3362 38075 3365
rect 36813 3360 38075 3362
rect 36813 3304 36818 3360
rect 36874 3304 37278 3360
rect 37334 3304 38014 3360
rect 38070 3304 38075 3360
rect 36813 3302 38075 3304
rect 36813 3299 36879 3302
rect 37273 3299 37339 3302
rect 38009 3299 38075 3302
rect 1302 3296 1618 3297
rect 1302 3232 1308 3296
rect 1372 3232 1388 3296
rect 1452 3232 1468 3296
rect 1532 3232 1548 3296
rect 1612 3232 1618 3296
rect 1302 3231 1618 3232
rect 9302 3296 9618 3297
rect 9302 3232 9308 3296
rect 9372 3232 9388 3296
rect 9452 3232 9468 3296
rect 9532 3232 9548 3296
rect 9612 3232 9618 3296
rect 9302 3231 9618 3232
rect 41302 3296 41618 3297
rect 41302 3232 41308 3296
rect 41372 3232 41388 3296
rect 41452 3232 41468 3296
rect 41532 3232 41548 3296
rect 41612 3232 41618 3296
rect 41302 3231 41618 3232
rect 30230 3164 30236 3228
rect 30300 3226 30306 3228
rect 38878 3226 38884 3228
rect 30300 3166 38884 3226
rect 30300 3164 30306 3166
rect 38878 3164 38884 3166
rect 38948 3164 38954 3228
rect 32673 3090 32739 3093
rect 33225 3090 33291 3093
rect 32673 3088 33291 3090
rect 32673 3032 32678 3088
rect 32734 3032 33230 3088
rect 33286 3032 33291 3088
rect 32673 3030 33291 3032
rect 32673 3027 32739 3030
rect 33225 3027 33291 3030
rect 35065 3090 35131 3093
rect 37457 3090 37523 3093
rect 35065 3088 37523 3090
rect 35065 3032 35070 3088
rect 35126 3032 37462 3088
rect 37518 3032 37523 3088
rect 35065 3030 37523 3032
rect 35065 3027 35131 3030
rect 37457 3027 37523 3030
rect 34881 2954 34947 2957
rect 38009 2954 38075 2957
rect 39113 2954 39179 2957
rect 34881 2952 38075 2954
rect 34881 2896 34886 2952
rect 34942 2896 38014 2952
rect 38070 2896 38075 2952
rect 34881 2894 38075 2896
rect 34881 2891 34947 2894
rect 38009 2891 38075 2894
rect 38150 2952 39179 2954
rect 38150 2896 39118 2952
rect 39174 2896 39179 2952
rect 38150 2894 39179 2896
rect 36261 2818 36327 2821
rect 36905 2818 36971 2821
rect 38150 2818 38210 2894
rect 39113 2891 39179 2894
rect 36261 2816 38210 2818
rect 36261 2760 36266 2816
rect 36322 2760 36910 2816
rect 36966 2760 38210 2816
rect 36261 2758 38210 2760
rect 38285 2818 38351 2821
rect 38285 2816 38394 2818
rect 38285 2760 38290 2816
rect 38346 2760 38394 2816
rect 36261 2755 36327 2758
rect 36905 2755 36971 2758
rect 38285 2755 38394 2760
rect 1942 2752 2258 2753
rect 1942 2688 1948 2752
rect 2012 2688 2028 2752
rect 2092 2688 2108 2752
rect 2172 2688 2188 2752
rect 2252 2688 2258 2752
rect 1942 2687 2258 2688
rect 9942 2752 10258 2753
rect 9942 2688 9948 2752
rect 10012 2688 10028 2752
rect 10092 2688 10108 2752
rect 10172 2688 10188 2752
rect 10252 2688 10258 2752
rect 9942 2687 10258 2688
rect 33942 2752 34258 2753
rect 33942 2688 33948 2752
rect 34012 2688 34028 2752
rect 34092 2688 34108 2752
rect 34172 2688 34188 2752
rect 34252 2688 34258 2752
rect 33942 2687 34258 2688
rect 38334 2685 38394 2755
rect 41942 2752 42258 2753
rect 41942 2688 41948 2752
rect 42012 2688 42028 2752
rect 42092 2688 42108 2752
rect 42172 2688 42188 2752
rect 42252 2688 42258 2752
rect 41942 2687 42258 2688
rect 16849 2684 16915 2685
rect 16798 2620 16804 2684
rect 16868 2682 16915 2684
rect 16868 2680 16960 2682
rect 16910 2624 16960 2680
rect 16868 2622 16960 2624
rect 16868 2620 16915 2622
rect 28206 2620 28212 2684
rect 28276 2682 28282 2684
rect 28533 2682 28599 2685
rect 28276 2680 28599 2682
rect 28276 2624 28538 2680
rect 28594 2624 28599 2680
rect 28276 2622 28599 2624
rect 28276 2620 28282 2622
rect 16849 2619 16915 2620
rect 28533 2619 28599 2622
rect 36813 2682 36879 2685
rect 38101 2682 38167 2685
rect 36813 2680 38167 2682
rect 36813 2624 36818 2680
rect 36874 2624 38106 2680
rect 38162 2624 38167 2680
rect 36813 2622 38167 2624
rect 36813 2619 36879 2622
rect 38101 2619 38167 2622
rect 38285 2680 38394 2685
rect 38285 2624 38290 2680
rect 38346 2624 38394 2680
rect 38285 2622 38394 2624
rect 38469 2682 38535 2685
rect 40033 2682 40099 2685
rect 38469 2680 40099 2682
rect 38469 2624 38474 2680
rect 38530 2624 40038 2680
rect 40094 2624 40099 2680
rect 38469 2622 40099 2624
rect 38285 2619 38351 2622
rect 38469 2619 38535 2622
rect 40033 2619 40099 2622
rect 16982 2484 16988 2548
rect 17052 2546 17058 2548
rect 17125 2546 17191 2549
rect 17052 2544 17191 2546
rect 17052 2488 17130 2544
rect 17186 2488 17191 2544
rect 17052 2486 17191 2488
rect 17052 2484 17058 2486
rect 17125 2483 17191 2486
rect 29678 2484 29684 2548
rect 29748 2546 29754 2548
rect 36261 2546 36327 2549
rect 29748 2544 36327 2546
rect 29748 2488 36266 2544
rect 36322 2488 36327 2544
rect 29748 2486 36327 2488
rect 29748 2484 29754 2486
rect 36261 2483 36327 2486
rect 38101 2546 38167 2549
rect 38561 2546 38627 2549
rect 38745 2548 38811 2549
rect 38101 2544 38627 2546
rect 38101 2488 38106 2544
rect 38162 2488 38566 2544
rect 38622 2488 38627 2544
rect 38101 2486 38627 2488
rect 38101 2483 38167 2486
rect 38561 2483 38627 2486
rect 38694 2484 38700 2548
rect 38764 2546 38811 2548
rect 38764 2544 38856 2546
rect 38806 2488 38856 2544
rect 38764 2486 38856 2488
rect 38764 2484 38811 2486
rect 38745 2483 38811 2484
rect 37549 2410 37615 2413
rect 39389 2410 39455 2413
rect 37549 2408 39455 2410
rect 37549 2352 37554 2408
rect 37610 2352 39394 2408
rect 39450 2352 39455 2408
rect 37549 2350 39455 2352
rect 37549 2347 37615 2350
rect 39389 2347 39455 2350
rect 37549 2274 37615 2277
rect 39665 2274 39731 2277
rect 37549 2272 39731 2274
rect 37549 2216 37554 2272
rect 37610 2216 39670 2272
rect 39726 2216 39731 2272
rect 37549 2214 39731 2216
rect 37549 2211 37615 2214
rect 39665 2211 39731 2214
rect 1302 2208 1618 2209
rect 1302 2144 1308 2208
rect 1372 2144 1388 2208
rect 1452 2144 1468 2208
rect 1532 2144 1548 2208
rect 1612 2144 1618 2208
rect 1302 2143 1618 2144
rect 9302 2208 9618 2209
rect 9302 2144 9308 2208
rect 9372 2144 9388 2208
rect 9452 2144 9468 2208
rect 9532 2144 9548 2208
rect 9612 2144 9618 2208
rect 9302 2143 9618 2144
rect 17302 2208 17618 2209
rect 17302 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17468 2208
rect 17532 2144 17548 2208
rect 17612 2144 17618 2208
rect 17302 2143 17618 2144
rect 25302 2208 25618 2209
rect 25302 2144 25308 2208
rect 25372 2144 25388 2208
rect 25452 2144 25468 2208
rect 25532 2144 25548 2208
rect 25612 2144 25618 2208
rect 25302 2143 25618 2144
rect 33302 2208 33618 2209
rect 33302 2144 33308 2208
rect 33372 2144 33388 2208
rect 33452 2144 33468 2208
rect 33532 2144 33548 2208
rect 33612 2144 33618 2208
rect 33302 2143 33618 2144
rect 41302 2208 41618 2209
rect 41302 2144 41308 2208
rect 41372 2144 41388 2208
rect 41452 2144 41468 2208
rect 41532 2144 41548 2208
rect 41612 2144 41618 2208
rect 41302 2143 41618 2144
rect 36537 2138 36603 2141
rect 39021 2138 39087 2141
rect 36537 2136 39087 2138
rect 36537 2080 36542 2136
rect 36598 2080 39026 2136
rect 39082 2080 39087 2136
rect 36537 2078 39087 2080
rect 36537 2075 36603 2078
rect 39021 2075 39087 2078
rect 22553 2002 22619 2005
rect 23790 2002 23796 2004
rect 22553 2000 23796 2002
rect 22553 1944 22558 2000
rect 22614 1944 23796 2000
rect 22553 1942 23796 1944
rect 22553 1939 22619 1942
rect 23790 1940 23796 1942
rect 23860 1940 23866 2004
rect 31150 1940 31156 2004
rect 31220 2002 31226 2004
rect 33317 2002 33383 2005
rect 31220 2000 33383 2002
rect 31220 1944 33322 2000
rect 33378 1944 33383 2000
rect 31220 1942 33383 1944
rect 31220 1940 31226 1942
rect 33317 1939 33383 1942
rect 38745 2002 38811 2005
rect 39205 2002 39271 2005
rect 38745 2000 39271 2002
rect 38745 1944 38750 2000
rect 38806 1944 39210 2000
rect 39266 1944 39271 2000
rect 38745 1942 39271 1944
rect 38745 1939 38811 1942
rect 39205 1939 39271 1942
rect 23657 1866 23723 1869
rect 24158 1866 24164 1868
rect 23657 1864 24164 1866
rect 23657 1808 23662 1864
rect 23718 1808 24164 1864
rect 23657 1806 24164 1808
rect 23657 1803 23723 1806
rect 24158 1804 24164 1806
rect 24228 1804 24234 1868
rect 24894 1804 24900 1868
rect 24964 1866 24970 1868
rect 25681 1866 25747 1869
rect 24964 1864 25747 1866
rect 24964 1808 25686 1864
rect 25742 1808 25747 1864
rect 24964 1806 25747 1808
rect 24964 1804 24970 1806
rect 25681 1803 25747 1806
rect 33961 1866 34027 1869
rect 36629 1866 36695 1869
rect 33961 1864 36695 1866
rect 33961 1808 33966 1864
rect 34022 1808 36634 1864
rect 36690 1808 36695 1864
rect 33961 1806 36695 1808
rect 33961 1803 34027 1806
rect 36629 1803 36695 1806
rect 38653 1868 38719 1869
rect 38929 1868 38995 1869
rect 38653 1864 38700 1868
rect 38764 1866 38770 1868
rect 38653 1808 38658 1864
rect 38653 1804 38700 1808
rect 38764 1806 38810 1866
rect 38764 1804 38770 1806
rect 38878 1804 38884 1868
rect 38948 1866 38995 1868
rect 38948 1864 39040 1866
rect 38990 1808 39040 1864
rect 38948 1806 39040 1808
rect 38948 1804 38995 1806
rect 38653 1803 38719 1804
rect 38929 1803 38995 1804
rect 31886 1668 31892 1732
rect 31956 1730 31962 1732
rect 33777 1730 33843 1733
rect 31956 1728 33843 1730
rect 31956 1672 33782 1728
rect 33838 1672 33843 1728
rect 31956 1670 33843 1672
rect 31956 1668 31962 1670
rect 33777 1667 33843 1670
rect 1942 1664 2258 1665
rect 1942 1600 1948 1664
rect 2012 1600 2028 1664
rect 2092 1600 2108 1664
rect 2172 1600 2188 1664
rect 2252 1600 2258 1664
rect 1942 1599 2258 1600
rect 9942 1664 10258 1665
rect 9942 1600 9948 1664
rect 10012 1600 10028 1664
rect 10092 1600 10108 1664
rect 10172 1600 10188 1664
rect 10252 1600 10258 1664
rect 9942 1599 10258 1600
rect 17942 1664 18258 1665
rect 17942 1600 17948 1664
rect 18012 1600 18028 1664
rect 18092 1600 18108 1664
rect 18172 1600 18188 1664
rect 18252 1600 18258 1664
rect 17942 1599 18258 1600
rect 25942 1664 26258 1665
rect 25942 1600 25948 1664
rect 26012 1600 26028 1664
rect 26092 1600 26108 1664
rect 26172 1600 26188 1664
rect 26252 1600 26258 1664
rect 25942 1599 26258 1600
rect 33942 1664 34258 1665
rect 33942 1600 33948 1664
rect 34012 1600 34028 1664
rect 34092 1600 34108 1664
rect 34172 1600 34188 1664
rect 34252 1600 34258 1664
rect 33942 1599 34258 1600
rect 41942 1664 42258 1665
rect 41942 1600 41948 1664
rect 42012 1600 42028 1664
rect 42092 1600 42108 1664
rect 42172 1600 42188 1664
rect 42252 1600 42258 1664
rect 41942 1599 42258 1600
rect 38745 1594 38811 1597
rect 39297 1594 39363 1597
rect 40401 1594 40467 1597
rect 38745 1592 40467 1594
rect 38745 1536 38750 1592
rect 38806 1536 39302 1592
rect 39358 1536 40406 1592
rect 40462 1536 40467 1592
rect 38745 1534 40467 1536
rect 38745 1531 38811 1534
rect 39297 1531 39363 1534
rect 40401 1531 40467 1534
rect 12433 1322 12499 1325
rect 14038 1322 14044 1324
rect 12433 1320 14044 1322
rect 12433 1264 12438 1320
rect 12494 1264 14044 1320
rect 12433 1262 14044 1264
rect 12433 1259 12499 1262
rect 14038 1260 14044 1262
rect 14108 1260 14114 1324
rect 15510 1260 15516 1324
rect 15580 1322 15586 1324
rect 15745 1322 15811 1325
rect 15580 1320 15811 1322
rect 15580 1264 15750 1320
rect 15806 1264 15811 1320
rect 15580 1262 15811 1264
rect 15580 1260 15586 1262
rect 15745 1259 15811 1262
rect 16021 1322 16087 1325
rect 17718 1322 17724 1324
rect 16021 1320 17724 1322
rect 16021 1264 16026 1320
rect 16082 1264 17724 1320
rect 16021 1262 17724 1264
rect 16021 1259 16087 1262
rect 17718 1260 17724 1262
rect 17788 1260 17794 1324
rect 18505 1322 18571 1325
rect 19742 1322 19748 1324
rect 18505 1320 19748 1322
rect 18505 1264 18510 1320
rect 18566 1264 19748 1320
rect 18505 1262 19748 1264
rect 18505 1259 18571 1262
rect 19742 1260 19748 1262
rect 19812 1260 19818 1324
rect 21817 1322 21883 1325
rect 21950 1322 21956 1324
rect 21817 1320 21956 1322
rect 21817 1264 21822 1320
rect 21878 1264 21956 1320
rect 21817 1262 21956 1264
rect 21817 1259 21883 1262
rect 21950 1260 21956 1262
rect 22020 1260 22026 1324
rect 22921 1322 22987 1325
rect 23054 1322 23060 1324
rect 22921 1320 23060 1322
rect 22921 1264 22926 1320
rect 22982 1264 23060 1320
rect 22921 1262 23060 1264
rect 22921 1259 22987 1262
rect 23054 1260 23060 1262
rect 23124 1260 23130 1324
rect 23289 1322 23355 1325
rect 24526 1322 24532 1324
rect 23289 1320 24532 1322
rect 23289 1264 23294 1320
rect 23350 1264 24532 1320
rect 23289 1262 24532 1264
rect 23289 1259 23355 1262
rect 24526 1260 24532 1262
rect 24596 1260 24602 1324
rect 24710 1260 24716 1324
rect 24780 1322 24786 1324
rect 25221 1322 25287 1325
rect 24780 1320 25287 1322
rect 24780 1264 25226 1320
rect 25282 1264 25287 1320
rect 24780 1262 25287 1264
rect 24780 1260 24786 1262
rect 25221 1259 25287 1262
rect 28073 1322 28139 1325
rect 30373 1324 30439 1325
rect 28390 1322 28396 1324
rect 28073 1320 28396 1322
rect 28073 1264 28078 1320
rect 28134 1264 28396 1320
rect 28073 1262 28396 1264
rect 28073 1259 28139 1262
rect 28390 1260 28396 1262
rect 28460 1260 28466 1324
rect 30373 1320 30420 1324
rect 30484 1322 30490 1324
rect 30373 1264 30378 1320
rect 30373 1260 30420 1264
rect 30484 1262 30530 1322
rect 30484 1260 30490 1262
rect 30598 1260 30604 1324
rect 30668 1322 30674 1324
rect 30741 1322 30807 1325
rect 30668 1320 30807 1322
rect 30668 1264 30746 1320
rect 30802 1264 30807 1320
rect 30668 1262 30807 1264
rect 30668 1260 30674 1262
rect 30373 1259 30439 1260
rect 30741 1259 30807 1262
rect 30925 1324 30991 1325
rect 32949 1324 33015 1325
rect 30925 1320 30972 1324
rect 31036 1322 31042 1324
rect 30925 1264 30930 1320
rect 30925 1260 30972 1264
rect 31036 1262 31082 1322
rect 32949 1320 32996 1324
rect 33060 1322 33066 1324
rect 32949 1264 32954 1320
rect 31036 1260 31042 1262
rect 32949 1260 32996 1264
rect 33060 1262 33106 1322
rect 33060 1260 33066 1262
rect 30925 1259 30991 1260
rect 32949 1259 33015 1260
rect 13813 1186 13879 1189
rect 15326 1186 15332 1188
rect 13813 1184 15332 1186
rect 13813 1128 13818 1184
rect 13874 1128 15332 1184
rect 13813 1126 15332 1128
rect 13813 1123 13879 1126
rect 15326 1124 15332 1126
rect 15396 1124 15402 1188
rect 19057 1186 19123 1189
rect 20294 1186 20300 1188
rect 19057 1184 20300 1186
rect 19057 1128 19062 1184
rect 19118 1128 20300 1184
rect 19057 1126 20300 1128
rect 19057 1123 19123 1126
rect 20294 1124 20300 1126
rect 20364 1124 20370 1188
rect 30649 1186 30715 1189
rect 30782 1186 30788 1188
rect 30649 1184 30788 1186
rect 30649 1128 30654 1184
rect 30710 1128 30788 1184
rect 30649 1126 30788 1128
rect 30649 1123 30715 1126
rect 30782 1124 30788 1126
rect 30852 1124 30858 1188
rect 1302 1120 1618 1121
rect 1302 1056 1308 1120
rect 1372 1056 1388 1120
rect 1452 1056 1468 1120
rect 1532 1056 1548 1120
rect 1612 1056 1618 1120
rect 1302 1055 1618 1056
rect 9302 1120 9618 1121
rect 9302 1056 9308 1120
rect 9372 1056 9388 1120
rect 9452 1056 9468 1120
rect 9532 1056 9548 1120
rect 9612 1056 9618 1120
rect 9302 1055 9618 1056
rect 17302 1120 17618 1121
rect 17302 1056 17308 1120
rect 17372 1056 17388 1120
rect 17452 1056 17468 1120
rect 17532 1056 17548 1120
rect 17612 1056 17618 1120
rect 17302 1055 17618 1056
rect 25302 1120 25618 1121
rect 25302 1056 25308 1120
rect 25372 1056 25388 1120
rect 25452 1056 25468 1120
rect 25532 1056 25548 1120
rect 25612 1056 25618 1120
rect 25302 1055 25618 1056
rect 33302 1120 33618 1121
rect 33302 1056 33308 1120
rect 33372 1056 33388 1120
rect 33452 1056 33468 1120
rect 33532 1056 33548 1120
rect 33612 1056 33618 1120
rect 33302 1055 33618 1056
rect 41302 1120 41618 1121
rect 41302 1056 41308 1120
rect 41372 1056 41388 1120
rect 41452 1056 41468 1120
rect 41532 1056 41548 1120
rect 41612 1056 41618 1120
rect 41302 1055 41618 1056
rect 14089 1050 14155 1053
rect 16062 1050 16068 1052
rect 14089 1048 16068 1050
rect 14089 992 14094 1048
rect 14150 992 16068 1048
rect 14089 990 16068 992
rect 14089 987 14155 990
rect 16062 988 16068 990
rect 16132 988 16138 1052
rect 19885 1050 19951 1053
rect 21398 1050 21404 1052
rect 19885 1048 21404 1050
rect 19885 992 19890 1048
rect 19946 992 21404 1048
rect 19885 990 21404 992
rect 19885 987 19951 990
rect 21398 988 21404 990
rect 21468 988 21474 1052
rect 22093 1050 22159 1053
rect 23422 1050 23428 1052
rect 22093 1048 23428 1050
rect 22093 992 22098 1048
rect 22154 992 23428 1048
rect 22093 990 23428 992
rect 22093 987 22159 990
rect 23422 988 23428 990
rect 23492 988 23498 1052
rect 17861 914 17927 917
rect 20110 914 20116 916
rect 17861 912 20116 914
rect 17861 856 17866 912
rect 17922 856 20116 912
rect 17861 854 20116 856
rect 17861 851 17927 854
rect 20110 852 20116 854
rect 20180 852 20186 916
rect 25681 914 25747 917
rect 25957 914 26023 917
rect 25681 912 26023 914
rect 25681 856 25686 912
rect 25742 856 25962 912
rect 26018 856 26023 912
rect 25681 854 26023 856
rect 25681 851 25747 854
rect 25957 851 26023 854
rect 36261 914 36327 917
rect 41781 914 41847 917
rect 36261 912 41847 914
rect 36261 856 36266 912
rect 36322 856 41786 912
rect 41842 856 41847 912
rect 36261 854 41847 856
rect 36261 851 36327 854
rect 41781 851 41847 854
rect 19609 778 19675 781
rect 21582 778 21588 780
rect 19609 776 21588 778
rect 19609 720 19614 776
rect 19670 720 21588 776
rect 19609 718 21588 720
rect 19609 715 19675 718
rect 21582 716 21588 718
rect 21652 716 21658 780
rect 38653 778 38719 781
rect 40493 778 40559 781
rect 42333 778 42399 781
rect 38653 776 42399 778
rect 38653 720 38658 776
rect 38714 720 40498 776
rect 40554 720 42338 776
rect 42394 720 42399 776
rect 38653 718 42399 720
rect 38653 715 38719 718
rect 40493 715 40559 718
rect 42333 715 42399 718
rect 40401 642 40467 645
rect 41321 642 41387 645
rect 40401 640 41387 642
rect 40401 584 40406 640
rect 40462 584 41326 640
rect 41382 584 41387 640
rect 40401 582 41387 584
rect 40401 579 40467 582
rect 41321 579 41387 582
rect 1942 576 2258 577
rect 1942 512 1948 576
rect 2012 512 2028 576
rect 2092 512 2108 576
rect 2172 512 2188 576
rect 2252 512 2258 576
rect 1942 511 2258 512
rect 9942 576 10258 577
rect 9942 512 9948 576
rect 10012 512 10028 576
rect 10092 512 10108 576
rect 10172 512 10188 576
rect 10252 512 10258 576
rect 9942 511 10258 512
rect 17942 576 18258 577
rect 17942 512 17948 576
rect 18012 512 18028 576
rect 18092 512 18108 576
rect 18172 512 18188 576
rect 18252 512 18258 576
rect 17942 511 18258 512
rect 25942 576 26258 577
rect 25942 512 25948 576
rect 26012 512 26028 576
rect 26092 512 26108 576
rect 26172 512 26188 576
rect 26252 512 26258 576
rect 25942 511 26258 512
rect 33942 576 34258 577
rect 33942 512 33948 576
rect 34012 512 34028 576
rect 34092 512 34108 576
rect 34172 512 34188 576
rect 34252 512 34258 576
rect 33942 511 34258 512
rect 41942 576 42258 577
rect 41942 512 41948 576
rect 42012 512 42028 576
rect 42092 512 42108 576
rect 42172 512 42188 576
rect 42252 512 42258 576
rect 41942 511 42258 512
<< via3 >>
rect 1948 11452 2012 11456
rect 1948 11396 1952 11452
rect 1952 11396 2008 11452
rect 2008 11396 2012 11452
rect 1948 11392 2012 11396
rect 2028 11452 2092 11456
rect 2028 11396 2032 11452
rect 2032 11396 2088 11452
rect 2088 11396 2092 11452
rect 2028 11392 2092 11396
rect 2108 11452 2172 11456
rect 2108 11396 2112 11452
rect 2112 11396 2168 11452
rect 2168 11396 2172 11452
rect 2108 11392 2172 11396
rect 2188 11452 2252 11456
rect 2188 11396 2192 11452
rect 2192 11396 2248 11452
rect 2248 11396 2252 11452
rect 2188 11392 2252 11396
rect 9948 11452 10012 11456
rect 9948 11396 9952 11452
rect 9952 11396 10008 11452
rect 10008 11396 10012 11452
rect 9948 11392 10012 11396
rect 10028 11452 10092 11456
rect 10028 11396 10032 11452
rect 10032 11396 10088 11452
rect 10088 11396 10092 11452
rect 10028 11392 10092 11396
rect 10108 11452 10172 11456
rect 10108 11396 10112 11452
rect 10112 11396 10168 11452
rect 10168 11396 10172 11452
rect 10108 11392 10172 11396
rect 10188 11452 10252 11456
rect 10188 11396 10192 11452
rect 10192 11396 10248 11452
rect 10248 11396 10252 11452
rect 10188 11392 10252 11396
rect 17948 11452 18012 11456
rect 17948 11396 17952 11452
rect 17952 11396 18008 11452
rect 18008 11396 18012 11452
rect 17948 11392 18012 11396
rect 18028 11452 18092 11456
rect 18028 11396 18032 11452
rect 18032 11396 18088 11452
rect 18088 11396 18092 11452
rect 18028 11392 18092 11396
rect 18108 11452 18172 11456
rect 18108 11396 18112 11452
rect 18112 11396 18168 11452
rect 18168 11396 18172 11452
rect 18108 11392 18172 11396
rect 18188 11452 18252 11456
rect 18188 11396 18192 11452
rect 18192 11396 18248 11452
rect 18248 11396 18252 11452
rect 18188 11392 18252 11396
rect 25948 11452 26012 11456
rect 25948 11396 25952 11452
rect 25952 11396 26008 11452
rect 26008 11396 26012 11452
rect 25948 11392 26012 11396
rect 26028 11452 26092 11456
rect 26028 11396 26032 11452
rect 26032 11396 26088 11452
rect 26088 11396 26092 11452
rect 26028 11392 26092 11396
rect 26108 11452 26172 11456
rect 26108 11396 26112 11452
rect 26112 11396 26168 11452
rect 26168 11396 26172 11452
rect 26108 11392 26172 11396
rect 26188 11452 26252 11456
rect 26188 11396 26192 11452
rect 26192 11396 26248 11452
rect 26248 11396 26252 11452
rect 26188 11392 26252 11396
rect 33948 11452 34012 11456
rect 33948 11396 33952 11452
rect 33952 11396 34008 11452
rect 34008 11396 34012 11452
rect 33948 11392 34012 11396
rect 34028 11452 34092 11456
rect 34028 11396 34032 11452
rect 34032 11396 34088 11452
rect 34088 11396 34092 11452
rect 34028 11392 34092 11396
rect 34108 11452 34172 11456
rect 34108 11396 34112 11452
rect 34112 11396 34168 11452
rect 34168 11396 34172 11452
rect 34108 11392 34172 11396
rect 34188 11452 34252 11456
rect 34188 11396 34192 11452
rect 34192 11396 34248 11452
rect 34248 11396 34252 11452
rect 34188 11392 34252 11396
rect 41948 11452 42012 11456
rect 41948 11396 41952 11452
rect 41952 11396 42008 11452
rect 42008 11396 42012 11452
rect 41948 11392 42012 11396
rect 42028 11452 42092 11456
rect 42028 11396 42032 11452
rect 42032 11396 42088 11452
rect 42088 11396 42092 11452
rect 42028 11392 42092 11396
rect 42108 11452 42172 11456
rect 42108 11396 42112 11452
rect 42112 11396 42168 11452
rect 42168 11396 42172 11452
rect 42108 11392 42172 11396
rect 42188 11452 42252 11456
rect 42188 11396 42192 11452
rect 42192 11396 42248 11452
rect 42248 11396 42252 11452
rect 42188 11392 42252 11396
rect 1308 10908 1372 10912
rect 1308 10852 1312 10908
rect 1312 10852 1368 10908
rect 1368 10852 1372 10908
rect 1308 10848 1372 10852
rect 1388 10908 1452 10912
rect 1388 10852 1392 10908
rect 1392 10852 1448 10908
rect 1448 10852 1452 10908
rect 1388 10848 1452 10852
rect 1468 10908 1532 10912
rect 1468 10852 1472 10908
rect 1472 10852 1528 10908
rect 1528 10852 1532 10908
rect 1468 10848 1532 10852
rect 1548 10908 1612 10912
rect 1548 10852 1552 10908
rect 1552 10852 1608 10908
rect 1608 10852 1612 10908
rect 1548 10848 1612 10852
rect 9308 10908 9372 10912
rect 9308 10852 9312 10908
rect 9312 10852 9368 10908
rect 9368 10852 9372 10908
rect 9308 10848 9372 10852
rect 9388 10908 9452 10912
rect 9388 10852 9392 10908
rect 9392 10852 9448 10908
rect 9448 10852 9452 10908
rect 9388 10848 9452 10852
rect 9468 10908 9532 10912
rect 9468 10852 9472 10908
rect 9472 10852 9528 10908
rect 9528 10852 9532 10908
rect 9468 10848 9532 10852
rect 9548 10908 9612 10912
rect 9548 10852 9552 10908
rect 9552 10852 9608 10908
rect 9608 10852 9612 10908
rect 9548 10848 9612 10852
rect 17308 10908 17372 10912
rect 17308 10852 17312 10908
rect 17312 10852 17368 10908
rect 17368 10852 17372 10908
rect 17308 10848 17372 10852
rect 17388 10908 17452 10912
rect 17388 10852 17392 10908
rect 17392 10852 17448 10908
rect 17448 10852 17452 10908
rect 17388 10848 17452 10852
rect 17468 10908 17532 10912
rect 17468 10852 17472 10908
rect 17472 10852 17528 10908
rect 17528 10852 17532 10908
rect 17468 10848 17532 10852
rect 17548 10908 17612 10912
rect 17548 10852 17552 10908
rect 17552 10852 17608 10908
rect 17608 10852 17612 10908
rect 17548 10848 17612 10852
rect 25308 10908 25372 10912
rect 25308 10852 25312 10908
rect 25312 10852 25368 10908
rect 25368 10852 25372 10908
rect 25308 10848 25372 10852
rect 25388 10908 25452 10912
rect 25388 10852 25392 10908
rect 25392 10852 25448 10908
rect 25448 10852 25452 10908
rect 25388 10848 25452 10852
rect 25468 10908 25532 10912
rect 25468 10852 25472 10908
rect 25472 10852 25528 10908
rect 25528 10852 25532 10908
rect 25468 10848 25532 10852
rect 25548 10908 25612 10912
rect 25548 10852 25552 10908
rect 25552 10852 25608 10908
rect 25608 10852 25612 10908
rect 25548 10848 25612 10852
rect 33308 10908 33372 10912
rect 33308 10852 33312 10908
rect 33312 10852 33368 10908
rect 33368 10852 33372 10908
rect 33308 10848 33372 10852
rect 33388 10908 33452 10912
rect 33388 10852 33392 10908
rect 33392 10852 33448 10908
rect 33448 10852 33452 10908
rect 33388 10848 33452 10852
rect 33468 10908 33532 10912
rect 33468 10852 33472 10908
rect 33472 10852 33528 10908
rect 33528 10852 33532 10908
rect 33468 10848 33532 10852
rect 33548 10908 33612 10912
rect 33548 10852 33552 10908
rect 33552 10852 33608 10908
rect 33608 10852 33612 10908
rect 33548 10848 33612 10852
rect 41308 10908 41372 10912
rect 41308 10852 41312 10908
rect 41312 10852 41368 10908
rect 41368 10852 41372 10908
rect 41308 10848 41372 10852
rect 41388 10908 41452 10912
rect 41388 10852 41392 10908
rect 41392 10852 41448 10908
rect 41448 10852 41452 10908
rect 41388 10848 41452 10852
rect 41468 10908 41532 10912
rect 41468 10852 41472 10908
rect 41472 10852 41528 10908
rect 41528 10852 41532 10908
rect 41468 10848 41532 10852
rect 41548 10908 41612 10912
rect 41548 10852 41552 10908
rect 41552 10852 41608 10908
rect 41608 10852 41612 10908
rect 41548 10848 41612 10852
rect 1948 10364 2012 10368
rect 1948 10308 1952 10364
rect 1952 10308 2008 10364
rect 2008 10308 2012 10364
rect 1948 10304 2012 10308
rect 2028 10364 2092 10368
rect 2028 10308 2032 10364
rect 2032 10308 2088 10364
rect 2088 10308 2092 10364
rect 2028 10304 2092 10308
rect 2108 10364 2172 10368
rect 2108 10308 2112 10364
rect 2112 10308 2168 10364
rect 2168 10308 2172 10364
rect 2108 10304 2172 10308
rect 2188 10364 2252 10368
rect 2188 10308 2192 10364
rect 2192 10308 2248 10364
rect 2248 10308 2252 10364
rect 2188 10304 2252 10308
rect 9948 10364 10012 10368
rect 9948 10308 9952 10364
rect 9952 10308 10008 10364
rect 10008 10308 10012 10364
rect 9948 10304 10012 10308
rect 10028 10364 10092 10368
rect 10028 10308 10032 10364
rect 10032 10308 10088 10364
rect 10088 10308 10092 10364
rect 10028 10304 10092 10308
rect 10108 10364 10172 10368
rect 10108 10308 10112 10364
rect 10112 10308 10168 10364
rect 10168 10308 10172 10364
rect 10108 10304 10172 10308
rect 10188 10364 10252 10368
rect 10188 10308 10192 10364
rect 10192 10308 10248 10364
rect 10248 10308 10252 10364
rect 10188 10304 10252 10308
rect 17948 10364 18012 10368
rect 17948 10308 17952 10364
rect 17952 10308 18008 10364
rect 18008 10308 18012 10364
rect 17948 10304 18012 10308
rect 18028 10364 18092 10368
rect 18028 10308 18032 10364
rect 18032 10308 18088 10364
rect 18088 10308 18092 10364
rect 18028 10304 18092 10308
rect 18108 10364 18172 10368
rect 18108 10308 18112 10364
rect 18112 10308 18168 10364
rect 18168 10308 18172 10364
rect 18108 10304 18172 10308
rect 18188 10364 18252 10368
rect 18188 10308 18192 10364
rect 18192 10308 18248 10364
rect 18248 10308 18252 10364
rect 18188 10304 18252 10308
rect 25948 10364 26012 10368
rect 25948 10308 25952 10364
rect 25952 10308 26008 10364
rect 26008 10308 26012 10364
rect 25948 10304 26012 10308
rect 26028 10364 26092 10368
rect 26028 10308 26032 10364
rect 26032 10308 26088 10364
rect 26088 10308 26092 10364
rect 26028 10304 26092 10308
rect 26108 10364 26172 10368
rect 26108 10308 26112 10364
rect 26112 10308 26168 10364
rect 26168 10308 26172 10364
rect 26108 10304 26172 10308
rect 26188 10364 26252 10368
rect 26188 10308 26192 10364
rect 26192 10308 26248 10364
rect 26248 10308 26252 10364
rect 26188 10304 26252 10308
rect 33948 10364 34012 10368
rect 33948 10308 33952 10364
rect 33952 10308 34008 10364
rect 34008 10308 34012 10364
rect 33948 10304 34012 10308
rect 34028 10364 34092 10368
rect 34028 10308 34032 10364
rect 34032 10308 34088 10364
rect 34088 10308 34092 10364
rect 34028 10304 34092 10308
rect 34108 10364 34172 10368
rect 34108 10308 34112 10364
rect 34112 10308 34168 10364
rect 34168 10308 34172 10364
rect 34108 10304 34172 10308
rect 34188 10364 34252 10368
rect 34188 10308 34192 10364
rect 34192 10308 34248 10364
rect 34248 10308 34252 10364
rect 34188 10304 34252 10308
rect 41948 10364 42012 10368
rect 41948 10308 41952 10364
rect 41952 10308 42008 10364
rect 42008 10308 42012 10364
rect 41948 10304 42012 10308
rect 42028 10364 42092 10368
rect 42028 10308 42032 10364
rect 42032 10308 42088 10364
rect 42088 10308 42092 10364
rect 42028 10304 42092 10308
rect 42108 10364 42172 10368
rect 42108 10308 42112 10364
rect 42112 10308 42168 10364
rect 42168 10308 42172 10364
rect 42108 10304 42172 10308
rect 42188 10364 42252 10368
rect 42188 10308 42192 10364
rect 42192 10308 42248 10364
rect 42248 10308 42252 10364
rect 42188 10304 42252 10308
rect 1308 9820 1372 9824
rect 1308 9764 1312 9820
rect 1312 9764 1368 9820
rect 1368 9764 1372 9820
rect 1308 9760 1372 9764
rect 1388 9820 1452 9824
rect 1388 9764 1392 9820
rect 1392 9764 1448 9820
rect 1448 9764 1452 9820
rect 1388 9760 1452 9764
rect 1468 9820 1532 9824
rect 1468 9764 1472 9820
rect 1472 9764 1528 9820
rect 1528 9764 1532 9820
rect 1468 9760 1532 9764
rect 1548 9820 1612 9824
rect 1548 9764 1552 9820
rect 1552 9764 1608 9820
rect 1608 9764 1612 9820
rect 1548 9760 1612 9764
rect 9308 9820 9372 9824
rect 9308 9764 9312 9820
rect 9312 9764 9368 9820
rect 9368 9764 9372 9820
rect 9308 9760 9372 9764
rect 9388 9820 9452 9824
rect 9388 9764 9392 9820
rect 9392 9764 9448 9820
rect 9448 9764 9452 9820
rect 9388 9760 9452 9764
rect 9468 9820 9532 9824
rect 9468 9764 9472 9820
rect 9472 9764 9528 9820
rect 9528 9764 9532 9820
rect 9468 9760 9532 9764
rect 9548 9820 9612 9824
rect 9548 9764 9552 9820
rect 9552 9764 9608 9820
rect 9608 9764 9612 9820
rect 9548 9760 9612 9764
rect 17308 9820 17372 9824
rect 17308 9764 17312 9820
rect 17312 9764 17368 9820
rect 17368 9764 17372 9820
rect 17308 9760 17372 9764
rect 17388 9820 17452 9824
rect 17388 9764 17392 9820
rect 17392 9764 17448 9820
rect 17448 9764 17452 9820
rect 17388 9760 17452 9764
rect 17468 9820 17532 9824
rect 17468 9764 17472 9820
rect 17472 9764 17528 9820
rect 17528 9764 17532 9820
rect 17468 9760 17532 9764
rect 17548 9820 17612 9824
rect 17548 9764 17552 9820
rect 17552 9764 17608 9820
rect 17608 9764 17612 9820
rect 17548 9760 17612 9764
rect 25308 9820 25372 9824
rect 25308 9764 25312 9820
rect 25312 9764 25368 9820
rect 25368 9764 25372 9820
rect 25308 9760 25372 9764
rect 25388 9820 25452 9824
rect 25388 9764 25392 9820
rect 25392 9764 25448 9820
rect 25448 9764 25452 9820
rect 25388 9760 25452 9764
rect 25468 9820 25532 9824
rect 25468 9764 25472 9820
rect 25472 9764 25528 9820
rect 25528 9764 25532 9820
rect 25468 9760 25532 9764
rect 25548 9820 25612 9824
rect 25548 9764 25552 9820
rect 25552 9764 25608 9820
rect 25608 9764 25612 9820
rect 25548 9760 25612 9764
rect 33308 9820 33372 9824
rect 33308 9764 33312 9820
rect 33312 9764 33368 9820
rect 33368 9764 33372 9820
rect 33308 9760 33372 9764
rect 33388 9820 33452 9824
rect 33388 9764 33392 9820
rect 33392 9764 33448 9820
rect 33448 9764 33452 9820
rect 33388 9760 33452 9764
rect 33468 9820 33532 9824
rect 33468 9764 33472 9820
rect 33472 9764 33528 9820
rect 33528 9764 33532 9820
rect 33468 9760 33532 9764
rect 33548 9820 33612 9824
rect 33548 9764 33552 9820
rect 33552 9764 33608 9820
rect 33608 9764 33612 9820
rect 33548 9760 33612 9764
rect 41308 9820 41372 9824
rect 41308 9764 41312 9820
rect 41312 9764 41368 9820
rect 41368 9764 41372 9820
rect 41308 9760 41372 9764
rect 41388 9820 41452 9824
rect 41388 9764 41392 9820
rect 41392 9764 41448 9820
rect 41448 9764 41452 9820
rect 41388 9760 41452 9764
rect 41468 9820 41532 9824
rect 41468 9764 41472 9820
rect 41472 9764 41528 9820
rect 41528 9764 41532 9820
rect 41468 9760 41532 9764
rect 41548 9820 41612 9824
rect 41548 9764 41552 9820
rect 41552 9764 41608 9820
rect 41608 9764 41612 9820
rect 41548 9760 41612 9764
rect 24532 9752 24596 9756
rect 24532 9696 24546 9752
rect 24546 9696 24596 9752
rect 24532 9692 24596 9696
rect 24716 9752 24780 9756
rect 24716 9696 24730 9752
rect 24730 9696 24780 9752
rect 24716 9692 24780 9696
rect 32996 9692 33060 9756
rect 14044 9480 14108 9484
rect 14044 9424 14094 9480
rect 14094 9424 14108 9480
rect 14044 9420 14108 9424
rect 14596 9420 14660 9484
rect 1948 9276 2012 9280
rect 1948 9220 1952 9276
rect 1952 9220 2008 9276
rect 2008 9220 2012 9276
rect 1948 9216 2012 9220
rect 2028 9276 2092 9280
rect 2028 9220 2032 9276
rect 2032 9220 2088 9276
rect 2088 9220 2092 9276
rect 2028 9216 2092 9220
rect 2108 9276 2172 9280
rect 2108 9220 2112 9276
rect 2112 9220 2168 9276
rect 2168 9220 2172 9276
rect 2108 9216 2172 9220
rect 2188 9276 2252 9280
rect 2188 9220 2192 9276
rect 2192 9220 2248 9276
rect 2248 9220 2252 9276
rect 2188 9216 2252 9220
rect 9948 9276 10012 9280
rect 9948 9220 9952 9276
rect 9952 9220 10008 9276
rect 10008 9220 10012 9276
rect 9948 9216 10012 9220
rect 10028 9276 10092 9280
rect 10028 9220 10032 9276
rect 10032 9220 10088 9276
rect 10088 9220 10092 9276
rect 10028 9216 10092 9220
rect 10108 9276 10172 9280
rect 10108 9220 10112 9276
rect 10112 9220 10168 9276
rect 10168 9220 10172 9276
rect 10108 9216 10172 9220
rect 10188 9276 10252 9280
rect 10188 9220 10192 9276
rect 10192 9220 10248 9276
rect 10248 9220 10252 9276
rect 10188 9216 10252 9220
rect 22324 9284 22388 9348
rect 33948 9276 34012 9280
rect 33948 9220 33952 9276
rect 33952 9220 34008 9276
rect 34008 9220 34012 9276
rect 33948 9216 34012 9220
rect 34028 9276 34092 9280
rect 34028 9220 34032 9276
rect 34032 9220 34088 9276
rect 34088 9220 34092 9276
rect 34028 9216 34092 9220
rect 34108 9276 34172 9280
rect 34108 9220 34112 9276
rect 34112 9220 34168 9276
rect 34168 9220 34172 9276
rect 34108 9216 34172 9220
rect 34188 9276 34252 9280
rect 34188 9220 34192 9276
rect 34192 9220 34248 9276
rect 34248 9220 34252 9276
rect 34188 9216 34252 9220
rect 41948 9276 42012 9280
rect 41948 9220 41952 9276
rect 41952 9220 42008 9276
rect 42008 9220 42012 9276
rect 41948 9216 42012 9220
rect 42028 9276 42092 9280
rect 42028 9220 42032 9276
rect 42032 9220 42088 9276
rect 42088 9220 42092 9276
rect 42028 9216 42092 9220
rect 42108 9276 42172 9280
rect 42108 9220 42112 9276
rect 42112 9220 42168 9276
rect 42168 9220 42172 9276
rect 42108 9216 42172 9220
rect 42188 9276 42252 9280
rect 42188 9220 42192 9276
rect 42192 9220 42248 9276
rect 42248 9220 42252 9276
rect 42188 9216 42252 9220
rect 23244 9148 23308 9212
rect 14412 9012 14476 9076
rect 22508 9012 22572 9076
rect 13676 8876 13740 8940
rect 16068 8876 16132 8940
rect 16436 8876 16500 8940
rect 19012 8876 19076 8940
rect 19748 8876 19812 8940
rect 19932 8936 19996 8940
rect 19932 8880 19982 8936
rect 19982 8880 19996 8936
rect 19932 8876 19996 8880
rect 20300 8876 20364 8940
rect 23612 8876 23676 8940
rect 30788 8876 30852 8940
rect 10548 8740 10612 8804
rect 15700 8740 15764 8804
rect 1308 8732 1372 8736
rect 1308 8676 1312 8732
rect 1312 8676 1368 8732
rect 1368 8676 1372 8732
rect 1308 8672 1372 8676
rect 1388 8732 1452 8736
rect 1388 8676 1392 8732
rect 1392 8676 1448 8732
rect 1448 8676 1452 8732
rect 1388 8672 1452 8676
rect 1468 8732 1532 8736
rect 1468 8676 1472 8732
rect 1472 8676 1528 8732
rect 1528 8676 1532 8732
rect 1468 8672 1532 8676
rect 1548 8732 1612 8736
rect 1548 8676 1552 8732
rect 1552 8676 1608 8732
rect 1608 8676 1612 8732
rect 1548 8672 1612 8676
rect 9308 8732 9372 8736
rect 9308 8676 9312 8732
rect 9312 8676 9368 8732
rect 9368 8676 9372 8732
rect 9308 8672 9372 8676
rect 9388 8732 9452 8736
rect 9388 8676 9392 8732
rect 9392 8676 9448 8732
rect 9448 8676 9452 8732
rect 9388 8672 9452 8676
rect 9468 8732 9532 8736
rect 9468 8676 9472 8732
rect 9472 8676 9528 8732
rect 9528 8676 9532 8732
rect 9468 8672 9532 8676
rect 9548 8732 9612 8736
rect 9548 8676 9552 8732
rect 9552 8676 9608 8732
rect 9608 8676 9612 8732
rect 9548 8672 9612 8676
rect 9812 8604 9876 8668
rect 10364 8604 10428 8668
rect 15516 8604 15580 8668
rect 30420 8740 30484 8804
rect 41308 8732 41372 8736
rect 41308 8676 41312 8732
rect 41312 8676 41368 8732
rect 41368 8676 41372 8732
rect 41308 8672 41372 8676
rect 41388 8732 41452 8736
rect 41388 8676 41392 8732
rect 41392 8676 41448 8732
rect 41448 8676 41452 8732
rect 41388 8672 41452 8676
rect 41468 8732 41532 8736
rect 41468 8676 41472 8732
rect 41472 8676 41528 8732
rect 41528 8676 41532 8732
rect 41468 8672 41532 8676
rect 41548 8732 41612 8736
rect 41548 8676 41552 8732
rect 41552 8676 41608 8732
rect 41608 8676 41612 8732
rect 41548 8672 41612 8676
rect 28396 8604 28460 8668
rect 16988 8468 17052 8532
rect 20852 8468 20916 8532
rect 21404 8468 21468 8532
rect 27844 8468 27908 8532
rect 30972 8468 31036 8532
rect 1948 8188 2012 8192
rect 1948 8132 1952 8188
rect 1952 8132 2008 8188
rect 2008 8132 2012 8188
rect 1948 8128 2012 8132
rect 2028 8188 2092 8192
rect 2028 8132 2032 8188
rect 2032 8132 2088 8188
rect 2088 8132 2092 8188
rect 2028 8128 2092 8132
rect 2108 8188 2172 8192
rect 2108 8132 2112 8188
rect 2112 8132 2168 8188
rect 2168 8132 2172 8188
rect 2108 8128 2172 8132
rect 2188 8188 2252 8192
rect 2188 8132 2192 8188
rect 2192 8132 2248 8188
rect 2248 8132 2252 8188
rect 2188 8128 2252 8132
rect 9948 8188 10012 8192
rect 9948 8132 9952 8188
rect 9952 8132 10008 8188
rect 10008 8132 10012 8188
rect 9948 8128 10012 8132
rect 10028 8188 10092 8192
rect 10028 8132 10032 8188
rect 10032 8132 10088 8188
rect 10088 8132 10092 8188
rect 10028 8128 10092 8132
rect 10108 8188 10172 8192
rect 10108 8132 10112 8188
rect 10112 8132 10168 8188
rect 10168 8132 10172 8188
rect 10108 8128 10172 8132
rect 10188 8188 10252 8192
rect 10188 8132 10192 8188
rect 10192 8132 10248 8188
rect 10248 8132 10252 8188
rect 10188 8128 10252 8132
rect 9812 8060 9876 8124
rect 13308 8332 13372 8396
rect 16068 8332 16132 8396
rect 16804 8332 16868 8396
rect 20116 8332 20180 8396
rect 20668 8392 20732 8396
rect 20668 8336 20718 8392
rect 20718 8336 20732 8392
rect 20668 8332 20732 8336
rect 21588 8332 21652 8396
rect 22876 8332 22940 8396
rect 23796 8332 23860 8396
rect 27660 8332 27724 8396
rect 28948 8392 29012 8396
rect 28948 8336 28998 8392
rect 28998 8336 29012 8392
rect 28948 8332 29012 8336
rect 29132 8392 29196 8396
rect 29132 8336 29182 8392
rect 29182 8336 29196 8392
rect 29132 8332 29196 8336
rect 14780 8256 14844 8260
rect 14780 8200 14794 8256
rect 14794 8200 14844 8256
rect 14780 8196 14844 8200
rect 15332 8256 15396 8260
rect 15332 8200 15382 8256
rect 15382 8200 15396 8256
rect 15332 8196 15396 8200
rect 15884 8196 15948 8260
rect 17172 8196 17236 8260
rect 12388 8060 12452 8124
rect 23428 8196 23492 8260
rect 30052 8196 30116 8260
rect 33948 8188 34012 8192
rect 33948 8132 33952 8188
rect 33952 8132 34008 8188
rect 34008 8132 34012 8188
rect 33948 8128 34012 8132
rect 34028 8188 34092 8192
rect 34028 8132 34032 8188
rect 34032 8132 34088 8188
rect 34088 8132 34092 8188
rect 34028 8128 34092 8132
rect 34108 8188 34172 8192
rect 34108 8132 34112 8188
rect 34112 8132 34168 8188
rect 34168 8132 34172 8188
rect 34108 8128 34172 8132
rect 34188 8188 34252 8192
rect 34188 8132 34192 8188
rect 34192 8132 34248 8188
rect 34248 8132 34252 8188
rect 34188 8128 34252 8132
rect 41948 8188 42012 8192
rect 41948 8132 41952 8188
rect 41952 8132 42008 8188
rect 42008 8132 42012 8188
rect 41948 8128 42012 8132
rect 42028 8188 42092 8192
rect 42028 8132 42032 8188
rect 42032 8132 42088 8188
rect 42088 8132 42092 8188
rect 42028 8128 42092 8132
rect 42108 8188 42172 8192
rect 42108 8132 42112 8188
rect 42112 8132 42168 8188
rect 42168 8132 42172 8188
rect 42108 8128 42172 8132
rect 42188 8188 42252 8192
rect 42188 8132 42192 8188
rect 42192 8132 42248 8188
rect 42248 8132 42252 8188
rect 42188 8128 42252 8132
rect 21036 8060 21100 8124
rect 21956 8060 22020 8124
rect 23980 8060 24044 8124
rect 16252 7924 16316 7988
rect 17724 7924 17788 7988
rect 25084 7848 25148 7852
rect 25084 7792 25134 7848
rect 25134 7792 25148 7848
rect 25084 7788 25148 7792
rect 28212 7788 28276 7852
rect 30604 7788 30668 7852
rect 24348 7652 24412 7716
rect 1308 7644 1372 7648
rect 1308 7588 1312 7644
rect 1312 7588 1368 7644
rect 1368 7588 1372 7644
rect 1308 7584 1372 7588
rect 1388 7644 1452 7648
rect 1388 7588 1392 7644
rect 1392 7588 1448 7644
rect 1448 7588 1452 7644
rect 1388 7584 1452 7588
rect 1468 7644 1532 7648
rect 1468 7588 1472 7644
rect 1472 7588 1528 7644
rect 1528 7588 1532 7644
rect 1468 7584 1532 7588
rect 1548 7644 1612 7648
rect 1548 7588 1552 7644
rect 1552 7588 1608 7644
rect 1608 7588 1612 7644
rect 1548 7584 1612 7588
rect 9308 7644 9372 7648
rect 9308 7588 9312 7644
rect 9312 7588 9368 7644
rect 9368 7588 9372 7644
rect 9308 7584 9372 7588
rect 9388 7644 9452 7648
rect 9388 7588 9392 7644
rect 9392 7588 9448 7644
rect 9448 7588 9452 7644
rect 9388 7584 9452 7588
rect 9468 7644 9532 7648
rect 9468 7588 9472 7644
rect 9472 7588 9528 7644
rect 9528 7588 9532 7644
rect 9468 7584 9532 7588
rect 9548 7644 9612 7648
rect 9548 7588 9552 7644
rect 9552 7588 9608 7644
rect 9608 7588 9612 7644
rect 9548 7584 9612 7588
rect 16620 7380 16684 7444
rect 24164 7576 24228 7580
rect 24164 7520 24214 7576
rect 24214 7520 24228 7576
rect 24164 7516 24228 7520
rect 24900 7576 24964 7580
rect 24900 7520 24914 7576
rect 24914 7520 24964 7576
rect 24900 7516 24964 7520
rect 26372 7576 26436 7580
rect 26372 7520 26422 7576
rect 26422 7520 26436 7576
rect 26372 7516 26436 7520
rect 23060 7380 23124 7444
rect 41308 7644 41372 7648
rect 41308 7588 41312 7644
rect 41312 7588 41368 7644
rect 41368 7588 41372 7644
rect 41308 7584 41372 7588
rect 41388 7644 41452 7648
rect 41388 7588 41392 7644
rect 41392 7588 41448 7644
rect 41448 7588 41452 7644
rect 41388 7584 41452 7588
rect 41468 7644 41532 7648
rect 41468 7588 41472 7644
rect 41472 7588 41528 7644
rect 41528 7588 41532 7644
rect 41468 7584 41532 7588
rect 41548 7644 41612 7648
rect 41548 7588 41552 7644
rect 41552 7588 41608 7644
rect 41608 7588 41612 7644
rect 41548 7584 41612 7588
rect 28580 7576 28644 7580
rect 28580 7520 28630 7576
rect 28630 7520 28644 7576
rect 28580 7516 28644 7520
rect 31892 7516 31956 7580
rect 31156 7380 31220 7444
rect 11100 7108 11164 7172
rect 1948 7100 2012 7104
rect 1948 7044 1952 7100
rect 1952 7044 2008 7100
rect 2008 7044 2012 7100
rect 1948 7040 2012 7044
rect 2028 7100 2092 7104
rect 2028 7044 2032 7100
rect 2032 7044 2088 7100
rect 2088 7044 2092 7100
rect 2028 7040 2092 7044
rect 2108 7100 2172 7104
rect 2108 7044 2112 7100
rect 2112 7044 2168 7100
rect 2168 7044 2172 7100
rect 2108 7040 2172 7044
rect 2188 7100 2252 7104
rect 2188 7044 2192 7100
rect 2192 7044 2248 7100
rect 2248 7044 2252 7100
rect 2188 7040 2252 7044
rect 9948 7100 10012 7104
rect 9948 7044 9952 7100
rect 9952 7044 10008 7100
rect 10008 7044 10012 7100
rect 9948 7040 10012 7044
rect 10028 7100 10092 7104
rect 10028 7044 10032 7100
rect 10032 7044 10088 7100
rect 10088 7044 10092 7100
rect 10028 7040 10092 7044
rect 10108 7100 10172 7104
rect 10108 7044 10112 7100
rect 10112 7044 10168 7100
rect 10168 7044 10172 7100
rect 10108 7040 10172 7044
rect 10188 7100 10252 7104
rect 10188 7044 10192 7100
rect 10192 7044 10248 7100
rect 10248 7044 10252 7100
rect 10188 7040 10252 7044
rect 12204 6972 12268 7036
rect 29684 7108 29748 7172
rect 14964 7100 15028 7104
rect 14964 7044 14968 7100
rect 14968 7044 15024 7100
rect 15024 7044 15028 7100
rect 14964 7040 15028 7044
rect 15148 7040 15212 7104
rect 28028 7100 28092 7104
rect 28028 7044 28032 7100
rect 28032 7044 28088 7100
rect 28088 7044 28092 7100
rect 28028 7040 28092 7044
rect 30236 7100 30300 7104
rect 30236 7044 30240 7100
rect 30240 7044 30296 7100
rect 30296 7044 30300 7100
rect 30236 7040 30300 7044
rect 33948 7100 34012 7104
rect 33948 7044 33952 7100
rect 33952 7044 34008 7100
rect 34008 7044 34012 7100
rect 33948 7040 34012 7044
rect 34028 7100 34092 7104
rect 34028 7044 34032 7100
rect 34032 7044 34088 7100
rect 34088 7044 34092 7100
rect 34028 7040 34092 7044
rect 34108 7100 34172 7104
rect 34108 7044 34112 7100
rect 34112 7044 34168 7100
rect 34168 7044 34172 7100
rect 34108 7040 34172 7044
rect 34188 7100 34252 7104
rect 34188 7044 34192 7100
rect 34192 7044 34248 7100
rect 34248 7044 34252 7100
rect 34188 7040 34252 7044
rect 41948 7100 42012 7104
rect 41948 7044 41952 7100
rect 41952 7044 42008 7100
rect 42008 7044 42012 7100
rect 41948 7040 42012 7044
rect 42028 7100 42092 7104
rect 42028 7044 42032 7100
rect 42032 7044 42088 7100
rect 42088 7044 42092 7100
rect 42028 7040 42092 7044
rect 42108 7100 42172 7104
rect 42108 7044 42112 7100
rect 42112 7044 42168 7100
rect 42168 7044 42172 7100
rect 42108 7040 42172 7044
rect 42188 7100 42252 7104
rect 42188 7044 42192 7100
rect 42192 7044 42248 7100
rect 42248 7044 42252 7100
rect 42188 7040 42252 7044
rect 11100 6700 11164 6764
rect 1308 6556 1372 6560
rect 1308 6500 1312 6556
rect 1312 6500 1368 6556
rect 1368 6500 1372 6556
rect 1308 6496 1372 6500
rect 1388 6556 1452 6560
rect 1388 6500 1392 6556
rect 1392 6500 1448 6556
rect 1448 6500 1452 6556
rect 1388 6496 1452 6500
rect 1468 6556 1532 6560
rect 1468 6500 1472 6556
rect 1472 6500 1528 6556
rect 1528 6500 1532 6556
rect 1468 6496 1532 6500
rect 1548 6556 1612 6560
rect 1548 6500 1552 6556
rect 1552 6500 1608 6556
rect 1608 6500 1612 6556
rect 1548 6496 1612 6500
rect 9308 6556 9372 6560
rect 9308 6500 9312 6556
rect 9312 6500 9368 6556
rect 9368 6500 9372 6556
rect 9308 6496 9372 6500
rect 9388 6556 9452 6560
rect 9388 6500 9392 6556
rect 9392 6500 9448 6556
rect 9448 6500 9452 6556
rect 9388 6496 9452 6500
rect 9468 6556 9532 6560
rect 9468 6500 9472 6556
rect 9472 6500 9528 6556
rect 9528 6500 9532 6556
rect 9468 6496 9532 6500
rect 9548 6556 9612 6560
rect 9548 6500 9552 6556
rect 9552 6500 9608 6556
rect 9608 6500 9612 6556
rect 9548 6496 9612 6500
rect 41308 6556 41372 6560
rect 41308 6500 41312 6556
rect 41312 6500 41368 6556
rect 41368 6500 41372 6556
rect 41308 6496 41372 6500
rect 41388 6556 41452 6560
rect 41388 6500 41392 6556
rect 41392 6500 41448 6556
rect 41448 6500 41452 6556
rect 41388 6496 41452 6500
rect 41468 6556 41532 6560
rect 41468 6500 41472 6556
rect 41472 6500 41528 6556
rect 41528 6500 41532 6556
rect 41468 6496 41532 6500
rect 41548 6556 41612 6560
rect 41548 6500 41552 6556
rect 41552 6500 41608 6556
rect 41608 6500 41612 6556
rect 41548 6496 41612 6500
rect 10548 6428 10612 6492
rect 15148 6292 15212 6356
rect 32628 6292 32692 6356
rect 14964 6156 15028 6220
rect 1948 6012 2012 6016
rect 1948 5956 1952 6012
rect 1952 5956 2008 6012
rect 2008 5956 2012 6012
rect 1948 5952 2012 5956
rect 2028 6012 2092 6016
rect 2028 5956 2032 6012
rect 2032 5956 2088 6012
rect 2088 5956 2092 6012
rect 2028 5952 2092 5956
rect 2108 6012 2172 6016
rect 2108 5956 2112 6012
rect 2112 5956 2168 6012
rect 2168 5956 2172 6012
rect 2108 5952 2172 5956
rect 2188 6012 2252 6016
rect 2188 5956 2192 6012
rect 2192 5956 2248 6012
rect 2248 5956 2252 6012
rect 2188 5952 2252 5956
rect 9948 6012 10012 6016
rect 9948 5956 9952 6012
rect 9952 5956 10008 6012
rect 10008 5956 10012 6012
rect 9948 5952 10012 5956
rect 10028 6012 10092 6016
rect 10028 5956 10032 6012
rect 10032 5956 10088 6012
rect 10088 5956 10092 6012
rect 10028 5952 10092 5956
rect 10108 6012 10172 6016
rect 10108 5956 10112 6012
rect 10112 5956 10168 6012
rect 10168 5956 10172 6012
rect 10108 5952 10172 5956
rect 10188 6012 10252 6016
rect 10188 5956 10192 6012
rect 10192 5956 10248 6012
rect 10248 5956 10252 6012
rect 10188 5952 10252 5956
rect 33948 6012 34012 6016
rect 33948 5956 33952 6012
rect 33952 5956 34008 6012
rect 34008 5956 34012 6012
rect 33948 5952 34012 5956
rect 34028 6012 34092 6016
rect 34028 5956 34032 6012
rect 34032 5956 34088 6012
rect 34088 5956 34092 6012
rect 34028 5952 34092 5956
rect 34108 6012 34172 6016
rect 34108 5956 34112 6012
rect 34112 5956 34168 6012
rect 34168 5956 34172 6012
rect 34108 5952 34172 5956
rect 34188 6012 34252 6016
rect 34188 5956 34192 6012
rect 34192 5956 34248 6012
rect 34248 5956 34252 6012
rect 34188 5952 34252 5956
rect 41948 6012 42012 6016
rect 41948 5956 41952 6012
rect 41952 5956 42008 6012
rect 42008 5956 42012 6012
rect 41948 5952 42012 5956
rect 42028 6012 42092 6016
rect 42028 5956 42032 6012
rect 42032 5956 42088 6012
rect 42088 5956 42092 6012
rect 42028 5952 42092 5956
rect 42108 6012 42172 6016
rect 42108 5956 42112 6012
rect 42112 5956 42168 6012
rect 42168 5956 42172 6012
rect 42108 5952 42172 5956
rect 42188 6012 42252 6016
rect 42188 5956 42192 6012
rect 42192 5956 42248 6012
rect 42248 5956 42252 6012
rect 42188 5952 42252 5956
rect 19228 5768 19292 5832
rect 19308 5768 19372 5832
rect 19388 5768 19452 5832
rect 19468 5768 19532 5832
rect 19228 5688 19292 5752
rect 19308 5688 19372 5752
rect 19388 5688 19452 5752
rect 19468 5688 19532 5752
rect 19228 5608 19292 5672
rect 19308 5608 19372 5672
rect 19388 5608 19452 5672
rect 19468 5608 19532 5672
rect 19228 5528 19292 5592
rect 19308 5528 19372 5592
rect 19388 5528 19452 5592
rect 19468 5528 19532 5592
rect 27228 5768 27292 5832
rect 27308 5768 27372 5832
rect 27388 5768 27452 5832
rect 27468 5768 27532 5832
rect 27228 5688 27292 5752
rect 27308 5688 27372 5752
rect 27388 5688 27452 5752
rect 27468 5688 27532 5752
rect 27228 5608 27292 5672
rect 27308 5608 27372 5672
rect 27388 5608 27452 5672
rect 27468 5608 27532 5672
rect 27228 5528 27292 5592
rect 27308 5528 27372 5592
rect 27388 5528 27452 5592
rect 27468 5528 27532 5592
rect 1308 5468 1372 5472
rect 1308 5412 1312 5468
rect 1312 5412 1368 5468
rect 1368 5412 1372 5468
rect 1308 5408 1372 5412
rect 1388 5468 1452 5472
rect 1388 5412 1392 5468
rect 1392 5412 1448 5468
rect 1448 5412 1452 5468
rect 1388 5408 1452 5412
rect 1468 5468 1532 5472
rect 1468 5412 1472 5468
rect 1472 5412 1528 5468
rect 1528 5412 1532 5468
rect 1468 5408 1532 5412
rect 1548 5468 1612 5472
rect 1548 5412 1552 5468
rect 1552 5412 1608 5468
rect 1608 5412 1612 5468
rect 1548 5408 1612 5412
rect 9308 5468 9372 5472
rect 9308 5412 9312 5468
rect 9312 5412 9368 5468
rect 9368 5412 9372 5468
rect 9308 5408 9372 5412
rect 9388 5468 9452 5472
rect 9388 5412 9392 5468
rect 9392 5412 9448 5468
rect 9448 5412 9452 5468
rect 9388 5408 9452 5412
rect 9468 5468 9532 5472
rect 9468 5412 9472 5468
rect 9472 5412 9528 5468
rect 9528 5412 9532 5468
rect 9468 5408 9532 5412
rect 9548 5468 9612 5472
rect 9548 5412 9552 5468
rect 9552 5412 9608 5468
rect 9608 5412 9612 5468
rect 9548 5408 9612 5412
rect 41308 5468 41372 5472
rect 41308 5412 41312 5468
rect 41312 5412 41368 5468
rect 41368 5412 41372 5468
rect 41308 5408 41372 5412
rect 41388 5468 41452 5472
rect 41388 5412 41392 5468
rect 41392 5412 41448 5468
rect 41448 5412 41452 5468
rect 41388 5408 41452 5412
rect 41468 5468 41532 5472
rect 41468 5412 41472 5468
rect 41472 5412 41528 5468
rect 41528 5412 41532 5468
rect 41468 5408 41532 5412
rect 41548 5468 41612 5472
rect 41548 5412 41552 5468
rect 41552 5412 41608 5468
rect 41608 5412 41612 5468
rect 41548 5408 41612 5412
rect 13308 5340 13372 5404
rect 18588 5128 18652 5192
rect 18668 5128 18732 5192
rect 18748 5128 18812 5192
rect 18828 5128 18892 5192
rect 18588 5048 18652 5112
rect 18668 5048 18732 5112
rect 18748 5048 18812 5112
rect 18828 5048 18892 5112
rect 18588 4968 18652 5032
rect 18668 4968 18732 5032
rect 18748 4968 18812 5032
rect 18828 4968 18892 5032
rect 1948 4924 2012 4928
rect 1948 4868 1952 4924
rect 1952 4868 2008 4924
rect 2008 4868 2012 4924
rect 1948 4864 2012 4868
rect 2028 4924 2092 4928
rect 2028 4868 2032 4924
rect 2032 4868 2088 4924
rect 2088 4868 2092 4924
rect 2028 4864 2092 4868
rect 2108 4924 2172 4928
rect 2108 4868 2112 4924
rect 2112 4868 2168 4924
rect 2168 4868 2172 4924
rect 2108 4864 2172 4868
rect 2188 4924 2252 4928
rect 2188 4868 2192 4924
rect 2192 4868 2248 4924
rect 2248 4868 2252 4924
rect 2188 4864 2252 4868
rect 18588 4888 18652 4952
rect 18668 4888 18732 4952
rect 18748 4888 18812 4952
rect 18828 4888 18892 4952
rect 26588 5128 26652 5192
rect 26668 5128 26732 5192
rect 26748 5128 26812 5192
rect 26828 5128 26892 5192
rect 26588 5048 26652 5112
rect 26668 5048 26732 5112
rect 26748 5048 26812 5112
rect 26828 5048 26892 5112
rect 26588 4968 26652 5032
rect 26668 4968 26732 5032
rect 26748 4968 26812 5032
rect 26828 4968 26892 5032
rect 26588 4888 26652 4952
rect 26668 4888 26732 4952
rect 26748 4888 26812 4952
rect 26828 4888 26892 4952
rect 33948 4924 34012 4928
rect 33948 4868 33952 4924
rect 33952 4868 34008 4924
rect 34008 4868 34012 4924
rect 33948 4864 34012 4868
rect 34028 4924 34092 4928
rect 34028 4868 34032 4924
rect 34032 4868 34088 4924
rect 34088 4868 34092 4924
rect 34028 4864 34092 4868
rect 34108 4924 34172 4928
rect 34108 4868 34112 4924
rect 34112 4868 34168 4924
rect 34168 4868 34172 4924
rect 34108 4864 34172 4868
rect 34188 4924 34252 4928
rect 34188 4868 34192 4924
rect 34192 4868 34248 4924
rect 34248 4868 34252 4924
rect 34188 4864 34252 4868
rect 41948 4924 42012 4928
rect 41948 4868 41952 4924
rect 41952 4868 42008 4924
rect 42008 4868 42012 4924
rect 41948 4864 42012 4868
rect 42028 4924 42092 4928
rect 42028 4868 42032 4924
rect 42032 4868 42088 4924
rect 42088 4868 42092 4924
rect 42028 4864 42092 4868
rect 42108 4924 42172 4928
rect 42108 4868 42112 4924
rect 42112 4868 42168 4924
rect 42168 4868 42172 4924
rect 42108 4864 42172 4868
rect 42188 4924 42252 4928
rect 42188 4868 42192 4924
rect 42192 4868 42248 4924
rect 42248 4868 42252 4924
rect 42188 4864 42252 4868
rect 14412 4524 14476 4588
rect 14780 4524 14844 4588
rect 15700 4660 15764 4724
rect 15884 4524 15948 4588
rect 16436 4524 16500 4588
rect 17172 4524 17236 4588
rect 19932 4524 19996 4588
rect 13676 4388 13740 4452
rect 14596 4388 14660 4452
rect 16252 4388 16316 4452
rect 16620 4388 16684 4452
rect 21036 4524 21100 4588
rect 22508 4524 22572 4588
rect 24900 4584 24964 4588
rect 24900 4528 24950 4584
rect 24950 4528 24964 4584
rect 24900 4524 24964 4528
rect 29132 4524 29196 4588
rect 22876 4388 22940 4452
rect 24348 4388 24412 4452
rect 24900 4388 24964 4452
rect 25084 4388 25148 4452
rect 26372 4388 26436 4452
rect 27844 4388 27908 4452
rect 1308 4380 1372 4384
rect 1308 4324 1312 4380
rect 1312 4324 1368 4380
rect 1368 4324 1372 4380
rect 1308 4320 1372 4324
rect 1388 4380 1452 4384
rect 1388 4324 1392 4380
rect 1392 4324 1448 4380
rect 1448 4324 1452 4380
rect 1388 4320 1452 4324
rect 1468 4380 1532 4384
rect 1468 4324 1472 4380
rect 1472 4324 1528 4380
rect 1528 4324 1532 4380
rect 1468 4320 1532 4324
rect 1548 4380 1612 4384
rect 1548 4324 1552 4380
rect 1552 4324 1608 4380
rect 1608 4324 1612 4380
rect 1548 4320 1612 4324
rect 9308 4380 9372 4384
rect 9308 4324 9312 4380
rect 9312 4324 9368 4380
rect 9368 4324 9372 4380
rect 9308 4320 9372 4324
rect 9388 4380 9452 4384
rect 9388 4324 9392 4380
rect 9392 4324 9448 4380
rect 9448 4324 9452 4380
rect 9388 4320 9452 4324
rect 9468 4380 9532 4384
rect 9468 4324 9472 4380
rect 9472 4324 9528 4380
rect 9528 4324 9532 4380
rect 9468 4320 9532 4324
rect 9548 4380 9612 4384
rect 9548 4324 9552 4380
rect 9552 4324 9608 4380
rect 9608 4324 9612 4380
rect 9548 4320 9612 4324
rect 41308 4380 41372 4384
rect 41308 4324 41312 4380
rect 41312 4324 41368 4380
rect 41368 4324 41372 4380
rect 41308 4320 41372 4324
rect 41388 4380 41452 4384
rect 41388 4324 41392 4380
rect 41392 4324 41448 4380
rect 41448 4324 41452 4380
rect 41388 4320 41452 4324
rect 41468 4380 41532 4384
rect 41468 4324 41472 4380
rect 41472 4324 41528 4380
rect 41528 4324 41532 4380
rect 41468 4320 41532 4324
rect 41548 4380 41612 4384
rect 41548 4324 41552 4380
rect 41552 4324 41608 4380
rect 41608 4324 41612 4380
rect 41548 4320 41612 4324
rect 20852 4252 20916 4316
rect 23244 4252 23308 4316
rect 19012 4116 19076 4180
rect 20668 4116 20732 4180
rect 23980 4116 24044 4180
rect 28580 4116 28644 4180
rect 28948 4116 29012 4180
rect 10364 3980 10428 4044
rect 22324 3980 22388 4044
rect 27660 3980 27724 4044
rect 30052 3980 30116 4044
rect 28028 3844 28092 3908
rect 1948 3836 2012 3840
rect 1948 3780 1952 3836
rect 1952 3780 2008 3836
rect 2008 3780 2012 3836
rect 1948 3776 2012 3780
rect 2028 3836 2092 3840
rect 2028 3780 2032 3836
rect 2032 3780 2088 3836
rect 2088 3780 2092 3836
rect 2028 3776 2092 3780
rect 2108 3836 2172 3840
rect 2108 3780 2112 3836
rect 2112 3780 2168 3836
rect 2168 3780 2172 3836
rect 2108 3776 2172 3780
rect 2188 3836 2252 3840
rect 2188 3780 2192 3836
rect 2192 3780 2248 3836
rect 2248 3780 2252 3836
rect 2188 3776 2252 3780
rect 9948 3836 10012 3840
rect 9948 3780 9952 3836
rect 9952 3780 10008 3836
rect 10008 3780 10012 3836
rect 9948 3776 10012 3780
rect 10028 3836 10092 3840
rect 10028 3780 10032 3836
rect 10032 3780 10088 3836
rect 10088 3780 10092 3836
rect 10028 3776 10092 3780
rect 10108 3836 10172 3840
rect 10108 3780 10112 3836
rect 10112 3780 10168 3836
rect 10168 3780 10172 3836
rect 10108 3776 10172 3780
rect 10188 3836 10252 3840
rect 10188 3780 10192 3836
rect 10192 3780 10248 3836
rect 10248 3780 10252 3836
rect 10188 3776 10252 3780
rect 32628 3708 32692 3772
rect 33948 3836 34012 3840
rect 33948 3780 33952 3836
rect 33952 3780 34008 3836
rect 34008 3780 34012 3836
rect 33948 3776 34012 3780
rect 34028 3836 34092 3840
rect 34028 3780 34032 3836
rect 34032 3780 34088 3836
rect 34088 3780 34092 3836
rect 34028 3776 34092 3780
rect 34108 3836 34172 3840
rect 34108 3780 34112 3836
rect 34112 3780 34168 3836
rect 34168 3780 34172 3836
rect 34108 3776 34172 3780
rect 34188 3836 34252 3840
rect 34188 3780 34192 3836
rect 34192 3780 34248 3836
rect 34248 3780 34252 3836
rect 34188 3776 34252 3780
rect 41948 3836 42012 3840
rect 41948 3780 41952 3836
rect 41952 3780 42008 3836
rect 42008 3780 42012 3836
rect 41948 3776 42012 3780
rect 42028 3836 42092 3840
rect 42028 3780 42032 3836
rect 42032 3780 42088 3836
rect 42088 3780 42092 3836
rect 42028 3776 42092 3780
rect 42108 3836 42172 3840
rect 42108 3780 42112 3836
rect 42112 3780 42168 3836
rect 42168 3780 42172 3836
rect 42108 3776 42172 3780
rect 42188 3836 42252 3840
rect 42188 3780 42192 3836
rect 42192 3780 42248 3836
rect 42248 3780 42252 3836
rect 42188 3776 42252 3780
rect 23612 3436 23676 3500
rect 1308 3292 1372 3296
rect 1308 3236 1312 3292
rect 1312 3236 1368 3292
rect 1368 3236 1372 3292
rect 1308 3232 1372 3236
rect 1388 3292 1452 3296
rect 1388 3236 1392 3292
rect 1392 3236 1448 3292
rect 1448 3236 1452 3292
rect 1388 3232 1452 3236
rect 1468 3292 1532 3296
rect 1468 3236 1472 3292
rect 1472 3236 1528 3292
rect 1528 3236 1532 3292
rect 1468 3232 1532 3236
rect 1548 3292 1612 3296
rect 1548 3236 1552 3292
rect 1552 3236 1608 3292
rect 1608 3236 1612 3292
rect 1548 3232 1612 3236
rect 9308 3292 9372 3296
rect 9308 3236 9312 3292
rect 9312 3236 9368 3292
rect 9368 3236 9372 3292
rect 9308 3232 9372 3236
rect 9388 3292 9452 3296
rect 9388 3236 9392 3292
rect 9392 3236 9448 3292
rect 9448 3236 9452 3292
rect 9388 3232 9452 3236
rect 9468 3292 9532 3296
rect 9468 3236 9472 3292
rect 9472 3236 9528 3292
rect 9528 3236 9532 3292
rect 9468 3232 9532 3236
rect 9548 3292 9612 3296
rect 9548 3236 9552 3292
rect 9552 3236 9608 3292
rect 9608 3236 9612 3292
rect 9548 3232 9612 3236
rect 41308 3292 41372 3296
rect 41308 3236 41312 3292
rect 41312 3236 41368 3292
rect 41368 3236 41372 3292
rect 41308 3232 41372 3236
rect 41388 3292 41452 3296
rect 41388 3236 41392 3292
rect 41392 3236 41448 3292
rect 41448 3236 41452 3292
rect 41388 3232 41452 3236
rect 41468 3292 41532 3296
rect 41468 3236 41472 3292
rect 41472 3236 41528 3292
rect 41528 3236 41532 3292
rect 41468 3232 41532 3236
rect 41548 3292 41612 3296
rect 41548 3236 41552 3292
rect 41552 3236 41608 3292
rect 41608 3236 41612 3292
rect 41548 3232 41612 3236
rect 30236 3164 30300 3228
rect 38884 3164 38948 3228
rect 1948 2748 2012 2752
rect 1948 2692 1952 2748
rect 1952 2692 2008 2748
rect 2008 2692 2012 2748
rect 1948 2688 2012 2692
rect 2028 2748 2092 2752
rect 2028 2692 2032 2748
rect 2032 2692 2088 2748
rect 2088 2692 2092 2748
rect 2028 2688 2092 2692
rect 2108 2748 2172 2752
rect 2108 2692 2112 2748
rect 2112 2692 2168 2748
rect 2168 2692 2172 2748
rect 2108 2688 2172 2692
rect 2188 2748 2252 2752
rect 2188 2692 2192 2748
rect 2192 2692 2248 2748
rect 2248 2692 2252 2748
rect 2188 2688 2252 2692
rect 9948 2748 10012 2752
rect 9948 2692 9952 2748
rect 9952 2692 10008 2748
rect 10008 2692 10012 2748
rect 9948 2688 10012 2692
rect 10028 2748 10092 2752
rect 10028 2692 10032 2748
rect 10032 2692 10088 2748
rect 10088 2692 10092 2748
rect 10028 2688 10092 2692
rect 10108 2748 10172 2752
rect 10108 2692 10112 2748
rect 10112 2692 10168 2748
rect 10168 2692 10172 2748
rect 10108 2688 10172 2692
rect 10188 2748 10252 2752
rect 10188 2692 10192 2748
rect 10192 2692 10248 2748
rect 10248 2692 10252 2748
rect 10188 2688 10252 2692
rect 33948 2748 34012 2752
rect 33948 2692 33952 2748
rect 33952 2692 34008 2748
rect 34008 2692 34012 2748
rect 33948 2688 34012 2692
rect 34028 2748 34092 2752
rect 34028 2692 34032 2748
rect 34032 2692 34088 2748
rect 34088 2692 34092 2748
rect 34028 2688 34092 2692
rect 34108 2748 34172 2752
rect 34108 2692 34112 2748
rect 34112 2692 34168 2748
rect 34168 2692 34172 2748
rect 34108 2688 34172 2692
rect 34188 2748 34252 2752
rect 34188 2692 34192 2748
rect 34192 2692 34248 2748
rect 34248 2692 34252 2748
rect 34188 2688 34252 2692
rect 41948 2748 42012 2752
rect 41948 2692 41952 2748
rect 41952 2692 42008 2748
rect 42008 2692 42012 2748
rect 41948 2688 42012 2692
rect 42028 2748 42092 2752
rect 42028 2692 42032 2748
rect 42032 2692 42088 2748
rect 42088 2692 42092 2748
rect 42028 2688 42092 2692
rect 42108 2748 42172 2752
rect 42108 2692 42112 2748
rect 42112 2692 42168 2748
rect 42168 2692 42172 2748
rect 42108 2688 42172 2692
rect 42188 2748 42252 2752
rect 42188 2692 42192 2748
rect 42192 2692 42248 2748
rect 42248 2692 42252 2748
rect 42188 2688 42252 2692
rect 16804 2680 16868 2684
rect 16804 2624 16854 2680
rect 16854 2624 16868 2680
rect 16804 2620 16868 2624
rect 28212 2620 28276 2684
rect 16988 2484 17052 2548
rect 29684 2484 29748 2548
rect 38700 2544 38764 2548
rect 38700 2488 38750 2544
rect 38750 2488 38764 2544
rect 38700 2484 38764 2488
rect 1308 2204 1372 2208
rect 1308 2148 1312 2204
rect 1312 2148 1368 2204
rect 1368 2148 1372 2204
rect 1308 2144 1372 2148
rect 1388 2204 1452 2208
rect 1388 2148 1392 2204
rect 1392 2148 1448 2204
rect 1448 2148 1452 2204
rect 1388 2144 1452 2148
rect 1468 2204 1532 2208
rect 1468 2148 1472 2204
rect 1472 2148 1528 2204
rect 1528 2148 1532 2204
rect 1468 2144 1532 2148
rect 1548 2204 1612 2208
rect 1548 2148 1552 2204
rect 1552 2148 1608 2204
rect 1608 2148 1612 2204
rect 1548 2144 1612 2148
rect 9308 2204 9372 2208
rect 9308 2148 9312 2204
rect 9312 2148 9368 2204
rect 9368 2148 9372 2204
rect 9308 2144 9372 2148
rect 9388 2204 9452 2208
rect 9388 2148 9392 2204
rect 9392 2148 9448 2204
rect 9448 2148 9452 2204
rect 9388 2144 9452 2148
rect 9468 2204 9532 2208
rect 9468 2148 9472 2204
rect 9472 2148 9528 2204
rect 9528 2148 9532 2204
rect 9468 2144 9532 2148
rect 9548 2204 9612 2208
rect 9548 2148 9552 2204
rect 9552 2148 9608 2204
rect 9608 2148 9612 2204
rect 9548 2144 9612 2148
rect 17308 2204 17372 2208
rect 17308 2148 17312 2204
rect 17312 2148 17368 2204
rect 17368 2148 17372 2204
rect 17308 2144 17372 2148
rect 17388 2204 17452 2208
rect 17388 2148 17392 2204
rect 17392 2148 17448 2204
rect 17448 2148 17452 2204
rect 17388 2144 17452 2148
rect 17468 2204 17532 2208
rect 17468 2148 17472 2204
rect 17472 2148 17528 2204
rect 17528 2148 17532 2204
rect 17468 2144 17532 2148
rect 17548 2204 17612 2208
rect 17548 2148 17552 2204
rect 17552 2148 17608 2204
rect 17608 2148 17612 2204
rect 17548 2144 17612 2148
rect 25308 2204 25372 2208
rect 25308 2148 25312 2204
rect 25312 2148 25368 2204
rect 25368 2148 25372 2204
rect 25308 2144 25372 2148
rect 25388 2204 25452 2208
rect 25388 2148 25392 2204
rect 25392 2148 25448 2204
rect 25448 2148 25452 2204
rect 25388 2144 25452 2148
rect 25468 2204 25532 2208
rect 25468 2148 25472 2204
rect 25472 2148 25528 2204
rect 25528 2148 25532 2204
rect 25468 2144 25532 2148
rect 25548 2204 25612 2208
rect 25548 2148 25552 2204
rect 25552 2148 25608 2204
rect 25608 2148 25612 2204
rect 25548 2144 25612 2148
rect 33308 2204 33372 2208
rect 33308 2148 33312 2204
rect 33312 2148 33368 2204
rect 33368 2148 33372 2204
rect 33308 2144 33372 2148
rect 33388 2204 33452 2208
rect 33388 2148 33392 2204
rect 33392 2148 33448 2204
rect 33448 2148 33452 2204
rect 33388 2144 33452 2148
rect 33468 2204 33532 2208
rect 33468 2148 33472 2204
rect 33472 2148 33528 2204
rect 33528 2148 33532 2204
rect 33468 2144 33532 2148
rect 33548 2204 33612 2208
rect 33548 2148 33552 2204
rect 33552 2148 33608 2204
rect 33608 2148 33612 2204
rect 33548 2144 33612 2148
rect 41308 2204 41372 2208
rect 41308 2148 41312 2204
rect 41312 2148 41368 2204
rect 41368 2148 41372 2204
rect 41308 2144 41372 2148
rect 41388 2204 41452 2208
rect 41388 2148 41392 2204
rect 41392 2148 41448 2204
rect 41448 2148 41452 2204
rect 41388 2144 41452 2148
rect 41468 2204 41532 2208
rect 41468 2148 41472 2204
rect 41472 2148 41528 2204
rect 41528 2148 41532 2204
rect 41468 2144 41532 2148
rect 41548 2204 41612 2208
rect 41548 2148 41552 2204
rect 41552 2148 41608 2204
rect 41608 2148 41612 2204
rect 41548 2144 41612 2148
rect 23796 1940 23860 2004
rect 31156 1940 31220 2004
rect 24164 1804 24228 1868
rect 24900 1804 24964 1868
rect 38700 1864 38764 1868
rect 38700 1808 38714 1864
rect 38714 1808 38764 1864
rect 38700 1804 38764 1808
rect 38884 1864 38948 1868
rect 38884 1808 38934 1864
rect 38934 1808 38948 1864
rect 38884 1804 38948 1808
rect 31892 1668 31956 1732
rect 1948 1660 2012 1664
rect 1948 1604 1952 1660
rect 1952 1604 2008 1660
rect 2008 1604 2012 1660
rect 1948 1600 2012 1604
rect 2028 1660 2092 1664
rect 2028 1604 2032 1660
rect 2032 1604 2088 1660
rect 2088 1604 2092 1660
rect 2028 1600 2092 1604
rect 2108 1660 2172 1664
rect 2108 1604 2112 1660
rect 2112 1604 2168 1660
rect 2168 1604 2172 1660
rect 2108 1600 2172 1604
rect 2188 1660 2252 1664
rect 2188 1604 2192 1660
rect 2192 1604 2248 1660
rect 2248 1604 2252 1660
rect 2188 1600 2252 1604
rect 9948 1660 10012 1664
rect 9948 1604 9952 1660
rect 9952 1604 10008 1660
rect 10008 1604 10012 1660
rect 9948 1600 10012 1604
rect 10028 1660 10092 1664
rect 10028 1604 10032 1660
rect 10032 1604 10088 1660
rect 10088 1604 10092 1660
rect 10028 1600 10092 1604
rect 10108 1660 10172 1664
rect 10108 1604 10112 1660
rect 10112 1604 10168 1660
rect 10168 1604 10172 1660
rect 10108 1600 10172 1604
rect 10188 1660 10252 1664
rect 10188 1604 10192 1660
rect 10192 1604 10248 1660
rect 10248 1604 10252 1660
rect 10188 1600 10252 1604
rect 17948 1660 18012 1664
rect 17948 1604 17952 1660
rect 17952 1604 18008 1660
rect 18008 1604 18012 1660
rect 17948 1600 18012 1604
rect 18028 1660 18092 1664
rect 18028 1604 18032 1660
rect 18032 1604 18088 1660
rect 18088 1604 18092 1660
rect 18028 1600 18092 1604
rect 18108 1660 18172 1664
rect 18108 1604 18112 1660
rect 18112 1604 18168 1660
rect 18168 1604 18172 1660
rect 18108 1600 18172 1604
rect 18188 1660 18252 1664
rect 18188 1604 18192 1660
rect 18192 1604 18248 1660
rect 18248 1604 18252 1660
rect 18188 1600 18252 1604
rect 25948 1660 26012 1664
rect 25948 1604 25952 1660
rect 25952 1604 26008 1660
rect 26008 1604 26012 1660
rect 25948 1600 26012 1604
rect 26028 1660 26092 1664
rect 26028 1604 26032 1660
rect 26032 1604 26088 1660
rect 26088 1604 26092 1660
rect 26028 1600 26092 1604
rect 26108 1660 26172 1664
rect 26108 1604 26112 1660
rect 26112 1604 26168 1660
rect 26168 1604 26172 1660
rect 26108 1600 26172 1604
rect 26188 1660 26252 1664
rect 26188 1604 26192 1660
rect 26192 1604 26248 1660
rect 26248 1604 26252 1660
rect 26188 1600 26252 1604
rect 33948 1660 34012 1664
rect 33948 1604 33952 1660
rect 33952 1604 34008 1660
rect 34008 1604 34012 1660
rect 33948 1600 34012 1604
rect 34028 1660 34092 1664
rect 34028 1604 34032 1660
rect 34032 1604 34088 1660
rect 34088 1604 34092 1660
rect 34028 1600 34092 1604
rect 34108 1660 34172 1664
rect 34108 1604 34112 1660
rect 34112 1604 34168 1660
rect 34168 1604 34172 1660
rect 34108 1600 34172 1604
rect 34188 1660 34252 1664
rect 34188 1604 34192 1660
rect 34192 1604 34248 1660
rect 34248 1604 34252 1660
rect 34188 1600 34252 1604
rect 41948 1660 42012 1664
rect 41948 1604 41952 1660
rect 41952 1604 42008 1660
rect 42008 1604 42012 1660
rect 41948 1600 42012 1604
rect 42028 1660 42092 1664
rect 42028 1604 42032 1660
rect 42032 1604 42088 1660
rect 42088 1604 42092 1660
rect 42028 1600 42092 1604
rect 42108 1660 42172 1664
rect 42108 1604 42112 1660
rect 42112 1604 42168 1660
rect 42168 1604 42172 1660
rect 42108 1600 42172 1604
rect 42188 1660 42252 1664
rect 42188 1604 42192 1660
rect 42192 1604 42248 1660
rect 42248 1604 42252 1660
rect 42188 1600 42252 1604
rect 14044 1260 14108 1324
rect 15516 1260 15580 1324
rect 17724 1260 17788 1324
rect 19748 1260 19812 1324
rect 21956 1260 22020 1324
rect 23060 1260 23124 1324
rect 24532 1260 24596 1324
rect 24716 1260 24780 1324
rect 28396 1260 28460 1324
rect 30420 1320 30484 1324
rect 30420 1264 30434 1320
rect 30434 1264 30484 1320
rect 30420 1260 30484 1264
rect 30604 1260 30668 1324
rect 30972 1320 31036 1324
rect 30972 1264 30986 1320
rect 30986 1264 31036 1320
rect 30972 1260 31036 1264
rect 32996 1320 33060 1324
rect 32996 1264 33010 1320
rect 33010 1264 33060 1320
rect 32996 1260 33060 1264
rect 15332 1124 15396 1188
rect 20300 1124 20364 1188
rect 30788 1124 30852 1188
rect 1308 1116 1372 1120
rect 1308 1060 1312 1116
rect 1312 1060 1368 1116
rect 1368 1060 1372 1116
rect 1308 1056 1372 1060
rect 1388 1116 1452 1120
rect 1388 1060 1392 1116
rect 1392 1060 1448 1116
rect 1448 1060 1452 1116
rect 1388 1056 1452 1060
rect 1468 1116 1532 1120
rect 1468 1060 1472 1116
rect 1472 1060 1528 1116
rect 1528 1060 1532 1116
rect 1468 1056 1532 1060
rect 1548 1116 1612 1120
rect 1548 1060 1552 1116
rect 1552 1060 1608 1116
rect 1608 1060 1612 1116
rect 1548 1056 1612 1060
rect 9308 1116 9372 1120
rect 9308 1060 9312 1116
rect 9312 1060 9368 1116
rect 9368 1060 9372 1116
rect 9308 1056 9372 1060
rect 9388 1116 9452 1120
rect 9388 1060 9392 1116
rect 9392 1060 9448 1116
rect 9448 1060 9452 1116
rect 9388 1056 9452 1060
rect 9468 1116 9532 1120
rect 9468 1060 9472 1116
rect 9472 1060 9528 1116
rect 9528 1060 9532 1116
rect 9468 1056 9532 1060
rect 9548 1116 9612 1120
rect 9548 1060 9552 1116
rect 9552 1060 9608 1116
rect 9608 1060 9612 1116
rect 9548 1056 9612 1060
rect 17308 1116 17372 1120
rect 17308 1060 17312 1116
rect 17312 1060 17368 1116
rect 17368 1060 17372 1116
rect 17308 1056 17372 1060
rect 17388 1116 17452 1120
rect 17388 1060 17392 1116
rect 17392 1060 17448 1116
rect 17448 1060 17452 1116
rect 17388 1056 17452 1060
rect 17468 1116 17532 1120
rect 17468 1060 17472 1116
rect 17472 1060 17528 1116
rect 17528 1060 17532 1116
rect 17468 1056 17532 1060
rect 17548 1116 17612 1120
rect 17548 1060 17552 1116
rect 17552 1060 17608 1116
rect 17608 1060 17612 1116
rect 17548 1056 17612 1060
rect 25308 1116 25372 1120
rect 25308 1060 25312 1116
rect 25312 1060 25368 1116
rect 25368 1060 25372 1116
rect 25308 1056 25372 1060
rect 25388 1116 25452 1120
rect 25388 1060 25392 1116
rect 25392 1060 25448 1116
rect 25448 1060 25452 1116
rect 25388 1056 25452 1060
rect 25468 1116 25532 1120
rect 25468 1060 25472 1116
rect 25472 1060 25528 1116
rect 25528 1060 25532 1116
rect 25468 1056 25532 1060
rect 25548 1116 25612 1120
rect 25548 1060 25552 1116
rect 25552 1060 25608 1116
rect 25608 1060 25612 1116
rect 25548 1056 25612 1060
rect 33308 1116 33372 1120
rect 33308 1060 33312 1116
rect 33312 1060 33368 1116
rect 33368 1060 33372 1116
rect 33308 1056 33372 1060
rect 33388 1116 33452 1120
rect 33388 1060 33392 1116
rect 33392 1060 33448 1116
rect 33448 1060 33452 1116
rect 33388 1056 33452 1060
rect 33468 1116 33532 1120
rect 33468 1060 33472 1116
rect 33472 1060 33528 1116
rect 33528 1060 33532 1116
rect 33468 1056 33532 1060
rect 33548 1116 33612 1120
rect 33548 1060 33552 1116
rect 33552 1060 33608 1116
rect 33608 1060 33612 1116
rect 33548 1056 33612 1060
rect 41308 1116 41372 1120
rect 41308 1060 41312 1116
rect 41312 1060 41368 1116
rect 41368 1060 41372 1116
rect 41308 1056 41372 1060
rect 41388 1116 41452 1120
rect 41388 1060 41392 1116
rect 41392 1060 41448 1116
rect 41448 1060 41452 1116
rect 41388 1056 41452 1060
rect 41468 1116 41532 1120
rect 41468 1060 41472 1116
rect 41472 1060 41528 1116
rect 41528 1060 41532 1116
rect 41468 1056 41532 1060
rect 41548 1116 41612 1120
rect 41548 1060 41552 1116
rect 41552 1060 41608 1116
rect 41608 1060 41612 1116
rect 41548 1056 41612 1060
rect 16068 988 16132 1052
rect 21404 988 21468 1052
rect 23428 988 23492 1052
rect 20116 852 20180 916
rect 21588 716 21652 780
rect 1948 572 2012 576
rect 1948 516 1952 572
rect 1952 516 2008 572
rect 2008 516 2012 572
rect 1948 512 2012 516
rect 2028 572 2092 576
rect 2028 516 2032 572
rect 2032 516 2088 572
rect 2088 516 2092 572
rect 2028 512 2092 516
rect 2108 572 2172 576
rect 2108 516 2112 572
rect 2112 516 2168 572
rect 2168 516 2172 572
rect 2108 512 2172 516
rect 2188 572 2252 576
rect 2188 516 2192 572
rect 2192 516 2248 572
rect 2248 516 2252 572
rect 2188 512 2252 516
rect 9948 572 10012 576
rect 9948 516 9952 572
rect 9952 516 10008 572
rect 10008 516 10012 572
rect 9948 512 10012 516
rect 10028 572 10092 576
rect 10028 516 10032 572
rect 10032 516 10088 572
rect 10088 516 10092 572
rect 10028 512 10092 516
rect 10108 572 10172 576
rect 10108 516 10112 572
rect 10112 516 10168 572
rect 10168 516 10172 572
rect 10108 512 10172 516
rect 10188 572 10252 576
rect 10188 516 10192 572
rect 10192 516 10248 572
rect 10248 516 10252 572
rect 10188 512 10252 516
rect 17948 572 18012 576
rect 17948 516 17952 572
rect 17952 516 18008 572
rect 18008 516 18012 572
rect 17948 512 18012 516
rect 18028 572 18092 576
rect 18028 516 18032 572
rect 18032 516 18088 572
rect 18088 516 18092 572
rect 18028 512 18092 516
rect 18108 572 18172 576
rect 18108 516 18112 572
rect 18112 516 18168 572
rect 18168 516 18172 572
rect 18108 512 18172 516
rect 18188 572 18252 576
rect 18188 516 18192 572
rect 18192 516 18248 572
rect 18248 516 18252 572
rect 18188 512 18252 516
rect 25948 572 26012 576
rect 25948 516 25952 572
rect 25952 516 26008 572
rect 26008 516 26012 572
rect 25948 512 26012 516
rect 26028 572 26092 576
rect 26028 516 26032 572
rect 26032 516 26088 572
rect 26088 516 26092 572
rect 26028 512 26092 516
rect 26108 572 26172 576
rect 26108 516 26112 572
rect 26112 516 26168 572
rect 26168 516 26172 572
rect 26108 512 26172 516
rect 26188 572 26252 576
rect 26188 516 26192 572
rect 26192 516 26248 572
rect 26248 516 26252 572
rect 26188 512 26252 516
rect 33948 572 34012 576
rect 33948 516 33952 572
rect 33952 516 34008 572
rect 34008 516 34012 572
rect 33948 512 34012 516
rect 34028 572 34092 576
rect 34028 516 34032 572
rect 34032 516 34088 572
rect 34088 516 34092 572
rect 34028 512 34092 516
rect 34108 572 34172 576
rect 34108 516 34112 572
rect 34112 516 34168 572
rect 34168 516 34172 572
rect 34108 512 34172 516
rect 34188 572 34252 576
rect 34188 516 34192 572
rect 34192 516 34248 572
rect 34248 516 34252 572
rect 34188 512 34252 516
rect 41948 572 42012 576
rect 41948 516 41952 572
rect 41952 516 42008 572
rect 42008 516 42012 572
rect 41948 512 42012 516
rect 42028 572 42092 576
rect 42028 516 42032 572
rect 42032 516 42088 572
rect 42088 516 42092 572
rect 42028 512 42092 516
rect 42108 572 42172 576
rect 42108 516 42112 572
rect 42112 516 42168 572
rect 42168 516 42172 572
rect 42108 512 42172 516
rect 42188 572 42252 576
rect 42188 516 42192 572
rect 42192 516 42248 572
rect 42248 516 42252 572
rect 42188 512 42252 516
<< metal4 >>
rect 1300 10912 1620 11472
rect 1300 10848 1308 10912
rect 1372 10848 1388 10912
rect 1452 10848 1468 10912
rect 1532 10848 1548 10912
rect 1612 10848 1620 10912
rect 1300 9824 1620 10848
rect 1300 9760 1308 9824
rect 1372 9760 1388 9824
rect 1452 9760 1468 9824
rect 1532 9760 1548 9824
rect 1612 9760 1620 9824
rect 1300 8736 1620 9760
rect 1300 8672 1308 8736
rect 1372 8672 1388 8736
rect 1452 8672 1468 8736
rect 1532 8672 1548 8736
rect 1612 8672 1620 8736
rect 1300 7648 1620 8672
rect 1300 7584 1308 7648
rect 1372 7584 1388 7648
rect 1452 7584 1468 7648
rect 1532 7584 1548 7648
rect 1612 7584 1620 7648
rect 1300 6560 1620 7584
rect 1300 6496 1308 6560
rect 1372 6496 1388 6560
rect 1452 6496 1468 6560
rect 1532 6496 1548 6560
rect 1612 6496 1620 6560
rect 1300 5472 1620 6496
rect 1300 5408 1308 5472
rect 1372 5408 1388 5472
rect 1452 5408 1468 5472
rect 1532 5408 1548 5472
rect 1612 5408 1620 5472
rect 1300 4384 1620 5408
rect 1300 4320 1308 4384
rect 1372 4320 1388 4384
rect 1452 4320 1468 4384
rect 1532 4320 1548 4384
rect 1612 4320 1620 4384
rect 1300 3296 1620 4320
rect 1300 3232 1308 3296
rect 1372 3232 1388 3296
rect 1452 3232 1468 3296
rect 1532 3232 1548 3296
rect 1612 3232 1620 3296
rect 1300 2208 1620 3232
rect 1300 2144 1308 2208
rect 1372 2144 1388 2208
rect 1452 2144 1468 2208
rect 1532 2144 1548 2208
rect 1612 2144 1620 2208
rect 1300 1120 1620 2144
rect 1300 1056 1308 1120
rect 1372 1056 1388 1120
rect 1452 1056 1468 1120
rect 1532 1056 1548 1120
rect 1612 1056 1620 1120
rect 1300 496 1620 1056
rect 1940 11456 2260 11472
rect 1940 11392 1948 11456
rect 2012 11392 2028 11456
rect 2092 11392 2108 11456
rect 2172 11392 2188 11456
rect 2252 11392 2260 11456
rect 1940 10368 2260 11392
rect 1940 10304 1948 10368
rect 2012 10304 2028 10368
rect 2092 10304 2108 10368
rect 2172 10304 2188 10368
rect 2252 10304 2260 10368
rect 1940 9280 2260 10304
rect 1940 9216 1948 9280
rect 2012 9216 2028 9280
rect 2092 9216 2108 9280
rect 2172 9216 2188 9280
rect 2252 9216 2260 9280
rect 1940 8192 2260 9216
rect 1940 8128 1948 8192
rect 2012 8128 2028 8192
rect 2092 8128 2108 8192
rect 2172 8128 2188 8192
rect 2252 8128 2260 8192
rect 1940 7104 2260 8128
rect 1940 7040 1948 7104
rect 2012 7040 2028 7104
rect 2092 7040 2108 7104
rect 2172 7040 2188 7104
rect 2252 7040 2260 7104
rect 1940 6016 2260 7040
rect 1940 5952 1948 6016
rect 2012 5952 2028 6016
rect 2092 5952 2108 6016
rect 2172 5952 2188 6016
rect 2252 5952 2260 6016
rect 1940 4928 2260 5952
rect 1940 4864 1948 4928
rect 2012 4864 2028 4928
rect 2092 4864 2108 4928
rect 2172 4864 2188 4928
rect 2252 4864 2260 4928
rect 1940 3840 2260 4864
rect 1940 3776 1948 3840
rect 2012 3776 2028 3840
rect 2092 3776 2108 3840
rect 2172 3776 2188 3840
rect 2252 3776 2260 3840
rect 1940 2752 2260 3776
rect 1940 2688 1948 2752
rect 2012 2688 2028 2752
rect 2092 2688 2108 2752
rect 2172 2688 2188 2752
rect 2252 2688 2260 2752
rect 1940 1664 2260 2688
rect 1940 1600 1948 1664
rect 2012 1600 2028 1664
rect 2092 1600 2108 1664
rect 2172 1600 2188 1664
rect 2252 1600 2260 1664
rect 1940 576 2260 1600
rect 1940 512 1948 576
rect 2012 512 2028 576
rect 2092 512 2108 576
rect 2172 512 2188 576
rect 2252 512 2260 576
rect 1940 496 2260 512
rect 9300 10912 9620 11472
rect 9300 10848 9308 10912
rect 9372 10848 9388 10912
rect 9452 10848 9468 10912
rect 9532 10848 9548 10912
rect 9612 10848 9620 10912
rect 9300 9824 9620 10848
rect 9300 9760 9308 9824
rect 9372 9760 9388 9824
rect 9452 9760 9468 9824
rect 9532 9760 9548 9824
rect 9612 9760 9620 9824
rect 9300 8736 9620 9760
rect 9300 8672 9308 8736
rect 9372 8672 9388 8736
rect 9452 8672 9468 8736
rect 9532 8672 9548 8736
rect 9612 8672 9620 8736
rect 9300 7648 9620 8672
rect 9940 11456 10260 11472
rect 9940 11392 9948 11456
rect 10012 11392 10028 11456
rect 10092 11392 10108 11456
rect 10172 11392 10188 11456
rect 10252 11392 10260 11456
rect 9940 10368 10260 11392
rect 9940 10304 9948 10368
rect 10012 10304 10028 10368
rect 10092 10304 10108 10368
rect 10172 10304 10188 10368
rect 10252 10304 10260 10368
rect 9940 9280 10260 10304
rect 17300 10912 17620 11472
rect 17300 10848 17308 10912
rect 17372 10848 17388 10912
rect 17452 10848 17468 10912
rect 17532 10848 17548 10912
rect 17612 10848 17620 10912
rect 17300 9824 17620 10848
rect 17300 9760 17308 9824
rect 17372 9760 17388 9824
rect 17452 9760 17468 9824
rect 17532 9760 17548 9824
rect 17612 9760 17620 9824
rect 14043 9484 14109 9485
rect 14043 9420 14044 9484
rect 14108 9420 14109 9484
rect 14043 9419 14109 9420
rect 14595 9484 14661 9485
rect 14595 9420 14596 9484
rect 14660 9420 14661 9484
rect 14595 9419 14661 9420
rect 9940 9216 9948 9280
rect 10012 9216 10028 9280
rect 10092 9216 10108 9280
rect 10172 9216 10188 9280
rect 10252 9216 10260 9280
rect 9811 8668 9877 8669
rect 9811 8604 9812 8668
rect 9876 8604 9877 8668
rect 9811 8603 9877 8604
rect 9814 8125 9874 8603
rect 9940 8192 10260 9216
rect 13675 8940 13741 8941
rect 13675 8876 13676 8940
rect 13740 8876 13741 8940
rect 13675 8875 13741 8876
rect 10547 8804 10613 8805
rect 10547 8740 10548 8804
rect 10612 8740 10613 8804
rect 10547 8739 10613 8740
rect 10363 8668 10429 8669
rect 10363 8604 10364 8668
rect 10428 8604 10429 8668
rect 10363 8603 10429 8604
rect 9940 8128 9948 8192
rect 10012 8128 10028 8192
rect 10092 8128 10108 8192
rect 10172 8128 10188 8192
rect 10252 8128 10260 8192
rect 9811 8124 9877 8125
rect 9811 8060 9812 8124
rect 9876 8060 9877 8124
rect 9811 8059 9877 8060
rect 9300 7584 9308 7648
rect 9372 7584 9388 7648
rect 9452 7584 9468 7648
rect 9532 7584 9548 7648
rect 9612 7584 9620 7648
rect 9300 6560 9620 7584
rect 9300 6496 9308 6560
rect 9372 6496 9388 6560
rect 9452 6496 9468 6560
rect 9532 6496 9548 6560
rect 9612 6496 9620 6560
rect 9300 5472 9620 6496
rect 9300 5408 9308 5472
rect 9372 5408 9388 5472
rect 9452 5408 9468 5472
rect 9532 5408 9548 5472
rect 9612 5408 9620 5472
rect 9300 4384 9620 5408
rect 9300 4320 9308 4384
rect 9372 4320 9388 4384
rect 9452 4320 9468 4384
rect 9532 4320 9548 4384
rect 9612 4320 9620 4384
rect 9300 3296 9620 4320
rect 9300 3232 9308 3296
rect 9372 3232 9388 3296
rect 9452 3232 9468 3296
rect 9532 3232 9548 3296
rect 9612 3232 9620 3296
rect 9300 2208 9620 3232
rect 9300 2144 9308 2208
rect 9372 2144 9388 2208
rect 9452 2144 9468 2208
rect 9532 2144 9548 2208
rect 9612 2144 9620 2208
rect 9300 1120 9620 2144
rect 9300 1056 9308 1120
rect 9372 1056 9388 1120
rect 9452 1056 9468 1120
rect 9532 1056 9548 1120
rect 9612 1056 9620 1120
rect 9300 496 9620 1056
rect 9940 7104 10260 8128
rect 9940 7040 9948 7104
rect 10012 7040 10028 7104
rect 10092 7040 10108 7104
rect 10172 7040 10188 7104
rect 10252 7040 10260 7104
rect 9940 6016 10260 7040
rect 9940 5952 9948 6016
rect 10012 5952 10028 6016
rect 10092 5952 10108 6016
rect 10172 5952 10188 6016
rect 10252 5952 10260 6016
rect 9940 3840 10260 5952
rect 10366 4045 10426 8603
rect 10550 6493 10610 8739
rect 13307 8396 13373 8397
rect 13307 8332 13308 8396
rect 13372 8332 13373 8396
rect 13307 8331 13373 8332
rect 12387 8124 12453 8125
rect 12387 8060 12388 8124
rect 12452 8060 12453 8124
rect 12387 8059 12453 8060
rect 12390 7850 12450 8059
rect 12206 7790 12450 7850
rect 11099 7172 11165 7173
rect 11099 7108 11100 7172
rect 11164 7108 11165 7172
rect 11099 7107 11165 7108
rect 11102 6765 11162 7107
rect 12206 7037 12266 7790
rect 12203 7036 12269 7037
rect 12203 6972 12204 7036
rect 12268 6972 12269 7036
rect 12203 6971 12269 6972
rect 11099 6764 11165 6765
rect 11099 6700 11100 6764
rect 11164 6700 11165 6764
rect 11099 6699 11165 6700
rect 10547 6492 10613 6493
rect 10547 6428 10548 6492
rect 10612 6428 10613 6492
rect 10547 6427 10613 6428
rect 13310 5405 13370 8331
rect 13307 5404 13373 5405
rect 13307 5340 13308 5404
rect 13372 5340 13373 5404
rect 13307 5339 13373 5340
rect 13678 4453 13738 8875
rect 13675 4452 13741 4453
rect 13675 4388 13676 4452
rect 13740 4388 13741 4452
rect 13675 4387 13741 4388
rect 10363 4044 10429 4045
rect 10363 3980 10364 4044
rect 10428 3980 10429 4044
rect 10363 3979 10429 3980
rect 9940 3776 9948 3840
rect 10012 3776 10028 3840
rect 10092 3776 10108 3840
rect 10172 3776 10188 3840
rect 10252 3776 10260 3840
rect 9940 2752 10260 3776
rect 9940 2688 9948 2752
rect 10012 2688 10028 2752
rect 10092 2688 10108 2752
rect 10172 2688 10188 2752
rect 10252 2688 10260 2752
rect 9940 1664 10260 2688
rect 9940 1600 9948 1664
rect 10012 1600 10028 1664
rect 10092 1600 10108 1664
rect 10172 1600 10188 1664
rect 10252 1600 10260 1664
rect 9940 576 10260 1600
rect 14046 1325 14106 9419
rect 14411 9076 14477 9077
rect 14411 9012 14412 9076
rect 14476 9012 14477 9076
rect 14411 9011 14477 9012
rect 14414 4589 14474 9011
rect 14411 4588 14477 4589
rect 14411 4524 14412 4588
rect 14476 4524 14477 4588
rect 14411 4523 14477 4524
rect 14598 4453 14658 9419
rect 16067 8940 16133 8941
rect 16067 8876 16068 8940
rect 16132 8876 16133 8940
rect 16067 8875 16133 8876
rect 16435 8940 16501 8941
rect 16435 8876 16436 8940
rect 16500 8876 16501 8940
rect 16435 8875 16501 8876
rect 15699 8804 15765 8805
rect 15699 8740 15700 8804
rect 15764 8740 15765 8804
rect 15699 8739 15765 8740
rect 15515 8668 15581 8669
rect 15515 8604 15516 8668
rect 15580 8604 15581 8668
rect 15515 8603 15581 8604
rect 14779 8260 14845 8261
rect 14779 8196 14780 8260
rect 14844 8196 14845 8260
rect 14779 8195 14845 8196
rect 15331 8260 15397 8261
rect 15331 8196 15332 8260
rect 15396 8196 15397 8260
rect 15331 8195 15397 8196
rect 14782 4589 14842 8195
rect 14963 7104 15029 7105
rect 14963 7040 14964 7104
rect 15028 7040 15029 7104
rect 14963 7039 15029 7040
rect 15147 7104 15213 7105
rect 15147 7040 15148 7104
rect 15212 7040 15213 7104
rect 15147 7039 15213 7040
rect 14966 6221 15026 7039
rect 15150 6357 15210 7039
rect 15147 6356 15213 6357
rect 15147 6292 15148 6356
rect 15212 6292 15213 6356
rect 15147 6291 15213 6292
rect 14963 6220 15029 6221
rect 14963 6156 14964 6220
rect 15028 6156 15029 6220
rect 14963 6155 15029 6156
rect 14779 4588 14845 4589
rect 14779 4524 14780 4588
rect 14844 4524 14845 4588
rect 14779 4523 14845 4524
rect 14595 4452 14661 4453
rect 14595 4388 14596 4452
rect 14660 4388 14661 4452
rect 14595 4387 14661 4388
rect 14043 1324 14109 1325
rect 14043 1260 14044 1324
rect 14108 1260 14109 1324
rect 14043 1259 14109 1260
rect 15334 1189 15394 8195
rect 15518 1325 15578 8603
rect 15702 4725 15762 8739
rect 16070 8397 16130 8875
rect 16067 8396 16133 8397
rect 16067 8332 16068 8396
rect 16132 8332 16133 8396
rect 16067 8331 16133 8332
rect 15883 8260 15949 8261
rect 15883 8196 15884 8260
rect 15948 8196 15949 8260
rect 15883 8195 15949 8196
rect 15699 4724 15765 4725
rect 15699 4660 15700 4724
rect 15764 4660 15765 4724
rect 15699 4659 15765 4660
rect 15886 4589 15946 8195
rect 15883 4588 15949 4589
rect 15883 4524 15884 4588
rect 15948 4524 15949 4588
rect 15883 4523 15949 4524
rect 15515 1324 15581 1325
rect 15515 1260 15516 1324
rect 15580 1260 15581 1324
rect 15515 1259 15581 1260
rect 15331 1188 15397 1189
rect 15331 1124 15332 1188
rect 15396 1124 15397 1188
rect 15331 1123 15397 1124
rect 16070 1053 16130 8331
rect 16251 7988 16317 7989
rect 16251 7924 16252 7988
rect 16316 7924 16317 7988
rect 16251 7923 16317 7924
rect 16254 4453 16314 7923
rect 16438 4589 16498 8875
rect 16987 8532 17053 8533
rect 16987 8468 16988 8532
rect 17052 8468 17053 8532
rect 16987 8467 17053 8468
rect 16803 8396 16869 8397
rect 16803 8332 16804 8396
rect 16868 8332 16869 8396
rect 16803 8331 16869 8332
rect 16619 7444 16685 7445
rect 16619 7380 16620 7444
rect 16684 7380 16685 7444
rect 16619 7379 16685 7380
rect 16435 4588 16501 4589
rect 16435 4524 16436 4588
rect 16500 4524 16501 4588
rect 16435 4523 16501 4524
rect 16622 4453 16682 7379
rect 16251 4452 16317 4453
rect 16251 4388 16252 4452
rect 16316 4388 16317 4452
rect 16251 4387 16317 4388
rect 16619 4452 16685 4453
rect 16619 4388 16620 4452
rect 16684 4388 16685 4452
rect 16619 4387 16685 4388
rect 16806 2685 16866 8331
rect 16803 2684 16869 2685
rect 16803 2620 16804 2684
rect 16868 2620 16869 2684
rect 16803 2619 16869 2620
rect 16990 2549 17050 8467
rect 17171 8260 17237 8261
rect 17171 8196 17172 8260
rect 17236 8196 17237 8260
rect 17171 8195 17237 8196
rect 17174 4589 17234 8195
rect 17171 4588 17237 4589
rect 17171 4524 17172 4588
rect 17236 4524 17237 4588
rect 17171 4523 17237 4524
rect 16987 2548 17053 2549
rect 16987 2484 16988 2548
rect 17052 2484 17053 2548
rect 16987 2483 17053 2484
rect 17300 2208 17620 9760
rect 17940 11456 18260 11472
rect 17940 11392 17948 11456
rect 18012 11392 18028 11456
rect 18092 11392 18108 11456
rect 18172 11392 18188 11456
rect 18252 11392 18260 11456
rect 17940 10368 18260 11392
rect 17940 10304 17948 10368
rect 18012 10304 18028 10368
rect 18092 10304 18108 10368
rect 18172 10304 18188 10368
rect 18252 10304 18260 10368
rect 17723 7988 17789 7989
rect 17723 7924 17724 7988
rect 17788 7924 17789 7988
rect 17723 7923 17789 7924
rect 17300 2144 17308 2208
rect 17372 2144 17388 2208
rect 17452 2144 17468 2208
rect 17532 2144 17548 2208
rect 17612 2144 17620 2208
rect 17300 1120 17620 2144
rect 17726 1325 17786 7923
rect 17940 1664 18260 10304
rect 17940 1600 17948 1664
rect 18012 1600 18028 1664
rect 18092 1600 18108 1664
rect 18172 1600 18188 1664
rect 18252 1600 18260 1664
rect 17723 1324 17789 1325
rect 17723 1260 17724 1324
rect 17788 1260 17789 1324
rect 17723 1259 17789 1260
rect 17300 1056 17308 1120
rect 17372 1056 17388 1120
rect 17452 1056 17468 1120
rect 17532 1056 17548 1120
rect 17612 1056 17620 1120
rect 16067 1052 16133 1053
rect 16067 988 16068 1052
rect 16132 988 16133 1052
rect 16067 987 16133 988
rect 9940 512 9948 576
rect 10012 512 10028 576
rect 10092 512 10108 576
rect 10172 512 10188 576
rect 10252 512 10260 576
rect 9940 496 10260 512
rect 17300 496 17620 1056
rect 17940 576 18260 1600
rect 17940 512 17948 576
rect 18012 512 18028 576
rect 18092 512 18108 576
rect 18172 512 18188 576
rect 18252 512 18260 576
rect 17940 496 18260 512
rect 18580 5192 18900 11472
rect 19011 8940 19077 8941
rect 19011 8876 19012 8940
rect 19076 8876 19077 8940
rect 19011 8875 19077 8876
rect 18580 5128 18588 5192
rect 18652 5128 18668 5192
rect 18732 5128 18748 5192
rect 18812 5128 18828 5192
rect 18892 5128 18900 5192
rect 18580 5112 18900 5128
rect 18580 5048 18588 5112
rect 18652 5048 18668 5112
rect 18732 5048 18748 5112
rect 18812 5048 18828 5112
rect 18892 5048 18900 5112
rect 18580 5032 18900 5048
rect 18580 4968 18588 5032
rect 18652 4968 18668 5032
rect 18732 4968 18748 5032
rect 18812 4968 18828 5032
rect 18892 4968 18900 5032
rect 18580 4952 18900 4968
rect 18580 4888 18588 4952
rect 18652 4888 18668 4952
rect 18732 4888 18748 4952
rect 18812 4888 18828 4952
rect 18892 4888 18900 4952
rect 18580 496 18900 4888
rect 19014 4181 19074 8875
rect 19220 5832 19540 11472
rect 25300 10912 25620 11472
rect 25300 10848 25308 10912
rect 25372 10848 25388 10912
rect 25452 10848 25468 10912
rect 25532 10848 25548 10912
rect 25612 10848 25620 10912
rect 25300 9824 25620 10848
rect 25300 9760 25308 9824
rect 25372 9760 25388 9824
rect 25452 9760 25468 9824
rect 25532 9760 25548 9824
rect 25612 9760 25620 9824
rect 24531 9756 24597 9757
rect 24531 9692 24532 9756
rect 24596 9692 24597 9756
rect 24531 9691 24597 9692
rect 24715 9756 24781 9757
rect 24715 9692 24716 9756
rect 24780 9692 24781 9756
rect 24715 9691 24781 9692
rect 22323 9348 22389 9349
rect 22323 9284 22324 9348
rect 22388 9284 22389 9348
rect 22323 9283 22389 9284
rect 19747 8940 19813 8941
rect 19747 8876 19748 8940
rect 19812 8876 19813 8940
rect 19747 8875 19813 8876
rect 19931 8940 19997 8941
rect 19931 8876 19932 8940
rect 19996 8876 19997 8940
rect 19931 8875 19997 8876
rect 20299 8940 20365 8941
rect 20299 8876 20300 8940
rect 20364 8876 20365 8940
rect 20299 8875 20365 8876
rect 19220 5768 19228 5832
rect 19292 5768 19308 5832
rect 19372 5768 19388 5832
rect 19452 5768 19468 5832
rect 19532 5768 19540 5832
rect 19220 5752 19540 5768
rect 19220 5688 19228 5752
rect 19292 5688 19308 5752
rect 19372 5688 19388 5752
rect 19452 5688 19468 5752
rect 19532 5688 19540 5752
rect 19220 5672 19540 5688
rect 19220 5608 19228 5672
rect 19292 5608 19308 5672
rect 19372 5608 19388 5672
rect 19452 5608 19468 5672
rect 19532 5608 19540 5672
rect 19220 5592 19540 5608
rect 19220 5528 19228 5592
rect 19292 5528 19308 5592
rect 19372 5528 19388 5592
rect 19452 5528 19468 5592
rect 19532 5528 19540 5592
rect 19011 4180 19077 4181
rect 19011 4116 19012 4180
rect 19076 4116 19077 4180
rect 19011 4115 19077 4116
rect 19220 496 19540 5528
rect 19750 1325 19810 8875
rect 19934 4589 19994 8875
rect 20115 8396 20181 8397
rect 20115 8332 20116 8396
rect 20180 8332 20181 8396
rect 20115 8331 20181 8332
rect 19931 4588 19997 4589
rect 19931 4524 19932 4588
rect 19996 4524 19997 4588
rect 19931 4523 19997 4524
rect 19747 1324 19813 1325
rect 19747 1260 19748 1324
rect 19812 1260 19813 1324
rect 19747 1259 19813 1260
rect 20118 917 20178 8331
rect 20302 1189 20362 8875
rect 20851 8532 20917 8533
rect 20851 8468 20852 8532
rect 20916 8468 20917 8532
rect 20851 8467 20917 8468
rect 21403 8532 21469 8533
rect 21403 8468 21404 8532
rect 21468 8468 21469 8532
rect 21403 8467 21469 8468
rect 20667 8396 20733 8397
rect 20667 8332 20668 8396
rect 20732 8332 20733 8396
rect 20667 8331 20733 8332
rect 20670 4181 20730 8331
rect 20854 4317 20914 8467
rect 21035 8124 21101 8125
rect 21035 8060 21036 8124
rect 21100 8060 21101 8124
rect 21035 8059 21101 8060
rect 21038 4589 21098 8059
rect 21035 4588 21101 4589
rect 21035 4524 21036 4588
rect 21100 4524 21101 4588
rect 21035 4523 21101 4524
rect 20851 4316 20917 4317
rect 20851 4252 20852 4316
rect 20916 4252 20917 4316
rect 20851 4251 20917 4252
rect 20667 4180 20733 4181
rect 20667 4116 20668 4180
rect 20732 4116 20733 4180
rect 20667 4115 20733 4116
rect 20299 1188 20365 1189
rect 20299 1124 20300 1188
rect 20364 1124 20365 1188
rect 20299 1123 20365 1124
rect 21406 1053 21466 8467
rect 21587 8396 21653 8397
rect 21587 8332 21588 8396
rect 21652 8332 21653 8396
rect 21587 8331 21653 8332
rect 21403 1052 21469 1053
rect 21403 988 21404 1052
rect 21468 988 21469 1052
rect 21403 987 21469 988
rect 20115 916 20181 917
rect 20115 852 20116 916
rect 20180 852 20181 916
rect 20115 851 20181 852
rect 21590 781 21650 8331
rect 21955 8124 22021 8125
rect 21955 8060 21956 8124
rect 22020 8060 22021 8124
rect 21955 8059 22021 8060
rect 21958 1325 22018 8059
rect 22326 4045 22386 9283
rect 23243 9212 23309 9213
rect 23243 9148 23244 9212
rect 23308 9148 23309 9212
rect 23243 9147 23309 9148
rect 22507 9076 22573 9077
rect 22507 9012 22508 9076
rect 22572 9012 22573 9076
rect 22507 9011 22573 9012
rect 22510 4589 22570 9011
rect 22875 8396 22941 8397
rect 22875 8332 22876 8396
rect 22940 8332 22941 8396
rect 22875 8331 22941 8332
rect 22507 4588 22573 4589
rect 22507 4524 22508 4588
rect 22572 4524 22573 4588
rect 22507 4523 22573 4524
rect 22878 4453 22938 8331
rect 23059 7444 23125 7445
rect 23059 7380 23060 7444
rect 23124 7380 23125 7444
rect 23059 7379 23125 7380
rect 22875 4452 22941 4453
rect 22875 4388 22876 4452
rect 22940 4388 22941 4452
rect 22875 4387 22941 4388
rect 22323 4044 22389 4045
rect 22323 3980 22324 4044
rect 22388 3980 22389 4044
rect 22323 3979 22389 3980
rect 23062 1325 23122 7379
rect 23246 4317 23306 9147
rect 23611 8940 23677 8941
rect 23611 8876 23612 8940
rect 23676 8876 23677 8940
rect 23611 8875 23677 8876
rect 23427 8260 23493 8261
rect 23427 8196 23428 8260
rect 23492 8196 23493 8260
rect 23427 8195 23493 8196
rect 23243 4316 23309 4317
rect 23243 4252 23244 4316
rect 23308 4252 23309 4316
rect 23243 4251 23309 4252
rect 21955 1324 22021 1325
rect 21955 1260 21956 1324
rect 22020 1260 22021 1324
rect 21955 1259 22021 1260
rect 23059 1324 23125 1325
rect 23059 1260 23060 1324
rect 23124 1260 23125 1324
rect 23059 1259 23125 1260
rect 23430 1053 23490 8195
rect 23614 3501 23674 8875
rect 23795 8396 23861 8397
rect 23795 8332 23796 8396
rect 23860 8332 23861 8396
rect 23795 8331 23861 8332
rect 23611 3500 23677 3501
rect 23611 3436 23612 3500
rect 23676 3436 23677 3500
rect 23611 3435 23677 3436
rect 23798 2005 23858 8331
rect 23979 8124 24045 8125
rect 23979 8060 23980 8124
rect 24044 8060 24045 8124
rect 23979 8059 24045 8060
rect 23982 4181 24042 8059
rect 24347 7716 24413 7717
rect 24347 7652 24348 7716
rect 24412 7652 24413 7716
rect 24347 7651 24413 7652
rect 24163 7580 24229 7581
rect 24163 7516 24164 7580
rect 24228 7516 24229 7580
rect 24163 7515 24229 7516
rect 23979 4180 24045 4181
rect 23979 4116 23980 4180
rect 24044 4116 24045 4180
rect 23979 4115 24045 4116
rect 23795 2004 23861 2005
rect 23795 1940 23796 2004
rect 23860 1940 23861 2004
rect 23795 1939 23861 1940
rect 24166 1869 24226 7515
rect 24350 4453 24410 7651
rect 24347 4452 24413 4453
rect 24347 4388 24348 4452
rect 24412 4388 24413 4452
rect 24347 4387 24413 4388
rect 24163 1868 24229 1869
rect 24163 1804 24164 1868
rect 24228 1804 24229 1868
rect 24163 1803 24229 1804
rect 24534 1325 24594 9691
rect 24718 1325 24778 9691
rect 25083 7852 25149 7853
rect 25083 7788 25084 7852
rect 25148 7788 25149 7852
rect 25083 7787 25149 7788
rect 24899 7580 24965 7581
rect 24899 7516 24900 7580
rect 24964 7516 24965 7580
rect 24899 7515 24965 7516
rect 24902 4589 24962 7515
rect 24899 4588 24965 4589
rect 24899 4524 24900 4588
rect 24964 4524 24965 4588
rect 24899 4523 24965 4524
rect 25086 4453 25146 7787
rect 24899 4452 24965 4453
rect 24899 4388 24900 4452
rect 24964 4388 24965 4452
rect 24899 4387 24965 4388
rect 25083 4452 25149 4453
rect 25083 4388 25084 4452
rect 25148 4388 25149 4452
rect 25083 4387 25149 4388
rect 24902 1869 24962 4387
rect 25300 2208 25620 9760
rect 25300 2144 25308 2208
rect 25372 2144 25388 2208
rect 25452 2144 25468 2208
rect 25532 2144 25548 2208
rect 25612 2144 25620 2208
rect 24899 1868 24965 1869
rect 24899 1804 24900 1868
rect 24964 1804 24965 1868
rect 24899 1803 24965 1804
rect 24531 1324 24597 1325
rect 24531 1260 24532 1324
rect 24596 1260 24597 1324
rect 24531 1259 24597 1260
rect 24715 1324 24781 1325
rect 24715 1260 24716 1324
rect 24780 1260 24781 1324
rect 24715 1259 24781 1260
rect 25300 1120 25620 2144
rect 25300 1056 25308 1120
rect 25372 1056 25388 1120
rect 25452 1056 25468 1120
rect 25532 1056 25548 1120
rect 25612 1056 25620 1120
rect 23427 1052 23493 1053
rect 23427 988 23428 1052
rect 23492 988 23493 1052
rect 23427 987 23493 988
rect 21587 780 21653 781
rect 21587 716 21588 780
rect 21652 716 21653 780
rect 21587 715 21653 716
rect 25300 496 25620 1056
rect 25940 11456 26260 11472
rect 25940 11392 25948 11456
rect 26012 11392 26028 11456
rect 26092 11392 26108 11456
rect 26172 11392 26188 11456
rect 26252 11392 26260 11456
rect 25940 10368 26260 11392
rect 25940 10304 25948 10368
rect 26012 10304 26028 10368
rect 26092 10304 26108 10368
rect 26172 10304 26188 10368
rect 26252 10304 26260 10368
rect 25940 1664 26260 10304
rect 26371 7580 26437 7581
rect 26371 7516 26372 7580
rect 26436 7516 26437 7580
rect 26371 7515 26437 7516
rect 26374 4453 26434 7515
rect 26580 5192 26900 11472
rect 26580 5128 26588 5192
rect 26652 5128 26668 5192
rect 26732 5128 26748 5192
rect 26812 5128 26828 5192
rect 26892 5128 26900 5192
rect 26580 5112 26900 5128
rect 26580 5048 26588 5112
rect 26652 5048 26668 5112
rect 26732 5048 26748 5112
rect 26812 5048 26828 5112
rect 26892 5048 26900 5112
rect 26580 5032 26900 5048
rect 26580 4968 26588 5032
rect 26652 4968 26668 5032
rect 26732 4968 26748 5032
rect 26812 4968 26828 5032
rect 26892 4968 26900 5032
rect 26580 4952 26900 4968
rect 26580 4888 26588 4952
rect 26652 4888 26668 4952
rect 26732 4888 26748 4952
rect 26812 4888 26828 4952
rect 26892 4888 26900 4952
rect 26371 4452 26437 4453
rect 26371 4388 26372 4452
rect 26436 4388 26437 4452
rect 26371 4387 26437 4388
rect 25940 1600 25948 1664
rect 26012 1600 26028 1664
rect 26092 1600 26108 1664
rect 26172 1600 26188 1664
rect 26252 1600 26260 1664
rect 25940 576 26260 1600
rect 25940 512 25948 576
rect 26012 512 26028 576
rect 26092 512 26108 576
rect 26172 512 26188 576
rect 26252 512 26260 576
rect 25940 496 26260 512
rect 26580 496 26900 4888
rect 27220 5832 27540 11472
rect 33300 10912 33620 11472
rect 33300 10848 33308 10912
rect 33372 10848 33388 10912
rect 33452 10848 33468 10912
rect 33532 10848 33548 10912
rect 33612 10848 33620 10912
rect 33300 9824 33620 10848
rect 33300 9760 33308 9824
rect 33372 9760 33388 9824
rect 33452 9760 33468 9824
rect 33532 9760 33548 9824
rect 33612 9760 33620 9824
rect 32995 9756 33061 9757
rect 32995 9692 32996 9756
rect 33060 9692 33061 9756
rect 32995 9691 33061 9692
rect 30787 8940 30853 8941
rect 30787 8876 30788 8940
rect 30852 8876 30853 8940
rect 30787 8875 30853 8876
rect 30419 8804 30485 8805
rect 30419 8740 30420 8804
rect 30484 8740 30485 8804
rect 30419 8739 30485 8740
rect 28395 8668 28461 8669
rect 28395 8604 28396 8668
rect 28460 8604 28461 8668
rect 28395 8603 28461 8604
rect 27843 8532 27909 8533
rect 27843 8468 27844 8532
rect 27908 8468 27909 8532
rect 27843 8467 27909 8468
rect 27659 8396 27725 8397
rect 27659 8332 27660 8396
rect 27724 8332 27725 8396
rect 27659 8331 27725 8332
rect 27220 5768 27228 5832
rect 27292 5768 27308 5832
rect 27372 5768 27388 5832
rect 27452 5768 27468 5832
rect 27532 5768 27540 5832
rect 27220 5752 27540 5768
rect 27220 5688 27228 5752
rect 27292 5688 27308 5752
rect 27372 5688 27388 5752
rect 27452 5688 27468 5752
rect 27532 5688 27540 5752
rect 27220 5672 27540 5688
rect 27220 5608 27228 5672
rect 27292 5608 27308 5672
rect 27372 5608 27388 5672
rect 27452 5608 27468 5672
rect 27532 5608 27540 5672
rect 27220 5592 27540 5608
rect 27220 5528 27228 5592
rect 27292 5528 27308 5592
rect 27372 5528 27388 5592
rect 27452 5528 27468 5592
rect 27532 5528 27540 5592
rect 27220 496 27540 5528
rect 27662 4045 27722 8331
rect 27846 4453 27906 8467
rect 28211 7852 28277 7853
rect 28211 7788 28212 7852
rect 28276 7788 28277 7852
rect 28211 7787 28277 7788
rect 28027 7104 28093 7105
rect 28027 7040 28028 7104
rect 28092 7040 28093 7104
rect 28027 7039 28093 7040
rect 27843 4452 27909 4453
rect 27843 4388 27844 4452
rect 27908 4388 27909 4452
rect 27843 4387 27909 4388
rect 27659 4044 27725 4045
rect 27659 3980 27660 4044
rect 27724 3980 27725 4044
rect 27659 3979 27725 3980
rect 28030 3909 28090 7039
rect 28027 3908 28093 3909
rect 28027 3844 28028 3908
rect 28092 3844 28093 3908
rect 28027 3843 28093 3844
rect 28214 2685 28274 7787
rect 28211 2684 28277 2685
rect 28211 2620 28212 2684
rect 28276 2620 28277 2684
rect 28211 2619 28277 2620
rect 28398 1325 28458 8603
rect 28947 8396 29013 8397
rect 28947 8332 28948 8396
rect 29012 8332 29013 8396
rect 28947 8331 29013 8332
rect 29131 8396 29197 8397
rect 29131 8332 29132 8396
rect 29196 8332 29197 8396
rect 29131 8331 29197 8332
rect 28579 7580 28645 7581
rect 28579 7516 28580 7580
rect 28644 7516 28645 7580
rect 28579 7515 28645 7516
rect 28582 4181 28642 7515
rect 28950 4181 29010 8331
rect 29134 4589 29194 8331
rect 30051 8260 30117 8261
rect 30051 8196 30052 8260
rect 30116 8196 30117 8260
rect 30051 8195 30117 8196
rect 29683 7172 29749 7173
rect 29683 7108 29684 7172
rect 29748 7108 29749 7172
rect 29683 7107 29749 7108
rect 29131 4588 29197 4589
rect 29131 4524 29132 4588
rect 29196 4524 29197 4588
rect 29131 4523 29197 4524
rect 28579 4180 28645 4181
rect 28579 4116 28580 4180
rect 28644 4116 28645 4180
rect 28579 4115 28645 4116
rect 28947 4180 29013 4181
rect 28947 4116 28948 4180
rect 29012 4116 29013 4180
rect 28947 4115 29013 4116
rect 29686 2549 29746 7107
rect 30054 4045 30114 8195
rect 30235 7104 30301 7105
rect 30235 7040 30236 7104
rect 30300 7040 30301 7104
rect 30235 7039 30301 7040
rect 30051 4044 30117 4045
rect 30051 3980 30052 4044
rect 30116 3980 30117 4044
rect 30051 3979 30117 3980
rect 30238 3229 30298 7039
rect 30235 3228 30301 3229
rect 30235 3164 30236 3228
rect 30300 3164 30301 3228
rect 30235 3163 30301 3164
rect 29683 2548 29749 2549
rect 29683 2484 29684 2548
rect 29748 2484 29749 2548
rect 29683 2483 29749 2484
rect 30422 1325 30482 8739
rect 30603 7852 30669 7853
rect 30603 7788 30604 7852
rect 30668 7788 30669 7852
rect 30603 7787 30669 7788
rect 30606 1325 30666 7787
rect 28395 1324 28461 1325
rect 28395 1260 28396 1324
rect 28460 1260 28461 1324
rect 28395 1259 28461 1260
rect 30419 1324 30485 1325
rect 30419 1260 30420 1324
rect 30484 1260 30485 1324
rect 30419 1259 30485 1260
rect 30603 1324 30669 1325
rect 30603 1260 30604 1324
rect 30668 1260 30669 1324
rect 30603 1259 30669 1260
rect 30790 1189 30850 8875
rect 30971 8532 31037 8533
rect 30971 8468 30972 8532
rect 31036 8468 31037 8532
rect 30971 8467 31037 8468
rect 30974 1325 31034 8467
rect 31891 7580 31957 7581
rect 31891 7516 31892 7580
rect 31956 7516 31957 7580
rect 31891 7515 31957 7516
rect 31155 7444 31221 7445
rect 31155 7380 31156 7444
rect 31220 7380 31221 7444
rect 31155 7379 31221 7380
rect 31158 2005 31218 7379
rect 31155 2004 31221 2005
rect 31155 1940 31156 2004
rect 31220 1940 31221 2004
rect 31155 1939 31221 1940
rect 31894 1733 31954 7515
rect 32627 6356 32693 6357
rect 32627 6292 32628 6356
rect 32692 6292 32693 6356
rect 32627 6291 32693 6292
rect 32630 3773 32690 6291
rect 32627 3772 32693 3773
rect 32627 3708 32628 3772
rect 32692 3708 32693 3772
rect 32627 3707 32693 3708
rect 31891 1732 31957 1733
rect 31891 1668 31892 1732
rect 31956 1668 31957 1732
rect 31891 1667 31957 1668
rect 32998 1325 33058 9691
rect 33300 2208 33620 9760
rect 33300 2144 33308 2208
rect 33372 2144 33388 2208
rect 33452 2144 33468 2208
rect 33532 2144 33548 2208
rect 33612 2144 33620 2208
rect 30971 1324 31037 1325
rect 30971 1260 30972 1324
rect 31036 1260 31037 1324
rect 30971 1259 31037 1260
rect 32995 1324 33061 1325
rect 32995 1260 32996 1324
rect 33060 1260 33061 1324
rect 32995 1259 33061 1260
rect 30787 1188 30853 1189
rect 30787 1124 30788 1188
rect 30852 1124 30853 1188
rect 30787 1123 30853 1124
rect 33300 1120 33620 2144
rect 33300 1056 33308 1120
rect 33372 1056 33388 1120
rect 33452 1056 33468 1120
rect 33532 1056 33548 1120
rect 33612 1056 33620 1120
rect 33300 496 33620 1056
rect 33940 11456 34260 11472
rect 33940 11392 33948 11456
rect 34012 11392 34028 11456
rect 34092 11392 34108 11456
rect 34172 11392 34188 11456
rect 34252 11392 34260 11456
rect 33940 10368 34260 11392
rect 33940 10304 33948 10368
rect 34012 10304 34028 10368
rect 34092 10304 34108 10368
rect 34172 10304 34188 10368
rect 34252 10304 34260 10368
rect 33940 9280 34260 10304
rect 33940 9216 33948 9280
rect 34012 9216 34028 9280
rect 34092 9216 34108 9280
rect 34172 9216 34188 9280
rect 34252 9216 34260 9280
rect 33940 8192 34260 9216
rect 33940 8128 33948 8192
rect 34012 8128 34028 8192
rect 34092 8128 34108 8192
rect 34172 8128 34188 8192
rect 34252 8128 34260 8192
rect 33940 7104 34260 8128
rect 33940 7040 33948 7104
rect 34012 7040 34028 7104
rect 34092 7040 34108 7104
rect 34172 7040 34188 7104
rect 34252 7040 34260 7104
rect 33940 6016 34260 7040
rect 33940 5952 33948 6016
rect 34012 5952 34028 6016
rect 34092 5952 34108 6016
rect 34172 5952 34188 6016
rect 34252 5952 34260 6016
rect 33940 4928 34260 5952
rect 33940 4864 33948 4928
rect 34012 4864 34028 4928
rect 34092 4864 34108 4928
rect 34172 4864 34188 4928
rect 34252 4864 34260 4928
rect 33940 3840 34260 4864
rect 33940 3776 33948 3840
rect 34012 3776 34028 3840
rect 34092 3776 34108 3840
rect 34172 3776 34188 3840
rect 34252 3776 34260 3840
rect 33940 2752 34260 3776
rect 41300 10912 41620 11472
rect 41300 10848 41308 10912
rect 41372 10848 41388 10912
rect 41452 10848 41468 10912
rect 41532 10848 41548 10912
rect 41612 10848 41620 10912
rect 41300 9824 41620 10848
rect 41300 9760 41308 9824
rect 41372 9760 41388 9824
rect 41452 9760 41468 9824
rect 41532 9760 41548 9824
rect 41612 9760 41620 9824
rect 41300 8736 41620 9760
rect 41300 8672 41308 8736
rect 41372 8672 41388 8736
rect 41452 8672 41468 8736
rect 41532 8672 41548 8736
rect 41612 8672 41620 8736
rect 41300 7648 41620 8672
rect 41300 7584 41308 7648
rect 41372 7584 41388 7648
rect 41452 7584 41468 7648
rect 41532 7584 41548 7648
rect 41612 7584 41620 7648
rect 41300 6560 41620 7584
rect 41300 6496 41308 6560
rect 41372 6496 41388 6560
rect 41452 6496 41468 6560
rect 41532 6496 41548 6560
rect 41612 6496 41620 6560
rect 41300 5472 41620 6496
rect 41300 5408 41308 5472
rect 41372 5408 41388 5472
rect 41452 5408 41468 5472
rect 41532 5408 41548 5472
rect 41612 5408 41620 5472
rect 41300 4384 41620 5408
rect 41300 4320 41308 4384
rect 41372 4320 41388 4384
rect 41452 4320 41468 4384
rect 41532 4320 41548 4384
rect 41612 4320 41620 4384
rect 41300 3296 41620 4320
rect 41300 3232 41308 3296
rect 41372 3232 41388 3296
rect 41452 3232 41468 3296
rect 41532 3232 41548 3296
rect 41612 3232 41620 3296
rect 38883 3228 38949 3229
rect 38883 3164 38884 3228
rect 38948 3164 38949 3228
rect 38883 3163 38949 3164
rect 33940 2688 33948 2752
rect 34012 2688 34028 2752
rect 34092 2688 34108 2752
rect 34172 2688 34188 2752
rect 34252 2688 34260 2752
rect 33940 1664 34260 2688
rect 38699 2548 38765 2549
rect 38699 2484 38700 2548
rect 38764 2484 38765 2548
rect 38699 2483 38765 2484
rect 38702 1869 38762 2483
rect 38886 1869 38946 3163
rect 41300 2208 41620 3232
rect 41300 2144 41308 2208
rect 41372 2144 41388 2208
rect 41452 2144 41468 2208
rect 41532 2144 41548 2208
rect 41612 2144 41620 2208
rect 38699 1868 38765 1869
rect 38699 1804 38700 1868
rect 38764 1804 38765 1868
rect 38699 1803 38765 1804
rect 38883 1868 38949 1869
rect 38883 1804 38884 1868
rect 38948 1804 38949 1868
rect 38883 1803 38949 1804
rect 33940 1600 33948 1664
rect 34012 1600 34028 1664
rect 34092 1600 34108 1664
rect 34172 1600 34188 1664
rect 34252 1600 34260 1664
rect 33940 576 34260 1600
rect 33940 512 33948 576
rect 34012 512 34028 576
rect 34092 512 34108 576
rect 34172 512 34188 576
rect 34252 512 34260 576
rect 33940 496 34260 512
rect 41300 1120 41620 2144
rect 41300 1056 41308 1120
rect 41372 1056 41388 1120
rect 41452 1056 41468 1120
rect 41532 1056 41548 1120
rect 41612 1056 41620 1120
rect 41300 496 41620 1056
rect 41940 11456 42260 11472
rect 41940 11392 41948 11456
rect 42012 11392 42028 11456
rect 42092 11392 42108 11456
rect 42172 11392 42188 11456
rect 42252 11392 42260 11456
rect 41940 10368 42260 11392
rect 41940 10304 41948 10368
rect 42012 10304 42028 10368
rect 42092 10304 42108 10368
rect 42172 10304 42188 10368
rect 42252 10304 42260 10368
rect 41940 9280 42260 10304
rect 41940 9216 41948 9280
rect 42012 9216 42028 9280
rect 42092 9216 42108 9280
rect 42172 9216 42188 9280
rect 42252 9216 42260 9280
rect 41940 8192 42260 9216
rect 41940 8128 41948 8192
rect 42012 8128 42028 8192
rect 42092 8128 42108 8192
rect 42172 8128 42188 8192
rect 42252 8128 42260 8192
rect 41940 7104 42260 8128
rect 41940 7040 41948 7104
rect 42012 7040 42028 7104
rect 42092 7040 42108 7104
rect 42172 7040 42188 7104
rect 42252 7040 42260 7104
rect 41940 6016 42260 7040
rect 41940 5952 41948 6016
rect 42012 5952 42028 6016
rect 42092 5952 42108 6016
rect 42172 5952 42188 6016
rect 42252 5952 42260 6016
rect 41940 4928 42260 5952
rect 41940 4864 41948 4928
rect 42012 4864 42028 4928
rect 42092 4864 42108 4928
rect 42172 4864 42188 4928
rect 42252 4864 42260 4928
rect 41940 3840 42260 4864
rect 41940 3776 41948 3840
rect 42012 3776 42028 3840
rect 42092 3776 42108 3840
rect 42172 3776 42188 3840
rect 42252 3776 42260 3840
rect 41940 2752 42260 3776
rect 41940 2688 41948 2752
rect 42012 2688 42028 2752
rect 42092 2688 42108 2752
rect 42172 2688 42188 2752
rect 42252 2688 42260 2752
rect 41940 1664 42260 2688
rect 41940 1600 41948 1664
rect 42012 1600 42028 1664
rect 42092 1600 42108 1664
rect 42172 1600 42188 1664
rect 42252 1600 42260 1664
rect 41940 576 42260 1600
rect 41940 512 41948 576
rect 42012 512 42028 576
rect 42092 512 42108 576
rect 42172 512 42188 576
rect 42252 512 42260 576
rect 41940 496 42260 512
use sky130_fd_sc_hd__inv_2  _000_
timestamp 21601
transform 1 0 35604 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _001_
timestamp 21601
transform 1 0 35972 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _002_
timestamp 21601
transform 1 0 35880 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _003_
timestamp 21601
transform 1 0 36156 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _004_
timestamp 21601
transform 1 0 39836 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _005_
timestamp 21601
transform 1 0 40112 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _006_
timestamp 21601
transform 1 0 40388 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _007_
timestamp 21601
transform 1 0 40664 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _008_
timestamp 21601
transform 1 0 38640 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _009_
timestamp 21601
transform 1 0 39192 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _010_
timestamp 21601
transform 1 0 39468 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _011_
timestamp 21601
transform 1 0 39744 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _012_
timestamp 21601
transform 1 0 40940 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _013_
timestamp 21601
transform 1 0 41216 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _014_
timestamp 21601
transform 1 0 40020 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _015_
timestamp 21601
transform 1 0 40756 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _016_
timestamp 21601
transform -1 0 23644 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _017_
timestamp 21601
transform -1 0 23368 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _018_
timestamp 21601
transform 1 0 25208 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _019_
timestamp 21601
transform 1 0 25484 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _020_
timestamp 21601
transform -1 0 25300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _021_
timestamp 21601
transform 1 0 25760 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _022_
timestamp 21601
transform -1 0 25760 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _023_
timestamp 21601
transform -1 0 26128 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _024_
timestamp 21601
transform 1 0 27784 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _025_
timestamp 21601
transform 1 0 28060 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _026_
timestamp 21601
transform 1 0 28336 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _027_
timestamp 21601
transform 1 0 28244 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _028_
timestamp 21601
transform 1 0 28520 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _029_
timestamp 21601
transform 1 0 30360 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _030_
timestamp 21601
transform 1 0 30636 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _031_
timestamp 21601
transform 1 0 30912 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _032_
timestamp 21601
transform -1 0 28520 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _033_
timestamp 21601
transform -1 0 28796 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _034_
timestamp 21601
transform 1 0 32936 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _035_
timestamp 21601
transform 1 0 30728 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _036_
timestamp 21601
transform 1 0 31004 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _037_
timestamp 21601
transform 1 0 30360 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _038_
timestamp 21601
transform 1 0 30636 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _039_
timestamp 21601
transform 1 0 30912 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _040_
timestamp 21601
transform 1 0 32936 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _041_
timestamp 21601
transform 1 0 33212 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _042_
timestamp 21601
transform 1 0 33488 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _043_
timestamp 21601
transform 1 0 32752 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _044_
timestamp 21601
transform 1 0 33028 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _045_
timestamp 21601
transform 1 0 34224 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _046_
timestamp 21601
transform 1 0 32752 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _047_
timestamp 21601
transform 1 0 34500 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _048_
timestamp 21601
transform 1 0 34040 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _049_
timestamp 21601
transform 1 0 35880 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _050_
timestamp 21601
transform 1 0 35512 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _051_
timestamp 21601
transform 1 0 35604 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _052_
timestamp 21601
transform 1 0 36248 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _053_
timestamp 21601
transform 1 0 37444 0 1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _054_
timestamp 21601
transform 1 0 36892 0 -1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _055_
timestamp 21601
transform 1 0 38272 0 -1 2720
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _056_
timestamp 21601
transform 1 0 39192 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _057_
timestamp 21601
transform 1 0 32752 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _058_
timestamp 21601
transform 1 0 3680 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _059_
timestamp 21601
transform -1 0 5336 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _060_
timestamp 21601
transform 1 0 4876 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _061_
timestamp 21601
transform -1 0 4968 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _062_
timestamp 21601
transform 1 0 4968 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _063_
timestamp 21601
transform 1 0 5704 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _064_
timestamp 21601
transform -1 0 6256 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _065_
timestamp 21601
transform 1 0 6256 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _066_
timestamp 21601
transform 1 0 6256 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _067_
timestamp 21601
transform 1 0 6808 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _068_
timestamp 21601
transform 1 0 7084 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _069_
timestamp 21601
transform 1 0 6900 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _070_
timestamp 21601
transform 1 0 7636 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _071_
timestamp 21601
transform 1 0 7544 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _072_
timestamp 21601
transform -1 0 8832 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _073_
timestamp 21601
transform 1 0 8464 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _074_
timestamp 21601
transform -1 0 9292 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _075_
timestamp 21601
transform 1 0 8924 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _076_
timestamp 21601
transform 1 0 8832 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _077_
timestamp 21601
transform -1 0 9936 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _078_
timestamp 21601
transform 1 0 9292 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _079_
timestamp 21601
transform 1 0 9752 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _080_
timestamp 21601
transform 1 0 9936 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _081_
timestamp 21601
transform 1 0 9476 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _082_
timestamp 21601
transform 1 0 10120 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _083_
timestamp 21601
transform -1 0 10764 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _084_
timestamp 21601
transform 1 0 10856 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _085_
timestamp 21601
transform 1 0 10120 0 -1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _086_
timestamp 21601
transform 1 0 11040 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _087_
timestamp 21601
transform 1 0 10672 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _088_
timestamp 21601
transform -1 0 11316 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _089_
timestamp 21601
transform 1 0 12420 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _090_
timestamp 21601
transform -1 0 12696 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _091_
timestamp 21601
transform -1 0 13892 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _092_
timestamp 21601
transform 1 0 12696 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _093_
timestamp 21601
transform 1 0 13984 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _094_
timestamp 21601
transform 1 0 13892 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _095_
timestamp 21601
transform -1 0 14628 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _096_
timestamp 21601
transform 1 0 14536 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _097_
timestamp 21601
transform -1 0 15824 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _098_
timestamp 21601
transform 1 0 15272 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _099_
timestamp 21601
transform -1 0 16652 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _100_
timestamp 21601
transform 1 0 16008 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _101_
timestamp 21601
transform 1 0 14628 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _102_
timestamp 21601
transform -1 0 17296 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _103_
timestamp 21601
transform -1 0 17204 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _104_
timestamp 21601
transform -1 0 17756 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _105_
timestamp 21601
transform 1 0 17480 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _106_
timestamp 21601
transform -1 0 18400 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _107_
timestamp 21601
transform 1 0 17204 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _108_
timestamp 21601
transform 1 0 17848 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _109_
timestamp 21601
transform 1 0 18676 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _110_
timestamp 21601
transform -1 0 19136 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _111_
timestamp 21601
transform 1 0 19320 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _112_
timestamp 21601
transform 1 0 19504 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _113_
timestamp 21601
transform -1 0 20608 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _114_
timestamp 21601
transform 1 0 19136 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _115_
timestamp 21601
transform 1 0 19780 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _116_
timestamp 21601
transform 1 0 20608 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _117_
timestamp 21601
transform 1 0 20424 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _118_
timestamp 21601
transform 1 0 21252 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _119_
timestamp 21601
transform -1 0 21896 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _120_
timestamp 21601
transform -1 0 22540 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _121_
timestamp 21601
transform 1 0 21896 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _122_
timestamp 21601
transform -1 0 23184 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _123_
timestamp 21601
transform 1 0 22632 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _124_
timestamp 21601
transform -1 0 25024 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _125_
timestamp 21601
transform -1 0 23920 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _126_
timestamp 21601
transform -1 0 24380 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _127_
timestamp 21601
transform -1 0 24564 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _128_
timestamp 21601
transform -1 0 25668 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _129_
timestamp 21601
transform -1 0 25484 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _130_
timestamp 21601
transform -1 0 26128 0 -1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _131_
timestamp 21601
transform -1 0 26956 0 1 8160
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _132_
timestamp 21601
transform 1 0 32844 0 -1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _133_
timestamp 21601
transform 1 0 33028 0 1 5984
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _134_
timestamp 21601
transform 1 0 33120 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _135_
timestamp 21601
transform 1 0 33396 0 1 3808
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _136_
timestamp 21601
transform 1 0 33304 0 1 544
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _137_
timestamp 21601
transform 1 0 33304 0 1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _138_
timestamp 21601
transform 1 0 35880 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _139_
timestamp 21601
transform 1 0 30728 0 -1 1632
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__000__Y
timestamp 21601
transform -1 0 36064 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__001__Y
timestamp 21601
transform -1 0 36432 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__002__Y
timestamp 21601
transform -1 0 36524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__003__Y
timestamp 21601
transform -1 0 37076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__004__Y
timestamp 21601
transform -1 0 42320 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__005__Y
timestamp 21601
transform -1 0 41400 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__006__Y
timestamp 21601
transform -1 0 42504 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__007__Y
timestamp 21601
transform -1 0 42688 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__008__Y
timestamp 21601
transform -1 0 40848 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__009__Y
timestamp 21601
transform -1 0 40204 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__010__Y
timestamp 21601
transform -1 0 40388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__011__Y
timestamp 21601
transform -1 0 41032 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__012__Y
timestamp 21601
transform -1 0 42136 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__013__Y
timestamp 21601
transform -1 0 42320 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__014__Y
timestamp 21601
transform -1 0 41216 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__015__Y
timestamp 21601
transform -1 0 41952 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__049__B
timestamp 21601
transform -1 0 38456 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__050__B
timestamp 21601
transform -1 0 35696 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__051__B
timestamp 21601
transform -1 0 35604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__052__B
timestamp 21601
transform -1 0 36708 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__053__B
timestamp 21601
transform -1 0 37904 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__054__B
timestamp 21601
transform -1 0 36892 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__055__B
timestamp 21601
transform -1 0 39008 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__056__B
timestamp 21601
transform -1 0 42136 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__057__B
timestamp 21601
transform -1 0 33580 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__B
timestamp 21601
transform -1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__058__X
timestamp 21601
transform 1 0 4324 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__B
timestamp 21601
transform 1 0 4140 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__059__X
timestamp 21601
transform -1 0 4692 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__B
timestamp 21601
transform 1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__060__X
timestamp 21601
transform -1 0 5704 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__B
timestamp 21601
transform 1 0 4140 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__X
timestamp 21601
transform -1 0 4692 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__B
timestamp 21601
transform 1 0 4324 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__062__X
timestamp 21601
transform 1 0 5428 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__B
timestamp 21601
transform -1 0 5888 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__X
timestamp 21601
transform 1 0 6348 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__B
timestamp 21601
transform -1 0 5612 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__064__X
timestamp 21601
transform -1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__B
timestamp 21601
transform 1 0 6072 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__X
timestamp 21601
transform -1 0 7084 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__B
timestamp 21601
transform 1 0 5704 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__066__X
timestamp 21601
transform -1 0 6808 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B
timestamp 21601
transform -1 0 6808 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__X
timestamp 21601
transform 1 0 7452 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__B
timestamp 21601
transform 1 0 6900 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__068__X
timestamp 21601
transform -1 0 7912 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__B
timestamp 21601
transform -1 0 6624 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__X
timestamp 21601
transform 1 0 7452 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__B
timestamp 21601
transform -1 0 7820 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__070__X
timestamp 21601
transform 1 0 8280 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__B
timestamp 21601
transform 1 0 7360 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__X
timestamp 21601
transform -1 0 8464 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__B
timestamp 21601
transform 1 0 7820 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__072__X
timestamp 21601
transform -1 0 8188 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__B
timestamp 21601
transform -1 0 8648 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__X
timestamp 21601
transform 1 0 9108 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__B
timestamp 21601
transform -1 0 8464 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__X
timestamp 21601
transform -1 0 8648 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__B
timestamp 21601
transform -1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__075__X
timestamp 21601
transform -1 0 9844 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__B
timestamp 21601
transform 1 0 8648 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__X
timestamp 21601
transform -1 0 9660 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__B
timestamp 21601
transform -1 0 9476 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__077__X
timestamp 21601
transform -1 0 9292 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__B
timestamp 21601
transform -1 0 8464 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__X
timestamp 21601
transform 1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__B
timestamp 21601
transform -1 0 10028 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__079__X
timestamp 21601
transform -1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__B
timestamp 21601
transform -1 0 9936 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__X
timestamp 21601
transform 1 0 10856 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__B
timestamp 21601
transform 1 0 9292 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__081__X
timestamp 21601
transform -1 0 10304 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__B
timestamp 21601
transform 1 0 9568 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__X
timestamp 21601
transform -1 0 11040 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__B
timestamp 21601
transform -1 0 9752 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__083__X
timestamp 21601
transform -1 0 10580 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__B
timestamp 21601
transform 1 0 10212 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__X
timestamp 21601
transform -1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__B
timestamp 21601
transform -1 0 10120 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__085__X
timestamp 21601
transform 1 0 10856 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__B
timestamp 21601
transform -1 0 10764 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__X
timestamp 21601
transform 1 0 11684 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__B
timestamp 21601
transform -1 0 10672 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__087__X
timestamp 21601
transform -1 0 11316 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__B
timestamp 21601
transform -1 0 11316 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__X
timestamp 21601
transform -1 0 11316 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__B
timestamp 21601
transform 1 0 12052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__089__X
timestamp 21601
transform 1 0 13064 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__B
timestamp 21601
transform -1 0 12052 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__X
timestamp 21601
transform -1 0 12052 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__B
timestamp 21601
transform 1 0 12236 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__091__X
timestamp 21601
transform -1 0 13248 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__B
timestamp 21601
transform -1 0 11868 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__X
timestamp 21601
transform 1 0 13432 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__B
timestamp 21601
transform -1 0 13984 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__093__X
timestamp 21601
transform -1 0 14904 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__B
timestamp 21601
transform -1 0 13892 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__X
timestamp 21601
transform 1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__B
timestamp 21601
transform -1 0 13616 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__X
timestamp 21601
transform -1 0 13800 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__B
timestamp 21601
transform -1 0 14536 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__096__X
timestamp 21601
transform -1 0 15088 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__B
timestamp 21601
transform -1 0 14904 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__X
timestamp 21601
transform -1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B
timestamp 21601
transform -1 0 15272 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__X
timestamp 21601
transform 1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__B
timestamp 21601
transform -1 0 15824 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__X
timestamp 21601
transform -1 0 16192 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__B
timestamp 21601
transform -1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__X
timestamp 21601
transform -1 0 16836 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__B
timestamp 21601
transform -1 0 13984 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__X
timestamp 21601
transform 1 0 15456 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__B
timestamp 21601
transform -1 0 17020 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__X
timestamp 21601
transform -1 0 17480 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__B
timestamp 21601
transform -1 0 16560 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__X
timestamp 21601
transform -1 0 16376 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__B
timestamp 21601
transform -1 0 16560 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__104__X
timestamp 21601
transform -1 0 16928 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__B
timestamp 21601
transform -1 0 17664 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__X
timestamp 21601
transform -1 0 18308 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__B
timestamp 21601
transform -1 0 17480 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__X
timestamp 21601
transform -1 0 17112 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__B
timestamp 21601
transform -1 0 17204 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__X
timestamp 21601
transform 1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__B
timestamp 21601
transform -1 0 17848 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__108__X
timestamp 21601
transform 1 0 18308 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__B
timestamp 21601
transform -1 0 18768 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__X
timestamp 21601
transform -1 0 19320 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__B
timestamp 21601
transform -1 0 18308 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__X
timestamp 21601
transform -1 0 18952 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__B
timestamp 21601
transform -1 0 19136 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__X
timestamp 21601
transform -1 0 20332 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__B
timestamp 21601
transform -1 0 19504 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__112__X
timestamp 21601
transform -1 0 20976 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__B
timestamp 21601
transform -1 0 19504 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__X
timestamp 21601
transform -1 0 21620 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__B
timestamp 21601
transform -1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__X
timestamp 21601
transform 1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__B
timestamp 21601
transform -1 0 19780 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__X
timestamp 21601
transform 1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__B
timestamp 21601
transform -1 0 20792 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__X
timestamp 21601
transform -1 0 22264 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__B
timestamp 21601
transform -1 0 20424 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__X
timestamp 21601
transform 1 0 21160 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__B
timestamp 21601
transform -1 0 20608 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__X
timestamp 21601
transform -1 0 22080 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__B
timestamp 21601
transform -1 0 21436 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__X
timestamp 21601
transform -1 0 21068 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__B
timestamp 21601
transform -1 0 21896 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__X
timestamp 21601
transform -1 0 22816 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__B
timestamp 21601
transform -1 0 20884 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__X
timestamp 21601
transform -1 0 23368 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__B
timestamp 21601
transform -1 0 23552 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__X
timestamp 21601
transform -1 0 23368 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__B
timestamp 21601
transform -1 0 22632 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__X
timestamp 21601
transform -1 0 24104 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__B
timestamp 21601
transform -1 0 24748 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__X
timestamp 21601
transform -1 0 26220 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__B
timestamp 21601
transform -1 0 23552 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__X
timestamp 21601
transform -1 0 24472 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__B
timestamp 21601
transform -1 0 23920 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__X
timestamp 21601
transform -1 0 25852 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__B
timestamp 21601
transform -1 0 24288 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__X
timestamp 21601
transform -1 0 24748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__B
timestamp 21601
transform -1 0 26036 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__X
timestamp 21601
transform -1 0 26496 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__B
timestamp 21601
transform -1 0 24932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__X
timestamp 21601
transform -1 0 25668 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__B
timestamp 21601
transform -1 0 25484 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__X
timestamp 21601
transform -1 0 26680 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__B
timestamp 21601
transform -1 0 27140 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__X
timestamp 21601
transform -1 0 27324 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__B
timestamp 21601
transform -1 0 33672 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__B
timestamp 21601
transform -1 0 33028 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__B
timestamp 21601
transform -1 0 33948 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__B
timestamp 21601
transform -1 0 35052 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__B
timestamp 21601
transform -1 0 34132 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__B
timestamp 21601
transform -1 0 35788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__B
timestamp 21601
transform -1 0 39468 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__B
timestamp 21601
transform -1 0 33120 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_hreadyout_ack_gate_A
timestamp 21601
transform -1 0 34224 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[0\]_A
timestamp 21601
transform -1 0 34960 0 -1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[1\]_A
timestamp 21601
transform -1 0 35328 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[2\]_A
timestamp 21601
transform -1 0 35512 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[3\]_A
timestamp 21601
transform -1 0 36340 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[4\]_A
timestamp 21601
transform -1 0 41952 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[5\]_A
timestamp 21601
transform 1 0 37076 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[6\]_A
timestamp 21601
transform -1 0 40020 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[7\]_A
timestamp 21601
transform -1 0 39652 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[8\]_A
timestamp 21601
transform -1 0 38824 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[9\]_A
timestamp 21601
transform -1 0 38088 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[10\]_A
timestamp 21601
transform -1 0 38272 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[11\]_A
timestamp 21601
transform -1 0 40480 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[12\]_A
timestamp 21601
transform -1 0 40664 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[13\]_A
timestamp 21601
transform -1 0 41584 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[14\]_A
timestamp 21601
transform -1 0 41400 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_irq_gates\[15\]_A
timestamp 21601
transform 1 0 40388 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output1_X
timestamp 21601
transform -1 0 23092 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output2_X
timestamp 21601
transform -1 0 23552 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output3_X
timestamp 21601
transform -1 0 27968 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output4_X
timestamp 21601
transform -1 0 36524 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output5_X
timestamp 21601
transform -1 0 31372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output6_X
timestamp 21601
transform -1 0 32936 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output7_X
timestamp 21601
transform -1 0 39100 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output8_X
timestamp 21601
transform -1 0 34500 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output9_X
timestamp 21601
transform -1 0 34684 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output10_X
timestamp 21601
transform -1 0 33948 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output11_X
timestamp 21601
transform -1 0 33488 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output12_X
timestamp 21601
transform -1 0 26220 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output13_X
timestamp 21601
transform -1 0 34132 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output14_X
timestamp 21601
transform -1 0 33304 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output15_X
timestamp 21601
transform -1 0 39100 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output16_X
timestamp 21601
transform -1 0 41676 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output17_X
timestamp 21601
transform -1 0 34868 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output18_X
timestamp 21601
transform -1 0 38640 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output19_X
timestamp 21601
transform -1 0 35328 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output20_X
timestamp 21601
transform -1 0 39284 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output21_X
timestamp 21601
transform -1 0 34408 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output22_X
timestamp 21601
transform -1 0 41216 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output23_X
timestamp 21601
transform -1 0 25484 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output24_X
timestamp 21601
transform -1 0 39100 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output25_X
timestamp 21601
transform -1 0 38272 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output26_X
timestamp 21601
transform -1 0 26220 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output27_X
timestamp 21601
transform -1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output28_X
timestamp 21601
transform -1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output29_X
timestamp 21601
transform -1 0 31372 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output30_X
timestamp 21601
transform -1 0 28796 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output31_X
timestamp 21601
transform -1 0 28152 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output32_X
timestamp 21601
transform -1 0 26036 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output33_X
timestamp 21601
transform -1 0 39836 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[0\]_A
timestamp 21601
transform -1 0 24564 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[1\]_A
timestamp 21601
transform 1 0 24564 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[2\]_A
timestamp 21601
transform -1 0 25024 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[3\]_A
timestamp 21601
transform 1 0 25300 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[4\]_A
timestamp 21601
transform 1 0 25484 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[5\]_A
timestamp 21601
transform -1 0 26772 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[6\]_A
timestamp 21601
transform -1 0 26956 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[7\]_A
timestamp 21601
transform -1 0 27140 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[8\]_A
timestamp 21601
transform -1 0 27140 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[9\]_A
timestamp 21601
transform -1 0 27876 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[10\]_A
timestamp 21601
transform -1 0 28060 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[11\]_A
timestamp 21601
transform -1 0 28244 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[12\]_A
timestamp 21601
transform 1 0 27784 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[13\]_A
timestamp 21601
transform -1 0 28520 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[14\]_A
timestamp 21601
transform -1 0 29072 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[15\]_A
timestamp 21601
transform 1 0 28428 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[16\]_A
timestamp 21601
transform -1 0 29256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[17\]_A
timestamp 21601
transform -1 0 29624 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[18\]_A
timestamp 21601
transform -1 0 29808 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[19\]_A
timestamp 21601
transform -1 0 30176 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[20\]_A
timestamp 21601
transform -1 0 30360 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[21\]_A
timestamp 21601
transform -1 0 30360 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[22\]_A
timestamp 21601
transform -1 0 31096 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[23\]_A
timestamp 21601
transform -1 0 31280 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[24\]_A
timestamp 21601
transform -1 0 31372 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[25\]_A
timestamp 21601
transform -1 0 31648 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[26\]_A
timestamp 21601
transform -1 0 31924 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[27\]_A
timestamp 21601
transform -1 0 32108 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[28\]_A
timestamp 21601
transform 1 0 32200 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[29\]_A
timestamp 21601
transform -1 0 33580 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[30\]_A
timestamp 21601
transform -1 0 33764 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_wb_hrdata_gates\[31\]_A
timestamp 21601
transform -1 0 33948 0 -1 11424
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3
timestamp 1636990056
transform 1 0 736 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15
timestamp 1636990056
transform 1 0 1840 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27
timestamp 21601
transform 1 0 2944 0 1 544
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1636990056
transform 1 0 3128 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1636990056
transform 1 0 4232 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 21601
transform 1 0 5336 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1636990056
transform 1 0 5704 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1636990056
transform 1 0 6808 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 21601
transform 1 0 7912 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1636990056
transform 1 0 8280 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1636990056
transform 1 0 9384 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 21601
transform 1 0 10488 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1636990056
transform 1 0 10856 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1636990056
transform 1 0 11960 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 21601
transform 1 0 13064 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1636990056
transform 1 0 13432 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1636990056
transform 1 0 14536 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 21601
transform 1 0 15640 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_169
timestamp 1636990056
transform 1 0 16008 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_181
timestamp 1636990056
transform 1 0 17112 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 21601
transform 1 0 18216 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1636990056
transform 1 0 18584 0 1 544
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1636990056
transform 1 0 19688 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 21601
transform 1 0 20792 0 1 544
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1636990056
transform 1 0 21160 0 1 544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_237
timestamp 21601
transform 1 0 22264 0 1 544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_243
timestamp 21601
transform 1 0 22816 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_356
timestamp 21601
transform 1 0 33212 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_459
timestamp 21601
transform 1 0 42688 0 1 544
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3
timestamp 1636990056
transform 1 0 736 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_15
timestamp 1636990056
transform 1 0 1840 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_27
timestamp 1636990056
transform 1 0 2944 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_39
timestamp 1636990056
transform 1 0 4048 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_51
timestamp 21601
transform 1 0 5152 0 -1 1632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 21601
transform 1 0 5520 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1636990056
transform 1 0 5704 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1636990056
transform 1 0 6808 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1636990056
transform 1 0 7912 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1636990056
transform 1 0 9016 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 21601
transform 1 0 10120 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 21601
transform 1 0 10672 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1636990056
transform 1 0 10856 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1636990056
transform 1 0 11960 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1636990056
transform 1 0 13064 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1636990056
transform 1 0 14168 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 21601
transform 1 0 15272 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 21601
transform 1 0 15824 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1636990056
transform 1 0 16008 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1636990056
transform 1 0 17112 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1636990056
transform 1 0 18216 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1636990056
transform 1 0 19320 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 21601
transform 1 0 20424 0 -1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 21601
transform 1 0 20976 0 -1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1636990056
transform 1 0 21160 0 -1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1636990056
transform 1 0 22264 0 -1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_275
timestamp 21601
transform 1 0 25760 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 21601
transform 1 0 26128 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_447
timestamp 21601
transform 1 0 41584 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_455
timestamp 21601
transform 1 0 42320 0 -1 1632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_463
timestamp 21601
transform 1 0 43056 0 -1 1632
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1636990056
transform 1 0 736 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1636990056
transform 1 0 1840 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 21601
transform 1 0 2944 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1636990056
transform 1 0 3128 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1636990056
transform 1 0 4232 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1636990056
transform 1 0 5336 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1636990056
transform 1 0 6440 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 21601
transform 1 0 7544 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 21601
transform 1 0 8096 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1636990056
transform 1 0 8280 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1636990056
transform 1 0 9384 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1636990056
transform 1 0 10488 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1636990056
transform 1 0 11592 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 21601
transform 1 0 12696 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 21601
transform 1 0 13248 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1636990056
transform 1 0 13432 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1636990056
transform 1 0 14536 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1636990056
transform 1 0 15640 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1636990056
transform 1 0 16744 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 21601
transform 1 0 17848 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 21601
transform 1 0 18400 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1636990056
transform 1 0 18584 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1636990056
transform 1 0 19688 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1636990056
transform 1 0 20792 0 1 1632
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1636990056
transform 1 0 21896 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 21601
transform 1 0 23000 0 1 1632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 21601
transform 1 0 23552 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_253
timestamp 21601
transform 1 0 23736 0 1 1632
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_445
timestamp 1636990056
transform 1 0 41400 0 1 1632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_457
timestamp 21601
transform 1 0 42504 0 1 1632
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1636990056
transform 1 0 736 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1636990056
transform 1 0 1840 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1636990056
transform 1 0 2944 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1636990056
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 21601
transform 1 0 5152 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 21601
transform 1 0 5520 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1636990056
transform 1 0 5704 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1636990056
transform 1 0 6808 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1636990056
transform 1 0 7912 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1636990056
transform 1 0 9016 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 21601
transform 1 0 10120 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 21601
transform 1 0 10672 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1636990056
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1636990056
transform 1 0 11960 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1636990056
transform 1 0 13064 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1636990056
transform 1 0 14168 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 21601
transform 1 0 15272 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 21601
transform 1 0 15824 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1636990056
transform 1 0 16008 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1636990056
transform 1 0 17112 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1636990056
transform 1 0 18216 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1636990056
transform 1 0 19320 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 21601
transform 1 0 20424 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 21601
transform 1 0 20976 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1636990056
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1636990056
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_249
timestamp 21601
transform 1 0 23368 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_257
timestamp 21601
transform 1 0 24104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 21601
transform 1 0 31280 0 -1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_436
timestamp 1636990056
transform 1 0 40572 0 -1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_449
timestamp 1636990056
transform 1 0 41768 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_461
timestamp 21601
transform 1 0 42872 0 -1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1636990056
transform 1 0 736 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1636990056
transform 1 0 1840 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 21601
transform 1 0 2944 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1636990056
transform 1 0 3128 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1636990056
transform 1 0 4232 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_53
timestamp 21601
transform 1 0 5336 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_57
timestamp 1636990056
transform 1 0 5704 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_69
timestamp 1636990056
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 21601
transform 1 0 7912 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1636990056
transform 1 0 8280 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1636990056
transform 1 0 9384 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_109
timestamp 21601
transform 1 0 10488 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_113
timestamp 1636990056
transform 1 0 10856 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_125
timestamp 1636990056
transform 1 0 11960 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_137
timestamp 21601
transform 1 0 13064 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1636990056
transform 1 0 13432 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1636990056
transform 1 0 14536 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 21601
transform 1 0 15640 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_169
timestamp 1636990056
transform 1 0 16008 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_181
timestamp 1636990056
transform 1 0 17112 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_193
timestamp 21601
transform 1 0 18216 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1636990056
transform 1 0 18584 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1636990056
transform 1 0 19688 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp 21601
transform 1 0 20792 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_225
timestamp 1636990056
transform 1 0 21160 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_237
timestamp 1636990056
transform 1 0 22264 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_249
timestamp 21601
transform 1 0 23368 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1636990056
transform 1 0 23736 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_265
timestamp 21601
transform 1 0 24840 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_273
timestamp 21601
transform 1 0 25576 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_301
timestamp 21601
transform 1 0 28152 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_391
timestamp 21601
transform 1 0 36432 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 21601
transform 1 0 39008 0 1 2720
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_421
timestamp 1636990056
transform 1 0 39192 0 1 2720
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_433
timestamp 1636990056
transform 1 0 40296 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_445
timestamp 21601
transform 1 0 41400 0 1 2720
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_4_449
timestamp 1636990056
transform 1 0 41768 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_461
timestamp 21601
transform 1 0 42872 0 1 2720
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1636990056
transform 1 0 736 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1636990056
transform 1 0 1840 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1636990056
transform 1 0 2944 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1636990056
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 21601
transform 1 0 5152 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 21601
transform 1 0 5520 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1636990056
transform 1 0 5704 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1636990056
transform 1 0 6808 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1636990056
transform 1 0 7912 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1636990056
transform 1 0 9016 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 21601
transform 1 0 10120 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 21601
transform 1 0 10672 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_113
timestamp 21601
transform 1 0 10856 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_117
timestamp 21601
transform 1 0 11224 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_403
timestamp 21601
transform 1 0 37536 0 -1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_411
timestamp 1636990056
transform 1 0 38272 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_423
timestamp 1636990056
transform 1 0 39376 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_435
timestamp 1636990056
transform 1 0 40480 0 -1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_447
timestamp 1636990056
transform 1 0 41584 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_459
timestamp 21601
transform 1 0 42688 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_461
timestamp 21601
transform 1 0 42872 0 -1 3808
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1636990056
transform 1 0 736 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1636990056
transform 1 0 1840 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 21601
transform 1 0 2944 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1636990056
transform 1 0 3128 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1636990056
transform 1 0 4232 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1636990056
transform 1 0 5336 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1636990056
transform 1 0 6440 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 21601
transform 1 0 7544 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 21601
transform 1 0 8096 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1636990056
transform 1 0 8280 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1636990056
transform 1 0 9384 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_109
timestamp 21601
transform 1 0 10488 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_117
timestamp 21601
transform 1 0 11224 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_357
timestamp 21601
transform 1 0 33304 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_379
timestamp 21601
transform 1 0 35328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_384
timestamp 21601
transform 1 0 35788 0 1 3808
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_400
timestamp 1636990056
transform 1 0 37260 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_412
timestamp 1636990056
transform 1 0 38364 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_424
timestamp 21601
transform 1 0 39468 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_6_433
timestamp 1636990056
transform 1 0 40296 0 1 3808
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_445
timestamp 1636990056
transform 1 0 41400 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_457
timestamp 21601
transform 1 0 42504 0 1 3808
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1636990056
transform 1 0 736 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1636990056
transform 1 0 1840 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1636990056
transform 1 0 2944 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1636990056
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 21601
transform 1 0 5152 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 21601
transform 1 0 5520 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1636990056
transform 1 0 5704 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1636990056
transform 1 0 6808 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1636990056
transform 1 0 7912 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1636990056
transform 1 0 9016 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 21601
transform 1 0 10120 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 21601
transform 1 0 10672 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_113
timestamp 21601
transform 1 0 10856 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_117
timestamp 21601
transform 1 0 11224 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_354
timestamp 21601
transform 1 0 33028 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_366
timestamp 21601
transform 1 0 34132 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_369
timestamp 21601
transform 1 0 34408 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_383
timestamp 1636990056
transform 1 0 35696 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_395
timestamp 21601
transform 1 0 36800 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_403
timestamp 21601
transform 1 0 37536 0 -1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_405
timestamp 1636990056
transform 1 0 37720 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_417
timestamp 1636990056
transform 1 0 38824 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_429
timestamp 1636990056
transform 1 0 39928 0 -1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_441
timestamp 1636990056
transform 1 0 41032 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_453
timestamp 21601
transform 1 0 42136 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_459
timestamp 21601
transform 1 0 42688 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_461
timestamp 21601
transform 1 0 42872 0 -1 4896
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1636990056
transform 1 0 736 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1636990056
transform 1 0 1840 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 21601
transform 1 0 2944 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1636990056
transform 1 0 3128 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1636990056
transform 1 0 4232 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1636990056
transform 1 0 5336 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1636990056
transform 1 0 6440 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 21601
transform 1 0 7544 0 1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 21601
transform 1 0 8096 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1636990056
transform 1 0 8280 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1636990056
transform 1 0 9384 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_109
timestamp 21601
transform 1 0 10488 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_117
timestamp 21601
transform 1 0 11224 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_359
timestamp 21601
transform 1 0 33488 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 21601
transform 1 0 33856 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_366
timestamp 21601
transform 1 0 34132 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_8_374
timestamp 21601
transform 1 0 34868 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_8_377
timestamp 21601
transform 1 0 35144 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_385
timestamp 21601
transform 1 0 35880 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_391
timestamp 1636990056
transform 1 0 36432 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_403
timestamp 1636990056
transform 1 0 37536 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_415
timestamp 1636990056
transform 1 0 38640 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_427
timestamp 21601
transform 1 0 39744 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_431
timestamp 21601
transform 1 0 40112 0 1 4896
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_433
timestamp 1636990056
transform 1 0 40296 0 1 4896
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_445
timestamp 1636990056
transform 1 0 41400 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_457
timestamp 21601
transform 1 0 42504 0 1 4896
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1636990056
transform 1 0 736 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1636990056
transform 1 0 1840 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1636990056
transform 1 0 2944 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1636990056
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 21601
transform 1 0 5152 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 21601
transform 1 0 5520 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1636990056
transform 1 0 5704 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1636990056
transform 1 0 6808 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1636990056
transform 1 0 7912 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_93
timestamp 21601
transform 1 0 9016 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_104
timestamp 21601
transform 1 0 10028 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_107
timestamp 21601
transform 1 0 10304 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 21601
transform 1 0 10580 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 21601
transform 1 0 10856 0 -1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_9_351
timestamp 1636990056
transform 1 0 32752 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_363
timestamp 1636990056
transform 1 0 33856 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_375
timestamp 1636990056
transform 1 0 34960 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_387
timestamp 1636990056
transform 1 0 36064 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_399
timestamp 21601
transform 1 0 37168 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_403
timestamp 21601
transform 1 0 37536 0 -1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_405
timestamp 1636990056
transform 1 0 37720 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_417
timestamp 1636990056
transform 1 0 38824 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_429
timestamp 1636990056
transform 1 0 39928 0 -1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_441
timestamp 1636990056
transform 1 0 41032 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_453
timestamp 21601
transform 1 0 42136 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_459
timestamp 21601
transform 1 0 42688 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_461
timestamp 21601
transform 1 0 42872 0 -1 5984
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1636990056
transform 1 0 736 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1636990056
transform 1 0 1840 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 21601
transform 1 0 2944 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1636990056
transform 1 0 3128 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1636990056
transform 1 0 4232 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_53
timestamp 21601
transform 1 0 5336 0 1 5984
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_57
timestamp 1636990056
transform 1 0 5704 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_69
timestamp 21601
transform 1 0 6808 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_72
timestamp 21601
transform 1 0 7084 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_77
timestamp 21601
transform 1 0 7544 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_81
timestamp 21601
transform 1 0 7912 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 21601
transform 1 0 8832 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_108
timestamp 21601
transform 1 0 10396 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_351
timestamp 21601
transform 1 0 32752 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_361
timestamp 21601
transform 1 0 33672 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_10_379
timestamp 21601
transform 1 0 35328 0 1 5984
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_387
timestamp 1636990056
transform 1 0 36064 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_399
timestamp 1636990056
transform 1 0 37168 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_411
timestamp 1636990056
transform 1 0 38272 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_423
timestamp 21601
transform 1 0 39376 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_431
timestamp 21601
transform 1 0 40112 0 1 5984
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_433
timestamp 1636990056
transform 1 0 40296 0 1 5984
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_445
timestamp 1636990056
transform 1 0 41400 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_457
timestamp 21601
transform 1 0 42504 0 1 5984
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1636990056
transform 1 0 736 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1636990056
transform 1 0 1840 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1636990056
transform 1 0 2944 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_39
timestamp 21601
transform 1 0 4048 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 21601
transform 1 0 5520 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_79
timestamp 21601
transform 1 0 7728 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_115
timestamp 21601
transform 1 0 11040 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_351
timestamp 21601
transform 1 0 32752 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_361
timestamp 21601
transform 1 0 33672 0 -1 7072
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_11_375
timestamp 1636990056
transform 1 0 34960 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_387
timestamp 1636990056
transform 1 0 36064 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_399
timestamp 21601
transform 1 0 37168 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_403
timestamp 21601
transform 1 0 37536 0 -1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_405
timestamp 1636990056
transform 1 0 37720 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_417
timestamp 1636990056
transform 1 0 38824 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_429
timestamp 1636990056
transform 1 0 39928 0 -1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_441
timestamp 1636990056
transform 1 0 41032 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_453
timestamp 21601
transform 1 0 42136 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_459
timestamp 21601
transform 1 0 42688 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_461
timestamp 21601
transform 1 0 42872 0 -1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1636990056
transform 1 0 736 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1636990056
transform 1 0 1840 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 21601
transform 1 0 2944 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_29
timestamp 21601
transform 1 0 3128 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_110
timestamp 21601
transform 1 0 10580 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_360
timestamp 1636990056
transform 1 0 33580 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_372
timestamp 21601
transform 1 0 34684 0 1 7072
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1636990056
transform 1 0 35144 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1636990056
transform 1 0 36248 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_401
timestamp 1636990056
transform 1 0 37352 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_413
timestamp 1636990056
transform 1 0 38456 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_425
timestamp 21601
transform 1 0 39560 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_431
timestamp 21601
transform 1 0 40112 0 1 7072
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_433
timestamp 1636990056
transform 1 0 40296 0 1 7072
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_445
timestamp 1636990056
transform 1 0 41400 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_457
timestamp 21601
transform 1 0 42504 0 1 7072
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1636990056
transform 1 0 736 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1636990056
transform 1 0 1840 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1636990056
transform 1 0 2944 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_39
timestamp 21601
transform 1 0 4048 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_53
timestamp 21601
transform 1 0 5336 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_64
timestamp 21601
transform 1 0 6348 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_115
timestamp 21601
transform 1 0 11040 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_351
timestamp 1636990056
transform 1 0 32752 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_363
timestamp 1636990056
transform 1 0 33856 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_375
timestamp 1636990056
transform 1 0 34960 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_387
timestamp 1636990056
transform 1 0 36064 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_399
timestamp 21601
transform 1 0 37168 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_403
timestamp 21601
transform 1 0 37536 0 -1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_405
timestamp 1636990056
transform 1 0 37720 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_417
timestamp 1636990056
transform 1 0 38824 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_429
timestamp 1636990056
transform 1 0 39928 0 -1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_441
timestamp 1636990056
transform 1 0 41032 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_453
timestamp 21601
transform 1 0 42136 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_459
timestamp 21601
transform 1 0 42688 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_461
timestamp 21601
transform 1 0 42872 0 -1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1636990056
transform 1 0 736 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1636990056
transform 1 0 1840 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 21601
transform 1 0 2944 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1636990056
transform 1 0 3128 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1636990056
transform 1 0 4232 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_53
timestamp 21601
transform 1 0 5336 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_59
timestamp 21601
transform 1 0 5888 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_63
timestamp 21601
transform 1 0 6256 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_66
timestamp 21601
transform 1 0 6532 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_69
timestamp 21601
transform 1 0 6808 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_75
timestamp 21601
transform 1 0 7360 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_80
timestamp 21601
transform 1 0 7820 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_89
timestamp 21601
transform 1 0 8648 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 21601
transform 1 0 9016 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_98
timestamp 21601
transform 1 0 9476 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_176
timestamp 21601
transform 1 0 16652 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 21601
transform 1 0 18400 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 21601
transform 1 0 18584 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_219
timestamp 21601
transform 1 0 20608 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_225
timestamp 21601
transform 1 0 21160 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 21601
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_292
timestamp 1636990056
transform 1 0 27324 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 21601
transform 1 0 28428 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1636990056
transform 1 0 28888 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1636990056
transform 1 0 29992 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_333
timestamp 21601
transform 1 0 31096 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_337
timestamp 1636990056
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_349
timestamp 1636990056
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_361
timestamp 21601
transform 1 0 33672 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1636990056
transform 1 0 34040 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1636990056
transform 1 0 35144 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_389
timestamp 21601
transform 1 0 36248 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_393
timestamp 1636990056
transform 1 0 36616 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_405
timestamp 1636990056
transform 1 0 37720 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_417
timestamp 21601
transform 1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_421
timestamp 1636990056
transform 1 0 39192 0 1 8160
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_433
timestamp 1636990056
transform 1 0 40296 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_445
timestamp 21601
transform 1 0 41400 0 1 8160
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_449
timestamp 1636990056
transform 1 0 41768 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_461
timestamp 21601
transform 1 0 42872 0 1 8160
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1636990056
transform 1 0 736 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1636990056
transform 1 0 1840 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1636990056
transform 1 0 2944 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1636990056
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 21601
transform 1 0 5152 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 21601
transform 1 0 5520 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1636990056
transform 1 0 5704 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1636990056
transform 1 0 6808 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1636990056
transform 1 0 7912 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1636990056
transform 1 0 9016 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_105
timestamp 21601
transform 1 0 10120 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 21601
transform 1 0 15824 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_225
timestamp 21601
transform 1 0 21160 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_240
timestamp 21601
transform 1 0 22540 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_264
timestamp 21601
transform 1 0 24748 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 21601
transform 1 0 26128 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_290
timestamp 1636990056
transform 1 0 27140 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_302
timestamp 1636990056
transform 1 0 28244 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_314
timestamp 1636990056
transform 1 0 29348 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_326
timestamp 21601
transform 1 0 30452 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_334
timestamp 21601
transform 1 0 31188 0 -1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1636990056
transform 1 0 31464 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1636990056
transform 1 0 32568 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1636990056
transform 1 0 33672 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1636990056
transform 1 0 34776 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 21601
transform 1 0 35880 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 21601
transform 1 0 36432 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1636990056
transform 1 0 36616 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_405
timestamp 1636990056
transform 1 0 37720 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_417
timestamp 1636990056
transform 1 0 38824 0 -1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_429
timestamp 1636990056
transform 1 0 39928 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 21601
transform 1 0 41032 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 21601
transform 1 0 41584 0 -1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_449
timestamp 1636990056
transform 1 0 41768 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_461
timestamp 21601
transform 1 0 42872 0 -1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1636990056
transform 1 0 736 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1636990056
transform 1 0 1840 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 21601
transform 1 0 2944 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1636990056
transform 1 0 3128 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1636990056
transform 1 0 4232 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1636990056
transform 1 0 5336 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1636990056
transform 1 0 6440 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 21601
transform 1 0 7544 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 21601
transform 1 0 8096 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1636990056
transform 1 0 8280 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1636990056
transform 1 0 9384 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1636990056
transform 1 0 10488 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1636990056
transform 1 0 11592 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_133
timestamp 21601
transform 1 0 12696 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 21601
transform 1 0 13248 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_143
timestamp 21601
transform 1 0 13616 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_146
timestamp 21601
transform 1 0 13892 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_154
timestamp 21601
transform 1 0 14628 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_216
timestamp 21601
transform 1 0 20332 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_230
timestamp 21601
transform 1 0 21620 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_237
timestamp 21601
transform 1 0 22264 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_243
timestamp 21601
transform 1 0 22816 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 21601
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_261
timestamp 21601
transform 1 0 24472 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_266
timestamp 21601
transform 1 0 24932 0 1 9248
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_274
timestamp 1636990056
transform 1 0 25668 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_286
timestamp 1636990056
transform 1 0 26772 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_298
timestamp 21601
transform 1 0 27876 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 21601
transform 1 0 28612 0 1 9248
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1636990056
transform 1 0 28888 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1636990056
transform 1 0 29992 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1636990056
transform 1 0 31096 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1636990056
transform 1 0 32200 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 21601
transform 1 0 33304 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 21601
transform 1 0 33856 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1636990056
transform 1 0 34040 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1636990056
transform 1 0 35144 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1636990056
transform 1 0 36248 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_401
timestamp 1636990056
transform 1 0 37352 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 21601
transform 1 0 38456 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 21601
transform 1 0 39008 0 1 9248
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_421
timestamp 1636990056
transform 1 0 39192 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_433
timestamp 1636990056
transform 1 0 40296 0 1 9248
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_445
timestamp 1636990056
transform 1 0 41400 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_457
timestamp 21601
transform 1 0 42504 0 1 9248
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1636990056
transform 1 0 736 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1636990056
transform 1 0 1840 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1636990056
transform 1 0 2944 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1636990056
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 21601
transform 1 0 5152 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 21601
transform 1 0 5520 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1636990056
transform 1 0 5704 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1636990056
transform 1 0 6808 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1636990056
transform 1 0 7912 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1636990056
transform 1 0 9016 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 21601
transform 1 0 10120 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 21601
transform 1 0 10672 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1636990056
transform 1 0 10856 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1636990056
transform 1 0 11960 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_137
timestamp 21601
transform 1 0 13064 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_17_147
timestamp 21601
transform 1 0 13984 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_157
timestamp 21601
transform 1 0 14904 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 21601
transform 1 0 15640 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_171
timestamp 21601
transform 1 0 16192 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_175
timestamp 21601
transform 1 0 16560 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 21601
transform 1 0 17204 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_191
timestamp 21601
transform 1 0 18032 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_194
timestamp 21601
transform 1 0 18308 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_200
timestamp 21601
transform 1 0 18860 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 21601
transform 1 0 19136 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_207
timestamp 21601
transform 1 0 19504 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_212
timestamp 21601
transform 1 0 19964 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 21601
transform 1 0 20976 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_227
timestamp 1636990056
transform 1 0 21344 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_239
timestamp 1636990056
transform 1 0 22448 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_251
timestamp 21601
transform 1 0 23552 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_259
timestamp 21601
transform 1 0 24288 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_267
timestamp 1636990056
transform 1 0 25024 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 21601
transform 1 0 26128 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_281
timestamp 21601
transform 1 0 26312 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_17_302
timestamp 21601
transform 1 0 28244 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_308
timestamp 21601
transform 1 0 28796 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_319
timestamp 21601
transform 1 0 29808 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_325
timestamp 21601
transform 1 0 30360 0 -1 10336
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_344
timestamp 1636990056
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_356
timestamp 1636990056
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_368
timestamp 1636990056
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_380
timestamp 1636990056
transform 1 0 35420 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1636990056
transform 1 0 36616 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_405
timestamp 1636990056
transform 1 0 37720 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_417
timestamp 1636990056
transform 1 0 38824 0 -1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_429
timestamp 1636990056
transform 1 0 39928 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 21601
transform 1 0 41032 0 -1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 21601
transform 1 0 41584 0 -1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_449
timestamp 1636990056
transform 1 0 41768 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_461
timestamp 21601
transform 1 0 42872 0 -1 10336
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1636990056
transform 1 0 736 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1636990056
transform 1 0 1840 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 21601
transform 1 0 2944 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1636990056
transform 1 0 3128 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1636990056
transform 1 0 4232 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1636990056
transform 1 0 5336 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1636990056
transform 1 0 6440 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 21601
transform 1 0 7544 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 21601
transform 1 0 8096 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1636990056
transform 1 0 8280 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1636990056
transform 1 0 9384 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1636990056
transform 1 0 10488 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1636990056
transform 1 0 11592 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 21601
transform 1 0 12696 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 21601
transform 1 0 13248 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1636990056
transform 1 0 13432 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1636990056
transform 1 0 14536 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1636990056
transform 1 0 15640 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1636990056
transform 1 0 16744 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 21601
transform 1 0 17848 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 21601
transform 1 0 18400 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1636990056
transform 1 0 18584 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1636990056
transform 1 0 19688 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1636990056
transform 1 0 20792 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1636990056
transform 1 0 21896 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 21601
transform 1 0 23000 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 21601
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 21601
transform 1 0 23736 0 1 10336
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_18_274
timestamp 1636990056
transform 1 0 25668 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_286
timestamp 21601
transform 1 0 26772 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_299
timestamp 21601
transform 1 0 27968 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 21601
transform 1 0 28704 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1636990056
transform 1 0 28888 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1636990056
transform 1 0 29992 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_333
timestamp 21601
transform 1 0 31096 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_341
timestamp 21601
transform 1 0 31832 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_347
timestamp 1636990056
transform 1 0 32384 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_359
timestamp 21601
transform 1 0 33488 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 21601
transform 1 0 33856 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1636990056
transform 1 0 34040 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1636990056
transform 1 0 35144 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_389
timestamp 1636990056
transform 1 0 36248 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_401
timestamp 1636990056
transform 1 0 37352 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 21601
transform 1 0 38456 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 21601
transform 1 0 39008 0 1 10336
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_421
timestamp 1636990056
transform 1 0 39192 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_433
timestamp 1636990056
transform 1 0 40296 0 1 10336
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_445
timestamp 1636990056
transform 1 0 41400 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_457
timestamp 21601
transform 1 0 42504 0 1 10336
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1636990056
transform 1 0 736 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1636990056
transform 1 0 1840 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_27
timestamp 21601
transform 1 0 2944 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_29
timestamp 1636990056
transform 1 0 3128 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_41
timestamp 1636990056
transform 1 0 4232 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_53
timestamp 21601
transform 1 0 5336 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1636990056
transform 1 0 5704 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1636990056
transform 1 0 6808 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_81
timestamp 21601
transform 1 0 7912 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_85
timestamp 1636990056
transform 1 0 8280 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_97
timestamp 1636990056
transform 1 0 9384 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 21601
transform 1 0 10488 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1636990056
transform 1 0 10856 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1636990056
transform 1 0 11960 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_137
timestamp 21601
transform 1 0 13064 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_141
timestamp 1636990056
transform 1 0 13432 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_153
timestamp 1636990056
transform 1 0 14536 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 21601
transform 1 0 15640 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1636990056
transform 1 0 16008 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1636990056
transform 1 0 17112 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_193
timestamp 21601
transform 1 0 18216 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_197
timestamp 1636990056
transform 1 0 18584 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_209
timestamp 1636990056
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_221
timestamp 21601
transform 1 0 20792 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1636990056
transform 1 0 21160 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1636990056
transform 1 0 22264 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_249
timestamp 21601
transform 1 0 23368 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_253
timestamp 21601
transform 1 0 23736 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_262
timestamp 21601
transform 1 0 24564 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_270
timestamp 21601
transform 1 0 25300 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_275
timestamp 21601
transform 1 0 25760 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 21601
transform 1 0 26128 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_290
timestamp 21601
transform 1 0 27140 0 -1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_296
timestamp 21601
transform 1 0 27692 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_313
timestamp 21601
transform 1 0 29256 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 21601
transform 1 0 31280 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_342
timestamp 21601
transform 1 0 31924 0 -1 11424
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_367
timestamp 1636990056
transform 1 0 34224 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_379
timestamp 1636990056
transform 1 0 35328 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 21601
transform 1 0 36432 0 -1 11424
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1636990056
transform 1 0 36616 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_405
timestamp 1636990056
transform 1 0 37720 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_417
timestamp 21601
transform 1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_421
timestamp 1636990056
transform 1 0 39192 0 -1 11424
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_433
timestamp 1636990056
transform 1 0 40296 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_445
timestamp 21601
transform 1 0 41400 0 -1 11424
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_449
timestamp 1636990056
transform 1 0 41768 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_461
timestamp 21601
transform 1 0 42872 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  hreadyout_ack_gate
timestamp 21601
transform 1 0 33120 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[0\]
timestamp 21601
transform 1 0 33948 0 -1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[1\]
timestamp 21601
transform 1 0 34224 0 1 5984
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[2\]
timestamp 21601
transform 1 0 34500 0 -1 4896
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[3\]
timestamp 21601
transform 1 0 34776 0 -1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[4\]
timestamp 21601
transform 1 0 35512 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[5\]
timestamp 21601
transform 1 0 36616 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[6\]
timestamp 21601
transform 1 0 37444 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[7\]
timestamp 21601
transform 1 0 36984 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[8\]
timestamp 21601
transform 1 0 36616 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[9\]
timestamp 21601
transform 1 0 36616 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[10\]
timestamp 21601
transform 1 0 37444 0 -1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[11\]
timestamp 21601
transform 1 0 37812 0 1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[12\]
timestamp 21601
transform 1 0 38272 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[13\]
timestamp 21601
transform 1 0 38088 0 1 544
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[14\]
timestamp 21601
transform 1 0 39100 0 -1 1632
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  irq_gates\[15\]
timestamp 21601
transform 1 0 39928 0 -1 1632
box -38 -48 866 592
use vccd1_tie_high  mprj_logic_high_inst
timestamp 0
transform 1 0 12000 0 1 4000
box 0 0 1 1
use sky130_fd_sc_hd__buf_12  output1
timestamp 21601
transform 1 0 23736 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output2
timestamp 21601
transform 1 0 28888 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output3
timestamp 21601
transform -1 0 27784 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output4
timestamp 21601
transform 1 0 29256 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output5
timestamp 21601
transform -1 0 29256 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output6
timestamp 21601
transform -1 0 30360 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output7
timestamp 21601
transform 1 0 31464 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output8
timestamp 21601
transform 1 0 29256 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output9
timestamp 21601
transform 1 0 30360 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output10
timestamp 21601
transform -1 0 30360 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output11
timestamp 21601
transform 1 0 31464 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output12
timestamp 21601
transform 1 0 23552 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output13
timestamp 21601
transform 1 0 31832 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output14
timestamp 21601
transform 1 0 31464 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output15
timestamp 21601
transform 1 0 32936 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output16
timestamp 21601
transform 1 0 34040 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output17
timestamp 21601
transform -1 0 32936 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output18
timestamp 21601
transform 1 0 34408 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output19
timestamp 21601
transform 1 0 32936 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output20
timestamp 21601
transform 1 0 34040 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 21601
transform 1 0 32752 0 -1 3808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 21601
transform 1 0 36616 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 21601
transform -1 0 25300 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 21601
transform 1 0 34408 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 21601
transform 1 0 34040 0 1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 21601
transform 1 0 26312 0 1 544
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 21601
transform -1 0 25852 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 21601
transform 1 0 25300 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 21601
transform 1 0 26312 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 21601
transform 1 0 26772 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 21601
transform -1 0 27784 0 -1 2720
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 21601
transform 1 0 27784 0 -1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 21601
transform 1 0 35512 0 1 1632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_20
timestamp 21601
transform 1 0 460 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 21601
transform -1 0 43516 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_21
timestamp 21601
transform 1 0 460 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 21601
transform -1 0 43516 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_22
timestamp 21601
transform 1 0 460 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 21601
transform -1 0 43516 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_23
timestamp 21601
transform 1 0 460 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 21601
transform -1 0 43516 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_24
timestamp 21601
transform 1 0 460 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 21601
transform -1 0 43516 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Left_39
timestamp 21601
transform 1 0 460 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_1_Right_57
timestamp 21601
transform -1 0 11592 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Left_40
timestamp 21601
transform 1 0 32476 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_2_Right_11
timestamp 21601
transform -1 0 43516 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Left_25
timestamp 21601
transform 1 0 460 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_1_Right_49
timestamp 21601
transform -1 0 11592 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Left_41
timestamp 21601
transform 1 0 32476 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_2_Right_12
timestamp 21601
transform -1 0 43516 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Left_26
timestamp 21601
transform 1 0 460 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_1_Right_50
timestamp 21601
transform -1 0 11592 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Left_42
timestamp 21601
transform 1 0 32476 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_2_Right_13
timestamp 21601
transform -1 0 43516 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Left_27
timestamp 21601
transform 1 0 460 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_1_Right_51
timestamp 21601
transform -1 0 11592 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Left_43
timestamp 21601
transform 1 0 32476 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_2_Right_14
timestamp 21601
transform -1 0 43516 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Left_28
timestamp 21601
transform 1 0 460 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_1_Right_52
timestamp 21601
transform -1 0 11592 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Left_44
timestamp 21601
transform 1 0 32476 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_2_Right_15
timestamp 21601
transform -1 0 43516 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Left_29
timestamp 21601
transform 1 0 460 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_1_Right_53
timestamp 21601
transform -1 0 11592 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Left_45
timestamp 21601
transform 1 0 32476 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_2_Right_16
timestamp 21601
transform -1 0 43516 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Left_30
timestamp 21601
transform 1 0 460 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_1_Right_54
timestamp 21601
transform -1 0 11592 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Left_46
timestamp 21601
transform 1 0 32476 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_2_Right_17
timestamp 21601
transform -1 0 43516 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Left_31
timestamp 21601
transform 1 0 460 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_1_Right_55
timestamp 21601
transform -1 0 11592 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Left_47
timestamp 21601
transform 1 0 32476 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_2_Right_18
timestamp 21601
transform -1 0 43516 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Left_32
timestamp 21601
transform 1 0 460 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_1_Right_56
timestamp 21601
transform -1 0 11592 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Left_48
timestamp 21601
transform 1 0 32476 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_2_Right_19
timestamp 21601
transform -1 0 43516 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_33
timestamp 21601
transform 1 0 460 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_5
timestamp 21601
transform -1 0 43516 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_34
timestamp 21601
transform 1 0 460 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_6
timestamp 21601
transform -1 0 43516 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_35
timestamp 21601
transform 1 0 460 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_7
timestamp 21601
transform -1 0 43516 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_36
timestamp 21601
transform 1 0 460 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_8
timestamp 21601
transform -1 0 43516 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_37
timestamp 21601
transform 1 0 460 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_9
timestamp 21601
transform -1 0 43516 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_38
timestamp 21601
transform 1 0 460 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_10
timestamp 21601
transform -1 0 43516 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_58
timestamp 21601
transform 1 0 3036 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_59
timestamp 21601
transform 1 0 5612 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_60
timestamp 21601
transform 1 0 8188 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_61
timestamp 21601
transform 1 0 10764 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62
timestamp 21601
transform 1 0 13340 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 21601
transform 1 0 15916 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 21601
transform 1 0 18492 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 21601
transform 1 0 21068 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 21601
transform 1 0 23644 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 21601
transform 1 0 26220 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp 21601
transform 1 0 28796 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 21601
transform 1 0 31372 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 21601
transform 1 0 33948 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 21601
transform 1 0 36524 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 21601
transform 1 0 39100 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_73
timestamp 21601
transform 1 0 41676 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_74
timestamp 21601
transform 1 0 5612 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 21601
transform 1 0 10764 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 21601
transform 1 0 15916 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_77
timestamp 21601
transform 1 0 21068 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_78
timestamp 21601
transform 1 0 26220 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_79
timestamp 21601
transform 1 0 31372 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_80
timestamp 21601
transform 1 0 36524 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_81
timestamp 21601
transform 1 0 41676 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_82
timestamp 21601
transform 1 0 3036 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_83
timestamp 21601
transform 1 0 8188 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_84
timestamp 21601
transform 1 0 13340 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_85
timestamp 21601
transform 1 0 18492 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_86
timestamp 21601
transform 1 0 23644 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_87
timestamp 21601
transform 1 0 28796 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_88
timestamp 21601
transform 1 0 33948 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_89
timestamp 21601
transform 1 0 39100 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_90
timestamp 21601
transform 1 0 5612 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_91
timestamp 21601
transform 1 0 10764 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_92
timestamp 21601
transform 1 0 15916 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_93
timestamp 21601
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_94
timestamp 21601
transform 1 0 26220 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_95
timestamp 21601
transform 1 0 31372 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_96
timestamp 21601
transform 1 0 36524 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_97
timestamp 21601
transform 1 0 41676 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_98
timestamp 21601
transform 1 0 3036 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_99
timestamp 21601
transform 1 0 5612 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_100
timestamp 21601
transform 1 0 8188 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_101
timestamp 21601
transform 1 0 10764 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_102
timestamp 21601
transform 1 0 13340 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_103
timestamp 21601
transform 1 0 15916 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_104
timestamp 21601
transform 1 0 18492 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_105
timestamp 21601
transform 1 0 21068 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_106
timestamp 21601
transform 1 0 23644 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_107
timestamp 21601
transform 1 0 26220 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_108
timestamp 21601
transform 1 0 28796 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_109
timestamp 21601
transform 1 0 31372 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_110
timestamp 21601
transform 1 0 33948 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_111
timestamp 21601
transform 1 0 36524 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_112
timestamp 21601
transform 1 0 39100 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_113
timestamp 21601
transform 1 0 41676 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1_194
timestamp 21601
transform 1 0 5612 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_1_195
timestamp 21601
transform 1 0 10764 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_2_196
timestamp 21601
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_2_197
timestamp 21601
transform 1 0 42780 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1_114
timestamp 21601
transform 1 0 3036 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_1_115
timestamp 21601
transform 1 0 8188 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_2_198
timestamp 21601
transform 1 0 35052 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_2_199
timestamp 21601
transform 1 0 40204 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1_116
timestamp 21601
transform 1 0 5612 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_1_117
timestamp 21601
transform 1 0 10764 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_2_200
timestamp 21601
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_2_201
timestamp 21601
transform 1 0 42780 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1_118
timestamp 21601
transform 1 0 3036 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_1_119
timestamp 21601
transform 1 0 8188 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_2_202
timestamp 21601
transform 1 0 35052 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_2_203
timestamp 21601
transform 1 0 40204 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1_120
timestamp 21601
transform 1 0 5612 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_1_121
timestamp 21601
transform 1 0 10764 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_2_204
timestamp 21601
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_2_205
timestamp 21601
transform 1 0 42780 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_122
timestamp 21601
transform 1 0 3036 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_1_123
timestamp 21601
transform 1 0 8188 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_206
timestamp 21601
transform 1 0 35052 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_2_207
timestamp 21601
transform 1 0 40204 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_1_124
timestamp 21601
transform 1 0 5612 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_1_125
timestamp 21601
transform 1 0 10764 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_208
timestamp 21601
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_2_209
timestamp 21601
transform 1 0 42780 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_126
timestamp 21601
transform 1 0 3036 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_1_127
timestamp 21601
transform 1 0 8188 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_210
timestamp 21601
transform 1 0 35052 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_2_211
timestamp 21601
transform 1 0 40204 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_1_128
timestamp 21601
transform 1 0 5612 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_1_129
timestamp 21601
transform 1 0 10764 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_212
timestamp 21601
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_2_213
timestamp 21601
transform 1 0 42780 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_130
timestamp 21601
transform 1 0 3036 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_131
timestamp 21601
transform 1 0 5612 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_132
timestamp 21601
transform 1 0 8188 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_133
timestamp 21601
transform 1 0 10764 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_134
timestamp 21601
transform 1 0 13340 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_135
timestamp 21601
transform 1 0 15916 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_136
timestamp 21601
transform 1 0 18492 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_137
timestamp 21601
transform 1 0 21068 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_138
timestamp 21601
transform 1 0 23644 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_139
timestamp 21601
transform 1 0 26220 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_140
timestamp 21601
transform 1 0 28796 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_141
timestamp 21601
transform 1 0 31372 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_142
timestamp 21601
transform 1 0 33948 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_143
timestamp 21601
transform 1 0 36524 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_144
timestamp 21601
transform 1 0 39100 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_145
timestamp 21601
transform 1 0 41676 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_146
timestamp 21601
transform 1 0 5612 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_147
timestamp 21601
transform 1 0 10764 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_148
timestamp 21601
transform 1 0 15916 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_149
timestamp 21601
transform 1 0 21068 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_150
timestamp 21601
transform 1 0 26220 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_151
timestamp 21601
transform 1 0 31372 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_152
timestamp 21601
transform 1 0 36524 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_153
timestamp 21601
transform 1 0 41676 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_154
timestamp 21601
transform 1 0 3036 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_155
timestamp 21601
transform 1 0 8188 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_156
timestamp 21601
transform 1 0 13340 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_157
timestamp 21601
transform 1 0 18492 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_158
timestamp 21601
transform 1 0 23644 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_159
timestamp 21601
transform 1 0 28796 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_160
timestamp 21601
transform 1 0 33948 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_161
timestamp 21601
transform 1 0 39100 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_162
timestamp 21601
transform 1 0 5612 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_163
timestamp 21601
transform 1 0 10764 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_164
timestamp 21601
transform 1 0 15916 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_165
timestamp 21601
transform 1 0 21068 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_166
timestamp 21601
transform 1 0 26220 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_167
timestamp 21601
transform 1 0 31372 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_168
timestamp 21601
transform 1 0 36524 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_169
timestamp 21601
transform 1 0 41676 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_170
timestamp 21601
transform 1 0 3036 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_171
timestamp 21601
transform 1 0 8188 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_172
timestamp 21601
transform 1 0 13340 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_173
timestamp 21601
transform 1 0 18492 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_174
timestamp 21601
transform 1 0 23644 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_175
timestamp 21601
transform 1 0 28796 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_176
timestamp 21601
transform 1 0 33948 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_177
timestamp 21601
transform 1 0 39100 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_178
timestamp 21601
transform 1 0 3036 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_179
timestamp 21601
transform 1 0 5612 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_180
timestamp 21601
transform 1 0 8188 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_181
timestamp 21601
transform 1 0 10764 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_182
timestamp 21601
transform 1 0 13340 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_183
timestamp 21601
transform 1 0 15916 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_184
timestamp 21601
transform 1 0 18492 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_185
timestamp 21601
transform 1 0 21068 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_186
timestamp 21601
transform 1 0 23644 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_187
timestamp 21601
transform 1 0 26220 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_188
timestamp 21601
transform 1 0 28796 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_189
timestamp 21601
transform 1 0 31372 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_190
timestamp 21601
transform 1 0 33948 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_191
timestamp 21601
transform 1 0 36524 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_192
timestamp 21601
transform 1 0 39100 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_193
timestamp 21601
transform 1 0 41676 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[0\]
timestamp 21601
transform -1 0 24380 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[1\]
timestamp 21601
transform 1 0 24288 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[2\]
timestamp 21601
transform 1 0 24564 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[3\]
timestamp 21601
transform 1 0 24748 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[4\]
timestamp 21601
transform 1 0 25024 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[5\]
timestamp 21601
transform 1 0 25484 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[6\]
timestamp 21601
transform 1 0 25852 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[7\]
timestamp 21601
transform 1 0 26312 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[8\]
timestamp 21601
transform 1 0 26680 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[9\]
timestamp 21601
transform 1 0 26864 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[10\]
timestamp 21601
transform 1 0 27140 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[11\]
timestamp 21601
transform 1 0 27416 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[12\]
timestamp 21601
transform 1 0 27508 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[13\]
timestamp 21601
transform 1 0 27784 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[14\]
timestamp 21601
transform 1 0 28060 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[15\]
timestamp 21601
transform 1 0 28152 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[16\]
timestamp 21601
transform 1 0 28520 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[17\]
timestamp 21601
transform 1 0 28888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[18\]
timestamp 21601
transform 1 0 29164 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[19\]
timestamp 21601
transform 1 0 29440 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[20\]
timestamp 21601
transform 1 0 29716 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[21\]
timestamp 21601
transform 1 0 29900 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[22\]
timestamp 21601
transform 1 0 30360 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[23\]
timestamp 21601
transform 1 0 30636 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[24\]
timestamp 21601
transform 1 0 30636 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[25\]
timestamp 21601
transform 1 0 30912 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[26\]
timestamp 21601
transform 1 0 31464 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[27\]
timestamp 21601
transform 1 0 31648 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[28\]
timestamp 21601
transform 1 0 31924 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[29\]
timestamp 21601
transform 1 0 32292 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[30\]
timestamp 21601
transform 1 0 32568 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  wb_hrdata_gates\[31\]
timestamp 21601
transform 1 0 32844 0 -1 11424
box -38 -48 314 592
<< labels >>
flabel metal2 s 3054 0 3110 400 0 FreeSans 224 90 0 0 frigate_HCLK
port 0 nsew signal input
flabel metal2 s 2778 0 2834 400 0 FreeSans 224 90 0 0 frigate_HRESETn
port 1 nsew signal input
flabel metal2 s 32310 0 32366 400 0 FreeSans 224 90 0 0 mprj_AHB_Ena
port 2 nsew signal input
flabel metal2 s 4986 0 5042 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[0]
port 3 nsew signal input
flabel metal2 s 7746 0 7802 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[10]
port 4 nsew signal input
flabel metal2 s 8022 0 8078 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[11]
port 5 nsew signal input
flabel metal2 s 8298 0 8354 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[12]
port 6 nsew signal input
flabel metal2 s 8574 0 8630 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[13]
port 7 nsew signal input
flabel metal2 s 8850 0 8906 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[14]
port 8 nsew signal input
flabel metal2 s 9126 0 9182 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[15]
port 9 nsew signal input
flabel metal2 s 9402 0 9458 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[16]
port 10 nsew signal input
flabel metal2 s 9678 0 9734 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[17]
port 11 nsew signal input
flabel metal2 s 9954 0 10010 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[18]
port 12 nsew signal input
flabel metal2 s 10230 0 10286 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[19]
port 13 nsew signal input
flabel metal2 s 5262 0 5318 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[1]
port 14 nsew signal input
flabel metal2 s 10506 0 10562 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[20]
port 15 nsew signal input
flabel metal2 s 10782 0 10838 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[21]
port 16 nsew signal input
flabel metal2 s 11058 0 11114 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[22]
port 17 nsew signal input
flabel metal2 s 11334 0 11390 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[23]
port 18 nsew signal input
flabel metal2 s 11610 0 11666 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[24]
port 19 nsew signal input
flabel metal2 s 11886 0 11942 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[25]
port 20 nsew signal input
flabel metal2 s 12162 0 12218 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[26]
port 21 nsew signal input
flabel metal2 s 12438 0 12494 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[27]
port 22 nsew signal input
flabel metal2 s 12714 0 12770 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[28]
port 23 nsew signal input
flabel metal2 s 12990 0 13046 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[29]
port 24 nsew signal input
flabel metal2 s 5538 0 5594 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[2]
port 25 nsew signal input
flabel metal2 s 13266 0 13322 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[30]
port 26 nsew signal input
flabel metal2 s 13542 0 13598 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[31]
port 27 nsew signal input
flabel metal2 s 5814 0 5870 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[3]
port 28 nsew signal input
flabel metal2 s 6090 0 6146 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[4]
port 29 nsew signal input
flabel metal2 s 6366 0 6422 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[5]
port 30 nsew signal input
flabel metal2 s 6642 0 6698 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[6]
port 31 nsew signal input
flabel metal2 s 6918 0 6974 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[7]
port 32 nsew signal input
flabel metal2 s 7194 0 7250 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[8]
port 33 nsew signal input
flabel metal2 s 7470 0 7526 400 0 FreeSans 224 90 0 0 mprj_HADDR_core[9]
port 34 nsew signal input
flabel metal2 s 7286 11600 7342 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[0]
port 35 nsew signal output
flabel metal2 s 10046 11600 10102 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[10]
port 36 nsew signal output
flabel metal2 s 10322 11600 10378 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[11]
port 37 nsew signal output
flabel metal2 s 10598 11600 10654 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[12]
port 38 nsew signal output
flabel metal2 s 10874 11600 10930 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[13]
port 39 nsew signal output
flabel metal2 s 11150 11600 11206 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[14]
port 40 nsew signal output
flabel metal2 s 11426 11600 11482 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[15]
port 41 nsew signal output
flabel metal2 s 11702 11600 11758 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[16]
port 42 nsew signal output
flabel metal2 s 11978 11600 12034 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[17]
port 43 nsew signal output
flabel metal2 s 12254 11600 12310 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[18]
port 44 nsew signal output
flabel metal2 s 12530 11600 12586 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[19]
port 45 nsew signal output
flabel metal2 s 7562 11600 7618 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[1]
port 46 nsew signal output
flabel metal2 s 12806 11600 12862 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[20]
port 47 nsew signal output
flabel metal2 s 13082 11600 13138 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[21]
port 48 nsew signal output
flabel metal2 s 13358 11600 13414 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[22]
port 49 nsew signal output
flabel metal2 s 13634 11600 13690 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[23]
port 50 nsew signal output
flabel metal2 s 13910 11600 13966 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[24]
port 51 nsew signal output
flabel metal2 s 14186 11600 14242 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[25]
port 52 nsew signal output
flabel metal2 s 14462 11600 14518 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[26]
port 53 nsew signal output
flabel metal2 s 14738 11600 14794 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[27]
port 54 nsew signal output
flabel metal2 s 15014 11600 15070 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[28]
port 55 nsew signal output
flabel metal2 s 15290 11600 15346 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[29]
port 56 nsew signal output
flabel metal2 s 7838 11600 7894 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[2]
port 57 nsew signal output
flabel metal2 s 15566 11600 15622 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[30]
port 58 nsew signal output
flabel metal2 s 15842 11600 15898 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[31]
port 59 nsew signal output
flabel metal2 s 8114 11600 8170 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[3]
port 60 nsew signal output
flabel metal2 s 8390 11600 8446 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[4]
port 61 nsew signal output
flabel metal2 s 8666 11600 8722 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[5]
port 62 nsew signal output
flabel metal2 s 8942 11600 8998 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[6]
port 63 nsew signal output
flabel metal2 s 9218 11600 9274 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[7]
port 64 nsew signal output
flabel metal2 s 9494 11600 9550 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[8]
port 65 nsew signal output
flabel metal2 s 9770 11600 9826 12000 0 FreeSans 224 90 0 0 mprj_HADDR_user[9]
port 66 nsew signal output
flabel metal2 s 23202 0 23258 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[0]
port 67 nsew signal output
flabel metal2 s 25962 0 26018 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[10]
port 68 nsew signal output
flabel metal2 s 26238 0 26294 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[11]
port 69 nsew signal output
flabel metal2 s 26514 0 26570 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[12]
port 70 nsew signal output
flabel metal2 s 26790 0 26846 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[13]
port 71 nsew signal output
flabel metal2 s 27066 0 27122 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[14]
port 72 nsew signal output
flabel metal2 s 27342 0 27398 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[15]
port 73 nsew signal output
flabel metal2 s 27618 0 27674 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[16]
port 74 nsew signal output
flabel metal2 s 27894 0 27950 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[17]
port 75 nsew signal output
flabel metal2 s 28170 0 28226 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[18]
port 76 nsew signal output
flabel metal2 s 28446 0 28502 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[19]
port 77 nsew signal output
flabel metal2 s 23478 0 23534 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[1]
port 78 nsew signal output
flabel metal2 s 28722 0 28778 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[20]
port 79 nsew signal output
flabel metal2 s 28998 0 29054 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[21]
port 80 nsew signal output
flabel metal2 s 29274 0 29330 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[22]
port 81 nsew signal output
flabel metal2 s 29550 0 29606 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[23]
port 82 nsew signal output
flabel metal2 s 29826 0 29882 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[24]
port 83 nsew signal output
flabel metal2 s 30102 0 30158 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[25]
port 84 nsew signal output
flabel metal2 s 30378 0 30434 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[26]
port 85 nsew signal output
flabel metal2 s 30654 0 30710 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[27]
port 86 nsew signal output
flabel metal2 s 30930 0 30986 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[28]
port 87 nsew signal output
flabel metal2 s 31206 0 31262 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[29]
port 88 nsew signal output
flabel metal2 s 23754 0 23810 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[2]
port 89 nsew signal output
flabel metal2 s 31482 0 31538 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[30]
port 90 nsew signal output
flabel metal2 s 31758 0 31814 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[31]
port 91 nsew signal output
flabel metal2 s 24030 0 24086 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[3]
port 92 nsew signal output
flabel metal2 s 24306 0 24362 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[4]
port 93 nsew signal output
flabel metal2 s 24582 0 24638 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[5]
port 94 nsew signal output
flabel metal2 s 24858 0 24914 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[6]
port 95 nsew signal output
flabel metal2 s 25134 0 25190 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[7]
port 96 nsew signal output
flabel metal2 s 25410 0 25466 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[8]
port 97 nsew signal output
flabel metal2 s 25686 0 25742 400 0 FreeSans 224 90 0 0 mprj_HRDATA_core[9]
port 98 nsew signal output
flabel metal2 s 25502 11600 25558 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[0]
port 99 nsew signal input
flabel metal2 s 28262 11600 28318 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[10]
port 100 nsew signal input
flabel metal2 s 28538 11600 28594 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[11]
port 101 nsew signal input
flabel metal2 s 28814 11600 28870 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[12]
port 102 nsew signal input
flabel metal2 s 29090 11600 29146 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[13]
port 103 nsew signal input
flabel metal2 s 29366 11600 29422 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[14]
port 104 nsew signal input
flabel metal2 s 29642 11600 29698 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[15]
port 105 nsew signal input
flabel metal2 s 29918 11600 29974 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[16]
port 106 nsew signal input
flabel metal2 s 30194 11600 30250 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[17]
port 107 nsew signal input
flabel metal2 s 30470 11600 30526 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[18]
port 108 nsew signal input
flabel metal2 s 30746 11600 30802 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[19]
port 109 nsew signal input
flabel metal2 s 25778 11600 25834 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[1]
port 110 nsew signal input
flabel metal2 s 31022 11600 31078 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[20]
port 111 nsew signal input
flabel metal2 s 31298 11600 31354 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[21]
port 112 nsew signal input
flabel metal2 s 31574 11600 31630 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[22]
port 113 nsew signal input
flabel metal2 s 31850 11600 31906 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[23]
port 114 nsew signal input
flabel metal2 s 32126 11600 32182 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[24]
port 115 nsew signal input
flabel metal2 s 32402 11600 32458 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[25]
port 116 nsew signal input
flabel metal2 s 32678 11600 32734 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[26]
port 117 nsew signal input
flabel metal2 s 32954 11600 33010 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[27]
port 118 nsew signal input
flabel metal2 s 33230 11600 33286 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[28]
port 119 nsew signal input
flabel metal2 s 33506 11600 33562 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[29]
port 120 nsew signal input
flabel metal2 s 26054 11600 26110 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[2]
port 121 nsew signal input
flabel metal2 s 33782 11600 33838 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[30]
port 122 nsew signal input
flabel metal2 s 34058 11600 34114 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[31]
port 123 nsew signal input
flabel metal2 s 26330 11600 26386 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[3]
port 124 nsew signal input
flabel metal2 s 26606 11600 26662 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[4]
port 125 nsew signal input
flabel metal2 s 26882 11600 26938 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[5]
port 126 nsew signal input
flabel metal2 s 27158 11600 27214 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[6]
port 127 nsew signal input
flabel metal2 s 27434 11600 27490 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[7]
port 128 nsew signal input
flabel metal2 s 27710 11600 27766 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[8]
port 129 nsew signal input
flabel metal2 s 27986 11600 28042 12000 0 FreeSans 224 90 0 0 mprj_HRDATA_user[9]
port 130 nsew signal input
flabel metal2 s 32034 0 32090 400 0 FreeSans 224 90 0 0 mprj_HREADYOUT_core
port 131 nsew signal output
flabel metal2 s 34334 11600 34390 12000 0 FreeSans 224 90 0 0 mprj_HREADYOUT_user
port 132 nsew signal input
flabel metal2 s 3606 0 3662 400 0 FreeSans 224 90 0 0 mprj_HREADY_core
port 133 nsew signal input
flabel metal2 s 5906 11600 5962 12000 0 FreeSans 224 90 0 0 mprj_HREADY_user
port 134 nsew signal output
flabel metal2 s 3330 0 3386 400 0 FreeSans 224 90 0 0 mprj_HSEL_core
port 135 nsew signal input
flabel metal2 s 5630 11600 5686 12000 0 FreeSans 224 90 0 0 mprj_HSEL_user
port 136 nsew signal output
flabel metal2 s 4158 0 4214 400 0 FreeSans 224 90 0 0 mprj_HSIZE_core[0]
port 137 nsew signal input
flabel metal2 s 4434 0 4490 400 0 FreeSans 224 90 0 0 mprj_HSIZE_core[1]
port 138 nsew signal input
flabel metal2 s 4710 0 4766 400 0 FreeSans 224 90 0 0 mprj_HSIZE_core[2]
port 139 nsew signal input
flabel metal2 s 6458 11600 6514 12000 0 FreeSans 224 90 0 0 mprj_HSIZE_user[0]
port 140 nsew signal output
flabel metal2 s 6734 11600 6790 12000 0 FreeSans 224 90 0 0 mprj_HSIZE_user[1]
port 141 nsew signal output
flabel metal2 s 7010 11600 7066 12000 0 FreeSans 224 90 0 0 mprj_HSIZE_user[2]
port 142 nsew signal output
flabel metal2 s 22650 0 22706 400 0 FreeSans 224 90 0 0 mprj_HTRANS_core[0]
port 143 nsew signal input
flabel metal2 s 22926 0 22982 400 0 FreeSans 224 90 0 0 mprj_HTRANS_core[1]
port 144 nsew signal input
flabel metal2 s 24950 11600 25006 12000 0 FreeSans 224 90 0 0 mprj_HTRANS_user[0]
port 145 nsew signal output
flabel metal2 s 25226 11600 25282 12000 0 FreeSans 224 90 0 0 mprj_HTRANS_user[1]
port 146 nsew signal output
flabel metal2 s 13818 0 13874 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[0]
port 147 nsew signal input
flabel metal2 s 16578 0 16634 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[10]
port 148 nsew signal input
flabel metal2 s 16854 0 16910 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[11]
port 149 nsew signal input
flabel metal2 s 17130 0 17186 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[12]
port 150 nsew signal input
flabel metal2 s 17406 0 17462 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[13]
port 151 nsew signal input
flabel metal2 s 17682 0 17738 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[14]
port 152 nsew signal input
flabel metal2 s 17958 0 18014 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[15]
port 153 nsew signal input
flabel metal2 s 18234 0 18290 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[16]
port 154 nsew signal input
flabel metal2 s 18510 0 18566 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[17]
port 155 nsew signal input
flabel metal2 s 18786 0 18842 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[18]
port 156 nsew signal input
flabel metal2 s 19062 0 19118 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[19]
port 157 nsew signal input
flabel metal2 s 14094 0 14150 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[1]
port 158 nsew signal input
flabel metal2 s 19338 0 19394 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[20]
port 159 nsew signal input
flabel metal2 s 19614 0 19670 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[21]
port 160 nsew signal input
flabel metal2 s 19890 0 19946 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[22]
port 161 nsew signal input
flabel metal2 s 20166 0 20222 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[23]
port 162 nsew signal input
flabel metal2 s 20442 0 20498 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[24]
port 163 nsew signal input
flabel metal2 s 20718 0 20774 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[25]
port 164 nsew signal input
flabel metal2 s 20994 0 21050 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[26]
port 165 nsew signal input
flabel metal2 s 21270 0 21326 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[27]
port 166 nsew signal input
flabel metal2 s 21546 0 21602 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[28]
port 167 nsew signal input
flabel metal2 s 21822 0 21878 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[29]
port 168 nsew signal input
flabel metal2 s 14370 0 14426 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[2]
port 169 nsew signal input
flabel metal2 s 22098 0 22154 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[30]
port 170 nsew signal input
flabel metal2 s 22374 0 22430 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[31]
port 171 nsew signal input
flabel metal2 s 14646 0 14702 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[3]
port 172 nsew signal input
flabel metal2 s 14922 0 14978 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[4]
port 173 nsew signal input
flabel metal2 s 15198 0 15254 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[5]
port 174 nsew signal input
flabel metal2 s 15474 0 15530 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[6]
port 175 nsew signal input
flabel metal2 s 15750 0 15806 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[7]
port 176 nsew signal input
flabel metal2 s 16026 0 16082 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[8]
port 177 nsew signal input
flabel metal2 s 16302 0 16358 400 0 FreeSans 224 90 0 0 mprj_HWDATA_core[9]
port 178 nsew signal input
flabel metal2 s 16118 11600 16174 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[0]
port 179 nsew signal output
flabel metal2 s 18878 11600 18934 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[10]
port 180 nsew signal output
flabel metal2 s 19154 11600 19210 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[11]
port 181 nsew signal output
flabel metal2 s 19430 11600 19486 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[12]
port 182 nsew signal output
flabel metal2 s 19706 11600 19762 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[13]
port 183 nsew signal output
flabel metal2 s 19982 11600 20038 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[14]
port 184 nsew signal output
flabel metal2 s 20258 11600 20314 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[15]
port 185 nsew signal output
flabel metal2 s 20534 11600 20590 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[16]
port 186 nsew signal output
flabel metal2 s 20810 11600 20866 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[17]
port 187 nsew signal output
flabel metal2 s 21086 11600 21142 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[18]
port 188 nsew signal output
flabel metal2 s 21362 11600 21418 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[19]
port 189 nsew signal output
flabel metal2 s 16394 11600 16450 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[1]
port 190 nsew signal output
flabel metal2 s 21638 11600 21694 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[20]
port 191 nsew signal output
flabel metal2 s 21914 11600 21970 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[21]
port 192 nsew signal output
flabel metal2 s 22190 11600 22246 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[22]
port 193 nsew signal output
flabel metal2 s 22466 11600 22522 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[23]
port 194 nsew signal output
flabel metal2 s 22742 11600 22798 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[24]
port 195 nsew signal output
flabel metal2 s 23018 11600 23074 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[25]
port 196 nsew signal output
flabel metal2 s 23294 11600 23350 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[26]
port 197 nsew signal output
flabel metal2 s 23570 11600 23626 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[27]
port 198 nsew signal output
flabel metal2 s 23846 11600 23902 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[28]
port 199 nsew signal output
flabel metal2 s 24122 11600 24178 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[29]
port 200 nsew signal output
flabel metal2 s 16670 11600 16726 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[2]
port 201 nsew signal output
flabel metal2 s 24398 11600 24454 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[30]
port 202 nsew signal output
flabel metal2 s 24674 11600 24730 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[31]
port 203 nsew signal output
flabel metal2 s 16946 11600 17002 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[3]
port 204 nsew signal output
flabel metal2 s 17222 11600 17278 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[4]
port 205 nsew signal output
flabel metal2 s 17498 11600 17554 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[5]
port 206 nsew signal output
flabel metal2 s 17774 11600 17830 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[6]
port 207 nsew signal output
flabel metal2 s 18050 11600 18106 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[7]
port 208 nsew signal output
flabel metal2 s 18326 11600 18382 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[8]
port 209 nsew signal output
flabel metal2 s 18602 11600 18658 12000 0 FreeSans 224 90 0 0 mprj_HWDATA_user[9]
port 210 nsew signal output
flabel metal2 s 3882 0 3938 400 0 FreeSans 224 90 0 0 mprj_HWRITE_core
port 211 nsew signal input
flabel metal2 s 6182 11600 6238 12000 0 FreeSans 224 90 0 0 mprj_HWRITE_user
port 212 nsew signal output
flabel metal2 s 5078 11600 5134 12000 0 FreeSans 224 90 0 0 user_HCLK
port 213 nsew signal output
flabel metal2 s 5354 11600 5410 12000 0 FreeSans 224 90 0 0 user_HRESETn
port 214 nsew signal output
flabel metal2 s 34610 11600 34666 12000 0 FreeSans 224 90 0 0 user_irq[0]
port 215 nsew signal input
flabel metal2 s 37370 11600 37426 12000 0 FreeSans 224 90 0 0 user_irq[10]
port 216 nsew signal input
flabel metal2 s 37646 11600 37702 12000 0 FreeSans 224 90 0 0 user_irq[11]
port 217 nsew signal input
flabel metal2 s 37922 11600 37978 12000 0 FreeSans 224 90 0 0 user_irq[12]
port 218 nsew signal input
flabel metal2 s 38198 11600 38254 12000 0 FreeSans 224 90 0 0 user_irq[13]
port 219 nsew signal input
flabel metal2 s 38474 11600 38530 12000 0 FreeSans 224 90 0 0 user_irq[14]
port 220 nsew signal input
flabel metal2 s 38750 11600 38806 12000 0 FreeSans 224 90 0 0 user_irq[15]
port 221 nsew signal input
flabel metal2 s 34886 11600 34942 12000 0 FreeSans 224 90 0 0 user_irq[1]
port 222 nsew signal input
flabel metal2 s 35162 11600 35218 12000 0 FreeSans 224 90 0 0 user_irq[2]
port 223 nsew signal input
flabel metal2 s 35438 11600 35494 12000 0 FreeSans 224 90 0 0 user_irq[3]
port 224 nsew signal input
flabel metal2 s 35714 11600 35770 12000 0 FreeSans 224 90 0 0 user_irq[4]
port 225 nsew signal input
flabel metal2 s 35990 11600 36046 12000 0 FreeSans 224 90 0 0 user_irq[5]
port 226 nsew signal input
flabel metal2 s 36266 11600 36322 12000 0 FreeSans 224 90 0 0 user_irq[6]
port 227 nsew signal input
flabel metal2 s 36542 11600 36598 12000 0 FreeSans 224 90 0 0 user_irq[7]
port 228 nsew signal input
flabel metal2 s 36818 11600 36874 12000 0 FreeSans 224 90 0 0 user_irq[8]
port 229 nsew signal input
flabel metal2 s 37094 11600 37150 12000 0 FreeSans 224 90 0 0 user_irq[9]
port 230 nsew signal input
flabel metal2 s 37002 0 37058 400 0 FreeSans 224 90 0 0 user_irq_core[0]
port 231 nsew signal output
flabel metal2 s 39762 0 39818 400 0 FreeSans 224 90 0 0 user_irq_core[10]
port 232 nsew signal output
flabel metal2 s 40038 0 40094 400 0 FreeSans 224 90 0 0 user_irq_core[11]
port 233 nsew signal output
flabel metal2 s 40314 0 40370 400 0 FreeSans 224 90 0 0 user_irq_core[12]
port 234 nsew signal output
flabel metal2 s 40590 0 40646 400 0 FreeSans 224 90 0 0 user_irq_core[13]
port 235 nsew signal output
flabel metal2 s 40866 0 40922 400 0 FreeSans 224 90 0 0 user_irq_core[14]
port 236 nsew signal output
flabel metal2 s 41142 0 41198 400 0 FreeSans 224 90 0 0 user_irq_core[15]
port 237 nsew signal output
flabel metal2 s 37278 0 37334 400 0 FreeSans 224 90 0 0 user_irq_core[1]
port 238 nsew signal output
flabel metal2 s 37554 0 37610 400 0 FreeSans 224 90 0 0 user_irq_core[2]
port 239 nsew signal output
flabel metal2 s 37830 0 37886 400 0 FreeSans 224 90 0 0 user_irq_core[3]
port 240 nsew signal output
flabel metal2 s 38106 0 38162 400 0 FreeSans 224 90 0 0 user_irq_core[4]
port 241 nsew signal output
flabel metal2 s 38382 0 38438 400 0 FreeSans 224 90 0 0 user_irq_core[5]
port 242 nsew signal output
flabel metal2 s 38658 0 38714 400 0 FreeSans 224 90 0 0 user_irq_core[6]
port 243 nsew signal output
flabel metal2 s 38934 0 38990 400 0 FreeSans 224 90 0 0 user_irq_core[7]
port 244 nsew signal output
flabel metal2 s 39210 0 39266 400 0 FreeSans 224 90 0 0 user_irq_core[8]
port 245 nsew signal output
flabel metal2 s 39486 0 39542 400 0 FreeSans 224 90 0 0 user_irq_core[9]
port 246 nsew signal output
flabel metal2 s 32586 0 32642 400 0 FreeSans 224 90 0 0 user_irq_ena[0]
port 247 nsew signal input
flabel metal2 s 35346 0 35402 400 0 FreeSans 224 90 0 0 user_irq_ena[10]
port 248 nsew signal input
flabel metal2 s 35622 0 35678 400 0 FreeSans 224 90 0 0 user_irq_ena[11]
port 249 nsew signal input
flabel metal2 s 35898 0 35954 400 0 FreeSans 224 90 0 0 user_irq_ena[12]
port 250 nsew signal input
flabel metal2 s 36174 0 36230 400 0 FreeSans 224 90 0 0 user_irq_ena[13]
port 251 nsew signal input
flabel metal2 s 36450 0 36506 400 0 FreeSans 224 90 0 0 user_irq_ena[14]
port 252 nsew signal input
flabel metal2 s 36726 0 36782 400 0 FreeSans 224 90 0 0 user_irq_ena[15]
port 253 nsew signal input
flabel metal2 s 32862 0 32918 400 0 FreeSans 224 90 0 0 user_irq_ena[1]
port 254 nsew signal input
flabel metal2 s 33138 0 33194 400 0 FreeSans 224 90 0 0 user_irq_ena[2]
port 255 nsew signal input
flabel metal2 s 33414 0 33470 400 0 FreeSans 224 90 0 0 user_irq_ena[3]
port 256 nsew signal input
flabel metal2 s 33690 0 33746 400 0 FreeSans 224 90 0 0 user_irq_ena[4]
port 257 nsew signal input
flabel metal2 s 33966 0 34022 400 0 FreeSans 224 90 0 0 user_irq_ena[5]
port 258 nsew signal input
flabel metal2 s 34242 0 34298 400 0 FreeSans 224 90 0 0 user_irq_ena[6]
port 259 nsew signal input
flabel metal2 s 34518 0 34574 400 0 FreeSans 224 90 0 0 user_irq_ena[7]
port 260 nsew signal input
flabel metal2 s 34794 0 34850 400 0 FreeSans 224 90 0 0 user_irq_ena[8]
port 261 nsew signal input
flabel metal2 s 35070 0 35126 400 0 FreeSans 224 90 0 0 user_irq_ena[9]
port 262 nsew signal input
flabel metal4 s 1300 496 1620 11472 0 FreeSans 1920 90 0 0 vccd0
port 263 nsew power bidirectional
flabel metal4 s 9300 496 9620 11472 0 FreeSans 1920 90 0 0 vccd0
port 263 nsew power bidirectional
flabel metal4 s 17300 496 17620 11472 0 FreeSans 1920 90 0 0 vccd0
port 263 nsew power bidirectional
flabel metal4 s 25300 496 25620 11472 0 FreeSans 1920 90 0 0 vccd0
port 263 nsew power bidirectional
flabel metal4 s 33300 496 33620 11472 0 FreeSans 1920 90 0 0 vccd0
port 263 nsew power bidirectional
flabel metal4 s 41300 496 41620 11472 0 FreeSans 1920 90 0 0 vccd0
port 263 nsew power bidirectional
flabel metal4 s 18580 496 18900 11472 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 26580 496 26900 11472 0 FreeSans 1920 90 0 0 vccd1
port 264 nsew power bidirectional
flabel metal4 s 1940 496 2260 11472 0 FreeSans 1920 90 0 0 vssd0
port 265 nsew ground bidirectional
flabel metal4 s 9940 496 10260 11472 0 FreeSans 1920 90 0 0 vssd0
port 265 nsew ground bidirectional
flabel metal4 s 17940 496 18260 11472 0 FreeSans 1920 90 0 0 vssd0
port 265 nsew ground bidirectional
flabel metal4 s 25940 496 26260 11472 0 FreeSans 1920 90 0 0 vssd0
port 265 nsew ground bidirectional
flabel metal4 s 33940 496 34260 11472 0 FreeSans 1920 90 0 0 vssd0
port 265 nsew ground bidirectional
flabel metal4 s 41940 496 42260 11472 0 FreeSans 1920 90 0 0 vssd0
port 265 nsew ground bidirectional
flabel metal4 s 19220 496 19540 11472 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
flabel metal4 s 27220 496 27540 11472 0 FreeSans 1920 90 0 0 vssd1
port 266 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 44000 12000
<< end >>
