magic
tech sky130A
magscale 1 2
timestamp 1750223503
<< viali >>
rect 4353 13413 4387 13447
rect 5825 13413 5859 13447
rect 10241 13413 10275 13447
rect 12357 13413 12391 13447
rect 3249 13345 3283 13379
rect 17969 13345 18003 13379
rect 3525 13277 3559 13311
rect 3801 13277 3835 13311
rect 4174 13277 4208 13311
rect 5089 13277 5123 13311
rect 5365 13277 5399 13311
rect 5549 13277 5583 13311
rect 6837 13277 6871 13311
rect 10793 13277 10827 13311
rect 11069 13277 11103 13311
rect 11161 13277 11195 13311
rect 11805 13277 11839 13311
rect 12225 13277 12259 13311
rect 14749 13277 14783 13311
rect 15485 13277 15519 13311
rect 16221 13277 16255 13311
rect 16681 13277 16715 13311
rect 17417 13277 17451 13311
rect 18153 13277 18187 13311
rect 19257 13277 19291 13311
rect 21557 13277 21591 13311
rect 2973 13209 3007 13243
rect 3985 13209 4019 13243
rect 4077 13209 4111 13243
rect 6193 13209 6227 13243
rect 7113 13209 7147 13243
rect 10609 13209 10643 13243
rect 11989 13209 12023 13243
rect 12081 13209 12115 13243
rect 20545 13209 20579 13243
rect 1501 13141 1535 13175
rect 3433 13141 3467 13175
rect 4997 13141 5031 13175
rect 5457 13141 5491 13175
rect 5733 13141 5767 13175
rect 8585 13141 8619 13175
rect 10149 13141 10183 13175
rect 10793 13141 10827 13175
rect 11253 13141 11287 13175
rect 14197 13141 14231 13175
rect 14933 13141 14967 13175
rect 15669 13141 15703 13175
rect 17233 13141 17267 13175
rect 18705 13141 18739 13175
rect 19809 13141 19843 13175
rect 6101 12937 6135 12971
rect 13277 12937 13311 12971
rect 14749 12937 14783 12971
rect 15485 12937 15519 12971
rect 16221 12937 16255 12971
rect 2513 12869 2547 12903
rect 7021 12869 7055 12903
rect 9781 12869 9815 12903
rect 16681 12869 16715 12903
rect 17877 12869 17911 12903
rect 18613 12869 18647 12903
rect 18889 12869 18923 12903
rect 4353 12801 4387 12835
rect 6561 12801 6595 12835
rect 6837 12801 6871 12835
rect 7113 12801 7147 12835
rect 7210 12801 7244 12835
rect 11529 12801 11563 12835
rect 13461 12801 13495 12835
rect 14197 12801 14231 12835
rect 14933 12801 14967 12835
rect 15669 12801 15703 12835
rect 17417 12801 17451 12835
rect 19625 12801 19659 12835
rect 19809 12801 19843 12835
rect 2145 12733 2179 12767
rect 2237 12733 2271 12767
rect 4629 12733 4663 12767
rect 7573 12733 7607 12767
rect 7849 12733 7883 12767
rect 9321 12733 9355 12767
rect 9505 12733 9539 12767
rect 11253 12733 11287 12767
rect 11805 12733 11839 12767
rect 14013 12733 14047 12767
rect 20085 12733 20119 12767
rect 21557 12733 21591 12767
rect 22385 12733 22419 12767
rect 1777 12665 1811 12699
rect 7389 12665 7423 12699
rect 1685 12597 1719 12631
rect 3985 12597 4019 12631
rect 6653 12597 6687 12631
rect 21833 12597 21867 12631
rect 1593 12393 1627 12427
rect 3985 12393 4019 12427
rect 4445 12393 4479 12427
rect 12633 12393 12667 12427
rect 13185 12393 13219 12427
rect 16589 12393 16623 12427
rect 17325 12393 17359 12427
rect 8493 12325 8527 12359
rect 1777 12257 1811 12291
rect 6193 12257 6227 12291
rect 10517 12257 10551 12291
rect 10793 12257 10827 12291
rect 15853 12257 15887 12291
rect 17785 12257 17819 12291
rect 20085 12257 20119 12291
rect 20545 12257 20579 12291
rect 22293 12257 22327 12291
rect 1685 12189 1719 12223
rect 4261 12189 4295 12223
rect 6285 12189 6319 12223
rect 10885 12189 10919 12223
rect 13737 12189 13771 12223
rect 14105 12189 14139 12223
rect 16037 12189 16071 12223
rect 16773 12189 16807 12223
rect 18337 12189 18371 12223
rect 18429 12189 18463 12223
rect 19257 12189 19291 12223
rect 20269 12189 20303 12223
rect 2053 12121 2087 12155
rect 3801 12121 3835 12155
rect 5917 12121 5951 12155
rect 6561 12121 6595 12155
rect 8217 12121 8251 12155
rect 11161 12121 11195 12155
rect 14381 12121 14415 12155
rect 3525 12053 3559 12087
rect 3985 12053 4019 12087
rect 8033 12053 8067 12087
rect 8677 12053 8711 12087
rect 9045 12053 9079 12087
rect 18981 12053 19015 12087
rect 2881 11849 2915 11883
rect 5089 11849 5123 11883
rect 5365 11849 5399 11883
rect 11253 11849 11287 11883
rect 15669 11849 15703 11883
rect 18705 11849 18739 11883
rect 19441 11849 19475 11883
rect 20913 11849 20947 11883
rect 3617 11781 3651 11815
rect 5917 11781 5951 11815
rect 7205 11781 7239 11815
rect 9873 11781 9907 11815
rect 1685 11713 1719 11747
rect 2881 11713 2915 11747
rect 3157 11713 3191 11747
rect 3341 11713 3375 11747
rect 5273 11713 5307 11747
rect 5773 11713 5807 11747
rect 6009 11713 6043 11747
rect 6193 11713 6227 11747
rect 6469 11713 6503 11747
rect 6745 11713 6779 11747
rect 6929 11713 6963 11747
rect 7113 11713 7147 11747
rect 7349 11713 7383 11747
rect 7665 11713 7699 11747
rect 9689 11713 9723 11747
rect 9965 11713 9999 11747
rect 10109 11713 10143 11747
rect 10649 11713 10683 11747
rect 10793 11713 10827 11747
rect 10885 11713 10919 11747
rect 11069 11713 11103 11747
rect 11161 11713 11195 11747
rect 11621 11713 11655 11747
rect 11897 11713 11931 11747
rect 13829 11713 13863 11747
rect 14565 11713 14599 11747
rect 14841 11713 14875 11747
rect 15761 11713 15795 11747
rect 16681 11713 16715 11747
rect 17417 11713 17451 11747
rect 18153 11713 18187 11747
rect 18889 11713 18923 11747
rect 21005 11713 21039 11747
rect 2697 11645 2731 11679
rect 7941 11645 7975 11679
rect 9413 11645 9447 11679
rect 12725 11645 12759 11679
rect 14381 11645 14415 11679
rect 17233 11645 17267 11679
rect 17969 11645 18003 11679
rect 5641 11577 5675 11611
rect 6469 11577 6503 11611
rect 7481 11577 7515 11611
rect 10241 11577 10275 11611
rect 11621 11577 11655 11611
rect 13001 11577 13035 11611
rect 14657 11577 14691 11611
rect 10517 11509 10551 11543
rect 13185 11509 13219 11543
rect 15393 11509 15427 11543
rect 1869 11305 1903 11339
rect 6745 11305 6779 11339
rect 7192 11305 7226 11339
rect 9413 11305 9447 11339
rect 13001 11305 13035 11339
rect 13737 11305 13771 11339
rect 16681 11305 16715 11339
rect 3341 11169 3375 11203
rect 3893 11169 3927 11203
rect 4353 11169 4387 11203
rect 4997 11169 5031 11203
rect 5273 11169 5307 11203
rect 6929 11169 6963 11203
rect 10885 11169 10919 11203
rect 11161 11169 11195 11203
rect 11253 11169 11287 11203
rect 11529 11169 11563 11203
rect 14289 11169 14323 11203
rect 3617 11101 3651 11135
rect 4077 11101 4111 11135
rect 4445 11101 4479 11135
rect 4629 11101 4663 11135
rect 4905 11101 4939 11135
rect 8953 11101 8987 11135
rect 13185 11101 13219 11135
rect 13461 11101 13495 11135
rect 13558 11101 13592 11135
rect 16037 11101 16071 11135
rect 16129 11101 16163 11135
rect 4537 11033 4571 11067
rect 13369 11033 13403 11067
rect 15761 11033 15795 11067
rect 8677 10965 8711 10999
rect 9045 10965 9079 10999
rect 3709 10761 3743 10795
rect 5917 10761 5951 10795
rect 14841 10761 14875 10795
rect 16773 10761 16807 10795
rect 1777 10693 1811 10727
rect 2237 10693 2271 10727
rect 4445 10693 4479 10727
rect 9965 10693 9999 10727
rect 10701 10693 10735 10727
rect 13369 10693 13403 10727
rect 15485 10693 15519 10727
rect 1685 10625 1719 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 9597 10625 9631 10659
rect 9781 10625 9815 10659
rect 10054 10625 10088 10659
rect 10201 10625 10235 10659
rect 10563 10625 10597 10659
rect 10793 10625 10827 10659
rect 10937 10625 10971 10659
rect 11529 10625 11563 10659
rect 11713 10625 11747 10659
rect 11805 10625 11839 10659
rect 11949 10625 11983 10659
rect 15296 10625 15330 10659
rect 15393 10625 15427 10659
rect 15669 10625 15703 10659
rect 16681 10625 16715 10659
rect 18797 10625 18831 10659
rect 1961 10557 1995 10591
rect 4169 10557 4203 10591
rect 6377 10557 6411 10591
rect 7849 10557 7883 10591
rect 9321 10557 9355 10591
rect 13093 10557 13127 10591
rect 15761 10557 15795 10591
rect 17049 10557 17083 10591
rect 18521 10557 18555 10591
rect 11069 10489 11103 10523
rect 16037 10489 16071 10523
rect 10333 10421 10367 10455
rect 12081 10421 12115 10455
rect 15117 10421 15151 10455
rect 16221 10421 16255 10455
rect 1869 10217 1903 10251
rect 3065 10217 3099 10251
rect 4353 10217 4387 10251
rect 7297 10217 7331 10251
rect 13277 10217 13311 10251
rect 16037 10217 16071 10251
rect 17969 10217 18003 10251
rect 5365 10149 5399 10183
rect 8401 10149 8435 10183
rect 5549 10081 5583 10115
rect 5825 10081 5859 10115
rect 9781 10081 9815 10115
rect 11529 10081 11563 10115
rect 11805 10081 11839 10115
rect 16497 10081 16531 10115
rect 2048 10013 2082 10047
rect 2145 10013 2179 10047
rect 2421 10013 2455 10047
rect 2513 10013 2547 10047
rect 2933 10013 2967 10047
rect 3801 10013 3835 10047
rect 4174 10013 4208 10047
rect 4813 10013 4847 10047
rect 5233 10013 5267 10047
rect 7573 10013 7607 10047
rect 7665 10013 7699 10047
rect 7849 10013 7883 10047
rect 8125 10013 8159 10047
rect 8222 10013 8256 10047
rect 10517 10013 10551 10047
rect 10890 10013 10924 10047
rect 13737 10013 13771 10047
rect 13921 10013 13955 10047
rect 14289 10013 14323 10047
rect 16221 10013 16255 10047
rect 2237 9945 2271 9979
rect 2697 9945 2731 9979
rect 2789 9945 2823 9979
rect 3985 9945 4019 9979
rect 4077 9945 4111 9979
rect 4997 9945 5031 9979
rect 5089 9945 5123 9979
rect 8033 9945 8067 9979
rect 8953 9945 8987 9979
rect 10701 9945 10735 9979
rect 10793 9945 10827 9979
rect 13553 9945 13587 9979
rect 14565 9945 14599 9979
rect 11086 9877 11120 9911
rect 1961 9605 1995 9639
rect 5733 9605 5767 9639
rect 8769 9605 8803 9639
rect 13461 9605 13495 9639
rect 15485 9605 15519 9639
rect 2053 9537 2087 9571
rect 4169 9537 4203 9571
rect 4445 9537 4479 9571
rect 5549 9537 5583 9571
rect 5825 9537 5859 9571
rect 5969 9537 6003 9571
rect 8493 9537 8527 9571
rect 10425 9537 10459 9571
rect 11529 9537 11563 9571
rect 11713 9537 11747 9571
rect 11805 9537 11839 9571
rect 11949 9537 11983 9571
rect 12265 9537 12299 9571
rect 12449 9537 12483 9571
rect 13185 9537 13219 9571
rect 15117 9537 15151 9571
rect 15393 9537 15427 9571
rect 16681 9537 16715 9571
rect 16865 9537 16899 9571
rect 2329 9469 2363 9503
rect 6377 9469 6411 9503
rect 6653 9469 6687 9503
rect 8125 9469 8159 9503
rect 10241 9469 10275 9503
rect 11161 9469 11195 9503
rect 12817 9469 12851 9503
rect 14933 9469 14967 9503
rect 16313 9469 16347 9503
rect 19165 9469 19199 9503
rect 19441 9469 19475 9503
rect 1593 9401 1627 9435
rect 4353 9401 4387 9435
rect 6101 9401 6135 9435
rect 12725 9401 12759 9435
rect 15301 9401 15335 9435
rect 15945 9401 15979 9435
rect 16957 9401 16991 9435
rect 1501 9333 1535 9367
rect 3801 9333 3835 9367
rect 4077 9333 4111 9367
rect 12081 9333 12115 9367
rect 15853 9333 15887 9367
rect 17693 9333 17727 9367
rect 2034 9129 2068 9163
rect 5733 9129 5767 9163
rect 17693 9129 17727 9163
rect 6561 9061 6595 9095
rect 13093 9061 13127 9095
rect 1777 8993 1811 9027
rect 3985 8993 4019 9027
rect 6929 8993 6963 9027
rect 8677 8993 8711 9027
rect 9229 8993 9263 9027
rect 11345 8993 11379 9027
rect 14657 8993 14691 9027
rect 6561 8925 6595 8959
rect 6837 8925 6871 8959
rect 8953 8925 8987 8959
rect 11069 8925 11103 8959
rect 11253 8925 11287 8959
rect 14933 8925 14967 8959
rect 15393 8925 15427 8959
rect 15485 8925 15519 8959
rect 15669 8925 15703 8959
rect 17601 8925 17635 8959
rect 4261 8857 4295 8891
rect 7205 8857 7239 8891
rect 11621 8857 11655 8891
rect 15945 8857 15979 8891
rect 3525 8789 3559 8823
rect 10701 8789 10735 8823
rect 11161 8789 11195 8823
rect 14105 8789 14139 8823
rect 17417 8789 17451 8823
rect 2605 8585 2639 8619
rect 5457 8585 5491 8619
rect 11989 8585 12023 8619
rect 14749 8585 14783 8619
rect 18429 8585 18463 8619
rect 3157 8517 3191 8551
rect 3985 8517 4019 8551
rect 11529 8517 11563 8551
rect 12173 8517 12207 8551
rect 12357 8517 12391 8551
rect 13277 8517 13311 8551
rect 16221 8517 16255 8551
rect 16313 8517 16347 8551
rect 2001 8449 2035 8483
rect 2145 8449 2179 8483
rect 2237 8449 2271 8483
rect 2421 8449 2455 8483
rect 2513 8449 2547 8483
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3249 8449 3283 8483
rect 3393 8449 3427 8483
rect 3709 8449 3743 8483
rect 9045 8449 9079 8483
rect 9137 8449 9171 8483
rect 9505 8449 9539 8483
rect 12725 8449 12759 8483
rect 13001 8449 13035 8483
rect 16124 8449 16158 8483
rect 16497 8449 16531 8483
rect 16681 8449 16715 8483
rect 6377 8381 6411 8415
rect 6653 8381 6687 8415
rect 8309 8381 8343 8415
rect 9781 8381 9815 8415
rect 16957 8381 16991 8415
rect 1869 8313 1903 8347
rect 3525 8313 3559 8347
rect 8585 8313 8619 8347
rect 11253 8313 11287 8347
rect 11805 8313 11839 8347
rect 12541 8313 12575 8347
rect 15945 8313 15979 8347
rect 8125 8245 8159 8279
rect 8769 8245 8803 8279
rect 12357 8245 12391 8279
rect 12817 8245 12851 8279
rect 3525 8041 3559 8075
rect 6193 8041 6227 8075
rect 8217 8041 8251 8075
rect 11621 8041 11655 8075
rect 16313 8041 16347 8075
rect 4077 7973 4111 8007
rect 3801 7905 3835 7939
rect 6745 7905 6779 7939
rect 13093 7905 13127 7939
rect 13369 7905 13403 7939
rect 14565 7905 14599 7939
rect 1501 7837 1535 7871
rect 1593 7837 1627 7871
rect 1777 7837 1811 7871
rect 4445 7837 4479 7871
rect 6469 7837 6503 7871
rect 11437 7837 11471 7871
rect 13461 7837 13495 7871
rect 13737 7837 13771 7871
rect 14289 7837 14323 7871
rect 2053 7769 2087 7803
rect 4721 7769 4755 7803
rect 11161 7769 11195 7803
rect 14841 7769 14875 7803
rect 4261 7701 4295 7735
rect 9689 7701 9723 7735
rect 13737 7701 13771 7735
rect 14197 7701 14231 7735
rect 3157 7497 3191 7531
rect 3433 7497 3467 7531
rect 5365 7497 5399 7531
rect 6561 7497 6595 7531
rect 6837 7497 6871 7531
rect 9965 7497 9999 7531
rect 10701 7497 10735 7531
rect 3893 7429 3927 7463
rect 7757 7429 7791 7463
rect 8493 7429 8527 7463
rect 13737 7429 13771 7463
rect 15577 7429 15611 7463
rect 1409 7361 1443 7395
rect 3341 7361 3375 7395
rect 3617 7361 3651 7395
rect 6653 7361 6687 7395
rect 6929 7361 6963 7395
rect 7021 7361 7055 7395
rect 7660 7361 7694 7395
rect 7849 7361 7883 7395
rect 8033 7361 8067 7395
rect 10149 7361 10183 7395
rect 10333 7361 10367 7395
rect 10609 7361 10643 7395
rect 11069 7361 11103 7395
rect 15393 7361 15427 7395
rect 15669 7361 15703 7395
rect 15807 7361 15841 7395
rect 16129 7361 16163 7395
rect 1685 7293 1719 7327
rect 8217 7293 8251 7327
rect 13369 7293 13403 7327
rect 13461 7293 13495 7327
rect 10425 7225 10459 7259
rect 13001 7225 13035 7259
rect 15945 7225 15979 7259
rect 7481 7157 7515 7191
rect 11161 7157 11195 7191
rect 12909 7157 12943 7191
rect 15209 7157 15243 7191
rect 16221 7157 16255 7191
rect 2040 6953 2074 6987
rect 9505 6953 9539 6987
rect 10412 6953 10446 6987
rect 12344 6953 12378 6987
rect 16294 6953 16328 6987
rect 3525 6885 3559 6919
rect 7113 6885 7147 6919
rect 1777 6817 1811 6851
rect 5365 6817 5399 6851
rect 10149 6817 10183 6851
rect 12081 6817 12115 6851
rect 14105 6817 14139 6851
rect 15853 6817 15887 6851
rect 16037 6817 16071 6851
rect 17785 6817 17819 6851
rect 4169 6749 4203 6783
rect 4542 6749 4576 6783
rect 4738 6749 4772 6783
rect 5089 6749 5123 6783
rect 7665 6749 7699 6783
rect 8125 6749 8159 6783
rect 9229 6749 9263 6783
rect 9321 6749 9355 6783
rect 9684 6749 9718 6783
rect 10057 6749 10091 6783
rect 4353 6681 4387 6715
rect 4445 6681 4479 6715
rect 5641 6681 5675 6715
rect 9781 6681 9815 6715
rect 9873 6681 9907 6715
rect 14381 6681 14415 6715
rect 4997 6613 5031 6647
rect 7297 6613 7331 6647
rect 11897 6613 11931 6647
rect 13829 6613 13863 6647
rect 1685 6409 1719 6443
rect 5549 6409 5583 6443
rect 6837 6409 6871 6443
rect 9229 6409 9263 6443
rect 11161 6409 11195 6443
rect 4077 6341 4111 6375
rect 5825 6341 5859 6375
rect 7757 6341 7791 6375
rect 1593 6273 1627 6307
rect 1777 6273 1811 6307
rect 2140 6273 2174 6307
rect 2237 6273 2271 6307
rect 2329 6273 2363 6307
rect 2513 6273 2547 6307
rect 2789 6273 2823 6307
rect 2881 6273 2915 6307
rect 3065 6273 3099 6307
rect 3157 6273 3191 6307
rect 3301 6273 3335 6307
rect 6009 6273 6043 6307
rect 6193 6273 6227 6307
rect 6837 6273 6871 6307
rect 7205 6273 7239 6307
rect 9413 6273 9447 6307
rect 11621 6273 11655 6307
rect 3801 6205 3835 6239
rect 6653 6205 6687 6239
rect 7481 6205 7515 6239
rect 9689 6205 9723 6239
rect 11897 6205 11931 6239
rect 1961 6137 1995 6171
rect 3433 6137 3467 6171
rect 2697 6069 2731 6103
rect 13369 6069 13403 6103
rect 4537 5865 4571 5899
rect 6837 5865 6871 5899
rect 7665 5865 7699 5899
rect 9597 5865 9631 5899
rect 12173 5865 12207 5899
rect 14105 5865 14139 5899
rect 6653 5797 6687 5831
rect 8493 5797 8527 5831
rect 9689 5797 9723 5831
rect 1777 5729 1811 5763
rect 3525 5729 3559 5763
rect 5549 5729 5583 5763
rect 10057 5729 10091 5763
rect 10425 5729 10459 5763
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 4358 5661 4392 5695
rect 6193 5661 6227 5695
rect 6469 5661 6503 5695
rect 7113 5661 7147 5695
rect 7297 5661 7331 5695
rect 7533 5661 7567 5695
rect 7849 5661 7883 5695
rect 8953 5661 8987 5695
rect 12449 5661 12483 5695
rect 12633 5661 12667 5695
rect 13001 5661 13035 5695
rect 14749 5661 14783 5695
rect 2053 5593 2087 5627
rect 4169 5593 4203 5627
rect 4721 5593 4755 5627
rect 7021 5593 7055 5627
rect 7389 5593 7423 5627
rect 8217 5593 8251 5627
rect 10701 5593 10735 5627
rect 6193 5525 6227 5559
rect 6837 5525 6871 5559
rect 7941 5525 7975 5559
rect 8677 5525 8711 5559
rect 9045 5525 9079 5559
rect 12633 5525 12667 5559
rect 13093 5525 13127 5559
rect 1501 5321 1535 5355
rect 6101 5321 6135 5355
rect 8861 5321 8895 5355
rect 10977 5321 11011 5355
rect 15117 5321 15151 5355
rect 3893 5253 3927 5287
rect 4629 5253 4663 5287
rect 12081 5253 12115 5287
rect 12725 5253 12759 5287
rect 3249 5185 3283 5219
rect 3341 5185 3375 5219
rect 3617 5185 3651 5219
rect 3801 5185 3835 5219
rect 3990 5185 4024 5219
rect 7113 5185 7147 5219
rect 9229 5185 9263 5219
rect 12357 5185 12391 5219
rect 12449 5185 12483 5219
rect 12633 5185 12667 5219
rect 12822 5185 12856 5219
rect 13369 5185 13403 5219
rect 2973 5117 3007 5151
rect 4353 5117 4387 5151
rect 6377 5117 6411 5151
rect 7389 5117 7423 5151
rect 9505 5117 9539 5151
rect 13645 5117 13679 5151
rect 4169 5049 4203 5083
rect 6653 5049 6687 5083
rect 11713 5049 11747 5083
rect 3433 4981 3467 5015
rect 6837 4981 6871 5015
rect 11621 4981 11655 5015
rect 12265 4981 12299 5015
rect 13001 4981 13035 5015
rect 5549 4777 5583 4811
rect 8125 4777 8159 4811
rect 12344 4777 12378 4811
rect 13829 4777 13863 4811
rect 3525 4709 3559 4743
rect 7757 4709 7791 4743
rect 9137 4709 9171 4743
rect 1777 4641 1811 4675
rect 3801 4641 3835 4675
rect 4077 4641 4111 4675
rect 6009 4641 6043 4675
rect 6285 4641 6319 4675
rect 10425 4641 10459 4675
rect 12081 4641 12115 4675
rect 5917 4573 5951 4607
rect 8263 4573 8297 4607
rect 8401 4573 8435 4607
rect 8677 4573 8711 4607
rect 9505 4573 9539 4607
rect 9781 4573 9815 4607
rect 10149 4573 10183 4607
rect 14289 4573 14323 4607
rect 2053 4505 2087 4539
rect 8493 4505 8527 4539
rect 5825 4437 5859 4471
rect 9045 4437 9079 4471
rect 9689 4437 9723 4471
rect 11897 4437 11931 4471
rect 14197 4437 14231 4471
rect 1593 4233 1627 4267
rect 5917 4233 5951 4267
rect 10149 4233 10183 4267
rect 13553 4233 13587 4267
rect 4169 4165 4203 4199
rect 12081 4165 12115 4199
rect 2053 4097 2087 4131
rect 3060 4097 3094 4131
rect 3157 4097 3191 4131
rect 3249 4097 3283 4131
rect 3433 4097 3467 4131
rect 3525 4097 3559 4131
rect 3893 4097 3927 4131
rect 5825 4097 5859 4131
rect 6009 4097 6043 4131
rect 8401 4097 8435 4131
rect 10333 4097 10367 4131
rect 11805 4097 11839 4131
rect 13921 4097 13955 4131
rect 2697 4029 2731 4063
rect 6469 4029 6503 4063
rect 6745 4029 6779 4063
rect 8677 4029 8711 4063
rect 14933 4029 14967 4063
rect 1777 3961 1811 3995
rect 2237 3961 2271 3995
rect 2421 3961 2455 3995
rect 2881 3961 2915 3995
rect 3617 3893 3651 3927
rect 5641 3893 5675 3927
rect 8217 3893 8251 3927
rect 10425 3893 10459 3927
rect 3893 3689 3927 3723
rect 11253 3689 11287 3723
rect 4813 3621 4847 3655
rect 11621 3621 11655 3655
rect 1593 3553 1627 3587
rect 1777 3553 1811 3587
rect 3525 3553 3559 3587
rect 4997 3553 5031 3587
rect 6745 3553 6779 3587
rect 6929 3553 6963 3587
rect 8677 3553 8711 3587
rect 9781 3553 9815 3587
rect 12081 3553 12115 3587
rect 14105 3553 14139 3587
rect 1685 3485 1719 3519
rect 4025 3485 4059 3519
rect 4169 3485 4203 3519
rect 4445 3485 4479 3519
rect 4537 3485 4571 3519
rect 4813 3485 4847 3519
rect 8953 3485 8987 3519
rect 9137 3485 9171 3519
rect 9505 3485 9539 3519
rect 2053 3417 2087 3451
rect 4261 3417 4295 3451
rect 5273 3417 5307 3451
rect 7205 3417 7239 3451
rect 11989 3417 12023 3451
rect 12357 3417 12391 3451
rect 14381 3417 14415 3451
rect 9045 3349 9079 3383
rect 11529 3349 11563 3383
rect 13829 3349 13863 3383
rect 15853 3349 15887 3383
rect 6101 3145 6135 3179
rect 8217 3145 8251 3179
rect 6745 3077 6779 3111
rect 15025 3077 15059 3111
rect 3704 3009 3738 3043
rect 3801 3009 3835 3043
rect 3893 3009 3927 3043
rect 4077 3009 4111 3043
rect 10241 3009 10275 3043
rect 10333 3009 10367 3043
rect 11069 3009 11103 3043
rect 11345 3009 11379 3043
rect 11621 3009 11655 3043
rect 14789 3009 14823 3043
rect 14933 3009 14967 3043
rect 15209 3009 15243 3043
rect 1593 2941 1627 2975
rect 3065 2941 3099 2975
rect 3341 2941 3375 2975
rect 4353 2941 4387 2975
rect 4629 2941 4663 2975
rect 6469 2941 6503 2975
rect 9965 2941 9999 2975
rect 10609 2941 10643 2975
rect 11713 2941 11747 2975
rect 11897 2941 11931 2975
rect 12173 2941 12207 2975
rect 14381 2941 14415 2975
rect 11069 2873 11103 2907
rect 14657 2873 14691 2907
rect 3525 2805 3559 2839
rect 8493 2805 8527 2839
rect 10425 2805 10459 2839
rect 13645 2805 13679 2839
rect 13829 2805 13863 2839
rect 7192 2601 7226 2635
rect 9597 2601 9631 2635
rect 12449 2601 12483 2635
rect 13645 2601 13679 2635
rect 10057 2533 10091 2567
rect 10241 2533 10275 2567
rect 1777 2465 1811 2499
rect 3893 2465 3927 2499
rect 6929 2465 6963 2499
rect 10977 2465 11011 2499
rect 14565 2465 14599 2499
rect 1501 2397 1535 2431
rect 5917 2397 5951 2431
rect 9045 2397 9079 2431
rect 9229 2397 9263 2431
rect 9418 2397 9452 2431
rect 9781 2397 9815 2431
rect 10609 2397 10643 2431
rect 10701 2397 10735 2431
rect 13369 2397 13403 2431
rect 13829 2397 13863 2431
rect 14105 2397 14139 2431
rect 21097 2397 21131 2431
rect 2053 2329 2087 2363
rect 4169 2329 4203 2363
rect 6745 2329 6779 2363
rect 9321 2329 9355 2363
rect 12633 2329 12667 2363
rect 22293 2329 22327 2363
rect 1593 2261 1627 2295
rect 3525 2261 3559 2295
rect 5641 2261 5675 2295
rect 8677 2261 8711 2295
rect 10425 2261 10459 2295
rect 1593 2057 1627 2091
rect 3893 2057 3927 2091
rect 4169 2057 4203 2091
rect 9321 2057 9355 2091
rect 6561 1989 6595 2023
rect 11805 1989 11839 2023
rect 11989 1989 12023 2023
rect 2053 1921 2087 1955
rect 2145 1921 2179 1955
rect 4077 1921 4111 1955
rect 6377 1921 6411 1955
rect 6653 1921 6687 1955
rect 6750 1921 6784 1955
rect 7297 1921 7331 1955
rect 11529 1921 11563 1955
rect 13921 1921 13955 1955
rect 14933 1921 14967 1955
rect 16773 1921 16807 1955
rect 18613 1921 18647 1955
rect 20269 1921 20303 1955
rect 22109 1921 22143 1955
rect 2421 1853 2455 1887
rect 4353 1853 4387 1887
rect 4629 1853 4663 1887
rect 6101 1853 6135 1887
rect 7389 1853 7423 1887
rect 7573 1853 7607 1887
rect 7849 1853 7883 1887
rect 9505 1853 9539 1887
rect 9781 1853 9815 1887
rect 12173 1853 12207 1887
rect 13645 1853 13679 1887
rect 14013 1853 14047 1887
rect 14565 1853 14599 1887
rect 15669 1853 15703 1887
rect 17509 1853 17543 1887
rect 19349 1853 19383 1887
rect 21189 1853 21223 1887
rect 1777 1785 1811 1819
rect 6929 1785 6963 1819
rect 11253 1785 11287 1819
rect 11805 1717 11839 1751
rect 1501 1513 1535 1547
rect 3893 1513 3927 1547
rect 5383 1513 5417 1547
rect 6929 1513 6963 1547
rect 11081 1513 11115 1547
rect 2973 1377 3007 1411
rect 8677 1377 8711 1411
rect 9597 1377 9631 1411
rect 11529 1377 11563 1411
rect 11805 1377 11839 1411
rect 3249 1309 3283 1343
rect 3617 1309 3651 1343
rect 5641 1309 5675 1343
rect 5733 1309 5767 1343
rect 5917 1309 5951 1343
rect 6469 1309 6503 1343
rect 6653 1309 6687 1343
rect 9229 1309 9263 1343
rect 9321 1309 9355 1343
rect 11345 1309 11379 1343
rect 14105 1309 14139 1343
rect 14657 1309 14691 1343
rect 3525 1241 3559 1275
rect 6377 1241 6411 1275
rect 8401 1241 8435 1275
rect 9045 1241 9079 1275
rect 5825 1173 5859 1207
rect 13277 1173 13311 1207
<< metal1 >>
rect 1104 13626 22816 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 20214 13626
rect 20266 13574 20278 13626
rect 20330 13574 20342 13626
rect 20394 13574 20406 13626
rect 20458 13574 20470 13626
rect 20522 13574 22816 13626
rect 1104 13552 22816 13574
rect 4341 13447 4399 13453
rect 4341 13413 4353 13447
rect 4387 13413 4399 13447
rect 4341 13407 4399 13413
rect 3237 13379 3295 13385
rect 3237 13345 3249 13379
rect 3283 13376 3295 13379
rect 3283 13348 4108 13376
rect 3283 13345 3295 13348
rect 3237 13339 3295 13345
rect 3513 13311 3571 13317
rect 3513 13277 3525 13311
rect 3559 13277 3571 13311
rect 3513 13271 3571 13277
rect 2530 13212 2917 13240
rect 1486 13132 1492 13184
rect 1544 13132 1550 13184
rect 2889 13172 2917 13212
rect 2958 13200 2964 13252
rect 3016 13200 3022 13252
rect 3528 13240 3556 13271
rect 3694 13268 3700 13320
rect 3752 13308 3758 13320
rect 3789 13311 3847 13317
rect 3789 13308 3801 13311
rect 3752 13280 3801 13308
rect 3752 13268 3758 13280
rect 3789 13277 3801 13280
rect 3835 13277 3847 13311
rect 3789 13271 3847 13277
rect 3878 13240 3884 13252
rect 3528 13212 3884 13240
rect 3878 13200 3884 13212
rect 3936 13240 3942 13252
rect 4080 13249 4108 13348
rect 4154 13268 4160 13320
rect 4212 13317 4218 13320
rect 4212 13308 4220 13317
rect 4356 13308 4384 13407
rect 5534 13404 5540 13456
rect 5592 13444 5598 13456
rect 5813 13447 5871 13453
rect 5813 13444 5825 13447
rect 5592 13416 5825 13444
rect 5592 13404 5598 13416
rect 5813 13413 5825 13416
rect 5859 13413 5871 13447
rect 5813 13407 5871 13413
rect 10226 13404 10232 13456
rect 10284 13404 10290 13456
rect 12345 13447 12403 13453
rect 12345 13413 12357 13447
rect 12391 13444 12403 13447
rect 12391 13416 19288 13444
rect 12391 13413 12403 13416
rect 12345 13407 12403 13413
rect 6178 13376 6184 13388
rect 5092 13348 6184 13376
rect 5092 13317 5120 13348
rect 6178 13336 6184 13348
rect 6236 13336 6242 13388
rect 17957 13379 18015 13385
rect 11072 13348 12296 13376
rect 5077 13311 5135 13317
rect 5077 13308 5089 13311
rect 4212 13280 4257 13308
rect 4356 13280 5089 13308
rect 4212 13271 4220 13280
rect 5077 13277 5089 13280
rect 5123 13277 5135 13311
rect 5077 13271 5135 13277
rect 5353 13311 5411 13317
rect 5353 13277 5365 13311
rect 5399 13277 5411 13311
rect 5353 13271 5411 13277
rect 4212 13268 4218 13271
rect 3973 13243 4031 13249
rect 3973 13240 3985 13243
rect 3936 13212 3985 13240
rect 3936 13200 3942 13212
rect 3973 13209 3985 13212
rect 4019 13209 4031 13243
rect 3973 13203 4031 13209
rect 4065 13243 4123 13249
rect 4065 13209 4077 13243
rect 4111 13209 4123 13243
rect 5368 13240 5396 13271
rect 5534 13268 5540 13320
rect 5592 13268 5598 13320
rect 5644 13280 6684 13308
rect 5644 13240 5672 13280
rect 5368 13212 5672 13240
rect 4065 13203 4123 13209
rect 3142 13172 3148 13184
rect 2889 13144 3148 13172
rect 3142 13132 3148 13144
rect 3200 13132 3206 13184
rect 3326 13132 3332 13184
rect 3384 13172 3390 13184
rect 3421 13175 3479 13181
rect 3421 13172 3433 13175
rect 3384 13144 3433 13172
rect 3384 13132 3390 13144
rect 3421 13141 3433 13144
rect 3467 13141 3479 13175
rect 3421 13135 3479 13141
rect 3786 13132 3792 13184
rect 3844 13172 3850 13184
rect 4080 13172 4108 13203
rect 6086 13200 6092 13252
rect 6144 13240 6150 13252
rect 6181 13243 6239 13249
rect 6181 13240 6193 13243
rect 6144 13212 6193 13240
rect 6144 13200 6150 13212
rect 6181 13209 6193 13212
rect 6227 13209 6239 13243
rect 6656 13240 6684 13280
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6788 13280 6837 13308
rect 6788 13268 6794 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 10226 13268 10232 13320
rect 10284 13308 10290 13320
rect 11072 13317 11100 13348
rect 10781 13311 10839 13317
rect 10781 13308 10793 13311
rect 10284 13280 10793 13308
rect 10284 13268 10290 13280
rect 10781 13277 10793 13280
rect 10827 13277 10839 13311
rect 10781 13271 10839 13277
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 11146 13268 11152 13320
rect 11204 13308 11210 13320
rect 11698 13308 11704 13320
rect 11204 13280 11704 13308
rect 11204 13268 11210 13280
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 12268 13317 12296 13348
rect 17957 13345 17969 13379
rect 18003 13376 18015 13379
rect 18003 13348 18184 13376
rect 18003 13345 18015 13348
rect 17957 13339 18015 13345
rect 11793 13311 11851 13317
rect 11793 13277 11805 13311
rect 11839 13302 11851 13311
rect 12213 13311 12296 13317
rect 12213 13308 12225 13311
rect 11839 13277 11856 13302
rect 12163 13280 12225 13308
rect 11793 13271 11856 13277
rect 12213 13277 12225 13280
rect 12259 13308 12296 13311
rect 13262 13308 13268 13320
rect 12259 13280 13268 13308
rect 12259 13277 12271 13280
rect 12213 13271 12271 13277
rect 7006 13240 7012 13252
rect 6656 13212 7012 13240
rect 6181 13203 6239 13209
rect 7006 13200 7012 13212
rect 7064 13200 7070 13252
rect 7101 13243 7159 13249
rect 7101 13209 7113 13243
rect 7147 13209 7159 13243
rect 7101 13203 7159 13209
rect 3844 13144 4108 13172
rect 3844 13132 3850 13144
rect 4338 13132 4344 13184
rect 4396 13172 4402 13184
rect 4985 13175 5043 13181
rect 4985 13172 4997 13175
rect 4396 13144 4997 13172
rect 4396 13132 4402 13144
rect 4985 13141 4997 13144
rect 5031 13141 5043 13175
rect 4985 13135 5043 13141
rect 5445 13175 5503 13181
rect 5445 13141 5457 13175
rect 5491 13172 5503 13175
rect 5626 13172 5632 13184
rect 5491 13144 5632 13172
rect 5491 13141 5503 13144
rect 5445 13135 5503 13141
rect 5626 13132 5632 13144
rect 5684 13132 5690 13184
rect 5721 13175 5779 13181
rect 5721 13141 5733 13175
rect 5767 13172 5779 13175
rect 7116 13172 7144 13203
rect 7558 13200 7564 13252
rect 7616 13200 7622 13252
rect 10597 13243 10655 13249
rect 10597 13209 10609 13243
rect 10643 13240 10655 13243
rect 10686 13240 10692 13252
rect 10643 13212 10692 13240
rect 10643 13209 10655 13212
rect 10597 13203 10655 13209
rect 10686 13200 10692 13212
rect 10744 13240 10750 13252
rect 11828 13240 11856 13271
rect 13262 13268 13268 13280
rect 13320 13268 13326 13320
rect 14734 13268 14740 13320
rect 14792 13268 14798 13320
rect 15470 13268 15476 13320
rect 15528 13268 15534 13320
rect 16114 13268 16120 13320
rect 16172 13308 16178 13320
rect 16209 13311 16267 13317
rect 16209 13308 16221 13311
rect 16172 13280 16221 13308
rect 16172 13268 16178 13280
rect 16209 13277 16221 13280
rect 16255 13277 16267 13311
rect 16209 13271 16267 13277
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 16669 13311 16727 13317
rect 16669 13308 16681 13311
rect 16632 13280 16681 13308
rect 16632 13268 16638 13280
rect 16669 13277 16681 13280
rect 16715 13277 16727 13311
rect 16669 13271 16727 13277
rect 17402 13268 17408 13320
rect 17460 13268 17466 13320
rect 18156 13317 18184 13348
rect 19260 13317 19288 13416
rect 18141 13311 18199 13317
rect 18141 13277 18153 13311
rect 18187 13277 18199 13311
rect 18141 13271 18199 13277
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 21545 13311 21603 13317
rect 19245 13271 19303 13277
rect 10744 13212 11856 13240
rect 10744 13200 10750 13212
rect 11974 13200 11980 13252
rect 12032 13200 12038 13252
rect 12069 13243 12127 13249
rect 12069 13209 12081 13243
rect 12115 13209 12127 13243
rect 12069 13203 12127 13209
rect 20533 13243 20591 13249
rect 20533 13209 20545 13243
rect 20579 13240 20591 13243
rect 20622 13240 20628 13252
rect 20579 13212 20628 13240
rect 20579 13209 20591 13212
rect 20533 13203 20591 13209
rect 5767 13144 7144 13172
rect 5767 13141 5779 13144
rect 5721 13135 5779 13141
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 9766 13132 9772 13184
rect 9824 13172 9830 13184
rect 10137 13175 10195 13181
rect 10137 13172 10149 13175
rect 9824 13144 10149 13172
rect 9824 13132 9830 13144
rect 10137 13141 10149 13144
rect 10183 13141 10195 13175
rect 10137 13135 10195 13141
rect 10502 13132 10508 13184
rect 10560 13172 10566 13184
rect 10781 13175 10839 13181
rect 10781 13172 10793 13175
rect 10560 13144 10793 13172
rect 10560 13132 10566 13144
rect 10781 13141 10793 13144
rect 10827 13141 10839 13175
rect 10781 13135 10839 13141
rect 11241 13175 11299 13181
rect 11241 13141 11253 13175
rect 11287 13172 11299 13175
rect 11514 13172 11520 13184
rect 11287 13144 11520 13172
rect 11287 13141 11299 13144
rect 11241 13135 11299 13141
rect 11514 13132 11520 13144
rect 11572 13132 11578 13184
rect 11698 13132 11704 13184
rect 11756 13172 11762 13184
rect 12084 13172 12112 13203
rect 20622 13200 20628 13212
rect 20680 13200 20686 13252
rect 21468 13240 21496 13294
rect 21545 13277 21557 13311
rect 21591 13308 21603 13311
rect 21818 13308 21824 13320
rect 21591 13280 21824 13308
rect 21591 13277 21603 13280
rect 21545 13271 21603 13277
rect 21818 13268 21824 13280
rect 21876 13268 21882 13320
rect 21726 13240 21732 13252
rect 21468 13212 21732 13240
rect 21726 13200 21732 13212
rect 21784 13240 21790 13252
rect 22278 13240 22284 13252
rect 21784 13212 22284 13240
rect 21784 13200 21790 13212
rect 22278 13200 22284 13212
rect 22336 13200 22342 13252
rect 11756 13144 12112 13172
rect 14185 13175 14243 13181
rect 11756 13132 11762 13144
rect 14185 13141 14197 13175
rect 14231 13172 14243 13175
rect 14826 13172 14832 13184
rect 14231 13144 14832 13172
rect 14231 13141 14243 13144
rect 14185 13135 14243 13141
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 14921 13175 14979 13181
rect 14921 13141 14933 13175
rect 14967 13172 14979 13175
rect 15562 13172 15568 13184
rect 14967 13144 15568 13172
rect 14967 13141 14979 13144
rect 14921 13135 14979 13141
rect 15562 13132 15568 13144
rect 15620 13132 15626 13184
rect 15657 13175 15715 13181
rect 15657 13141 15669 13175
rect 15703 13172 15715 13175
rect 16666 13172 16672 13184
rect 15703 13144 16672 13172
rect 15703 13141 15715 13144
rect 15657 13135 15715 13141
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 16758 13132 16764 13184
rect 16816 13172 16822 13184
rect 17221 13175 17279 13181
rect 17221 13172 17233 13175
rect 16816 13144 17233 13172
rect 16816 13132 16822 13144
rect 17221 13141 17233 13144
rect 17267 13141 17279 13175
rect 17221 13135 17279 13141
rect 18598 13132 18604 13184
rect 18656 13172 18662 13184
rect 18693 13175 18751 13181
rect 18693 13172 18705 13175
rect 18656 13144 18705 13172
rect 18656 13132 18662 13144
rect 18693 13141 18705 13144
rect 18739 13141 18751 13175
rect 18693 13135 18751 13141
rect 19794 13132 19800 13184
rect 19852 13132 19858 13184
rect 1104 13082 22816 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 22816 13082
rect 1104 13008 22816 13030
rect 6086 12928 6092 12980
rect 6144 12968 6150 12980
rect 6144 12940 7144 12968
rect 6144 12928 6150 12940
rect 1486 12860 1492 12912
rect 1544 12900 1550 12912
rect 2501 12903 2559 12909
rect 2501 12900 2513 12903
rect 1544 12872 2513 12900
rect 1544 12860 1550 12872
rect 2501 12869 2513 12872
rect 2547 12869 2559 12903
rect 5074 12900 5080 12912
rect 3726 12886 5080 12900
rect 2501 12863 2559 12869
rect 3712 12872 5080 12886
rect 2133 12767 2191 12773
rect 2133 12733 2145 12767
rect 2179 12733 2191 12767
rect 2133 12727 2191 12733
rect 1762 12656 1768 12708
rect 1820 12656 1826 12708
rect 1673 12631 1731 12637
rect 1673 12597 1685 12631
rect 1719 12628 1731 12631
rect 2038 12628 2044 12640
rect 1719 12600 2044 12628
rect 1719 12597 1731 12600
rect 1673 12591 1731 12597
rect 2038 12588 2044 12600
rect 2096 12588 2102 12640
rect 2148 12628 2176 12727
rect 2222 12724 2228 12776
rect 2280 12724 2286 12776
rect 3142 12724 3148 12776
rect 3200 12764 3206 12776
rect 3712 12764 3740 12872
rect 5074 12860 5080 12872
rect 5132 12860 5138 12912
rect 5166 12860 5172 12912
rect 5224 12860 5230 12912
rect 6730 12900 6736 12912
rect 6564 12872 6736 12900
rect 4338 12792 4344 12844
rect 4396 12792 4402 12844
rect 6362 12792 6368 12844
rect 6420 12832 6426 12844
rect 6564 12841 6592 12872
rect 6730 12860 6736 12872
rect 6788 12900 6794 12912
rect 7009 12903 7067 12909
rect 7009 12900 7021 12903
rect 6788 12872 7021 12900
rect 6788 12860 6794 12872
rect 7009 12869 7021 12872
rect 7055 12869 7067 12903
rect 7009 12863 7067 12869
rect 6549 12835 6607 12841
rect 6549 12832 6561 12835
rect 6420 12804 6561 12832
rect 6420 12792 6426 12804
rect 6549 12801 6561 12804
rect 6595 12801 6607 12835
rect 6549 12795 6607 12801
rect 6825 12835 6883 12841
rect 6825 12801 6837 12835
rect 6871 12832 6883 12835
rect 6914 12832 6920 12844
rect 6871 12804 6920 12832
rect 6871 12801 6883 12804
rect 6825 12795 6883 12801
rect 6914 12792 6920 12804
rect 6972 12792 6978 12844
rect 7116 12841 7144 12940
rect 7190 12928 7196 12980
rect 7248 12968 7254 12980
rect 9398 12968 9404 12980
rect 7248 12940 9404 12968
rect 7248 12928 7254 12940
rect 9398 12928 9404 12940
rect 9456 12928 9462 12980
rect 9674 12928 9680 12980
rect 9732 12968 9738 12980
rect 9732 12940 9904 12968
rect 9732 12928 9738 12940
rect 9490 12900 9496 12912
rect 9062 12872 9496 12900
rect 9490 12860 9496 12872
rect 9548 12860 9554 12912
rect 9766 12860 9772 12912
rect 9824 12860 9830 12912
rect 9876 12900 9904 12940
rect 13262 12928 13268 12980
rect 13320 12928 13326 12980
rect 14734 12928 14740 12980
rect 14792 12928 14798 12980
rect 15470 12928 15476 12980
rect 15528 12928 15534 12980
rect 16114 12928 16120 12980
rect 16172 12968 16178 12980
rect 16209 12971 16267 12977
rect 16209 12968 16221 12971
rect 16172 12940 16221 12968
rect 16172 12928 16178 12940
rect 16209 12937 16221 12940
rect 16255 12937 16267 12971
rect 16209 12931 16267 12937
rect 13814 12900 13820 12912
rect 9876 12872 10258 12900
rect 13018 12872 13820 12900
rect 13814 12860 13820 12872
rect 13872 12860 13878 12912
rect 16666 12860 16672 12912
rect 16724 12860 16730 12912
rect 17862 12860 17868 12912
rect 17920 12860 17926 12912
rect 18598 12860 18604 12912
rect 18656 12860 18662 12912
rect 18874 12860 18880 12912
rect 18932 12860 18938 12912
rect 19978 12900 19984 12912
rect 19812 12872 19984 12900
rect 7101 12835 7159 12841
rect 7101 12801 7113 12835
rect 7147 12801 7159 12835
rect 7101 12795 7159 12801
rect 7198 12835 7256 12841
rect 7198 12801 7210 12835
rect 7244 12832 7256 12835
rect 7244 12804 7328 12832
rect 7244 12801 7256 12804
rect 7198 12795 7256 12801
rect 3200 12736 3740 12764
rect 3200 12724 3206 12736
rect 4614 12724 4620 12776
rect 4672 12724 4678 12776
rect 6178 12724 6184 12776
rect 6236 12764 6242 12776
rect 7300 12764 7328 12804
rect 11514 12792 11520 12844
rect 11572 12792 11578 12844
rect 13446 12792 13452 12844
rect 13504 12792 13510 12844
rect 14185 12835 14243 12841
rect 14185 12832 14197 12835
rect 14016 12804 14197 12832
rect 6236 12736 7328 12764
rect 6236 12724 6242 12736
rect 7466 12724 7472 12776
rect 7524 12764 7530 12776
rect 7561 12767 7619 12773
rect 7561 12764 7573 12767
rect 7524 12736 7573 12764
rect 7524 12724 7530 12736
rect 7561 12733 7573 12736
rect 7607 12733 7619 12767
rect 7837 12767 7895 12773
rect 7837 12764 7849 12767
rect 7561 12727 7619 12733
rect 7668 12736 7849 12764
rect 7377 12699 7435 12705
rect 7377 12665 7389 12699
rect 7423 12696 7435 12699
rect 7668 12696 7696 12736
rect 7837 12733 7849 12736
rect 7883 12733 7895 12767
rect 7837 12727 7895 12733
rect 9309 12767 9367 12773
rect 9309 12733 9321 12767
rect 9355 12764 9367 12767
rect 9493 12767 9551 12773
rect 9493 12764 9505 12767
rect 9355 12736 9505 12764
rect 9355 12733 9367 12736
rect 9309 12727 9367 12733
rect 9493 12733 9505 12736
rect 9539 12764 9551 12767
rect 11146 12764 11152 12776
rect 9539 12736 11152 12764
rect 9539 12733 9551 12736
rect 9493 12727 9551 12733
rect 11146 12724 11152 12736
rect 11204 12724 11210 12776
rect 14016 12773 14044 12804
rect 14185 12801 14197 12804
rect 14231 12801 14243 12835
rect 14185 12795 14243 12801
rect 14826 12792 14832 12844
rect 14884 12832 14890 12844
rect 14921 12835 14979 12841
rect 14921 12832 14933 12835
rect 14884 12804 14933 12832
rect 14884 12792 14890 12804
rect 14921 12801 14933 12804
rect 14967 12801 14979 12835
rect 14921 12795 14979 12801
rect 15562 12792 15568 12844
rect 15620 12832 15626 12844
rect 15657 12835 15715 12841
rect 15657 12832 15669 12835
rect 15620 12804 15669 12832
rect 15620 12792 15626 12804
rect 15657 12801 15669 12804
rect 15703 12801 15715 12835
rect 15657 12795 15715 12801
rect 16022 12792 16028 12844
rect 16080 12832 16086 12844
rect 17405 12835 17463 12841
rect 17405 12832 17417 12835
rect 16080 12804 17417 12832
rect 16080 12792 16086 12804
rect 17405 12801 17417 12804
rect 17451 12801 17463 12835
rect 17405 12795 17463 12801
rect 19610 12792 19616 12844
rect 19668 12792 19674 12844
rect 19812 12841 19840 12872
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 22094 12900 22100 12912
rect 21298 12872 22100 12900
rect 22094 12860 22100 12872
rect 22152 12900 22158 12912
rect 22646 12900 22652 12912
rect 22152 12872 22652 12900
rect 22152 12860 22158 12872
rect 22646 12860 22652 12872
rect 22704 12860 22710 12912
rect 19797 12835 19855 12841
rect 19797 12801 19809 12835
rect 19843 12801 19855 12835
rect 19797 12795 19855 12801
rect 11241 12767 11299 12773
rect 11241 12733 11253 12767
rect 11287 12764 11299 12767
rect 11793 12767 11851 12773
rect 11793 12764 11805 12767
rect 11287 12736 11805 12764
rect 11287 12733 11299 12736
rect 11241 12727 11299 12733
rect 11793 12733 11805 12736
rect 11839 12733 11851 12767
rect 11793 12727 11851 12733
rect 14001 12767 14059 12773
rect 14001 12733 14013 12767
rect 14047 12733 14059 12767
rect 14001 12727 14059 12733
rect 20073 12767 20131 12773
rect 20073 12733 20085 12767
rect 20119 12764 20131 12767
rect 20806 12764 20812 12776
rect 20119 12736 20812 12764
rect 20119 12733 20131 12736
rect 20073 12727 20131 12733
rect 20806 12724 20812 12736
rect 20864 12724 20870 12776
rect 21545 12767 21603 12773
rect 21545 12733 21557 12767
rect 21591 12764 21603 12767
rect 22373 12767 22431 12773
rect 22373 12764 22385 12767
rect 21591 12736 22385 12764
rect 21591 12733 21603 12736
rect 21545 12727 21603 12733
rect 22373 12733 22385 12736
rect 22419 12733 22431 12767
rect 22373 12727 22431 12733
rect 7423 12668 7696 12696
rect 7423 12665 7435 12668
rect 7377 12659 7435 12665
rect 3973 12631 4031 12637
rect 3973 12628 3985 12631
rect 2148 12600 3985 12628
rect 3973 12597 3985 12600
rect 4019 12628 4031 12631
rect 4154 12628 4160 12640
rect 4019 12600 4160 12628
rect 4019 12597 4031 12600
rect 3973 12591 4031 12597
rect 4154 12588 4160 12600
rect 4212 12588 4218 12640
rect 6641 12631 6699 12637
rect 6641 12597 6653 12631
rect 6687 12628 6699 12631
rect 7650 12628 7656 12640
rect 6687 12600 7656 12628
rect 6687 12597 6699 12600
rect 6641 12591 6699 12597
rect 7650 12588 7656 12600
rect 7708 12588 7714 12640
rect 21818 12588 21824 12640
rect 21876 12588 21882 12640
rect 1104 12538 22816 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 20214 12538
rect 20266 12486 20278 12538
rect 20330 12486 20342 12538
rect 20394 12486 20406 12538
rect 20458 12486 20470 12538
rect 20522 12486 22816 12538
rect 1104 12464 22816 12486
rect 1581 12427 1639 12433
rect 1581 12393 1593 12427
rect 1627 12424 1639 12427
rect 2222 12424 2228 12436
rect 1627 12396 2228 12424
rect 1627 12393 1639 12396
rect 1581 12387 1639 12393
rect 2222 12384 2228 12396
rect 2280 12384 2286 12436
rect 2406 12384 2412 12436
rect 2464 12424 2470 12436
rect 2464 12396 3832 12424
rect 2464 12384 2470 12396
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12288 1823 12291
rect 2774 12288 2780 12300
rect 1811 12260 2780 12288
rect 1811 12257 1823 12260
rect 1765 12251 1823 12257
rect 2774 12248 2780 12260
rect 2832 12248 2838 12300
rect 1670 12180 1676 12232
rect 1728 12180 1734 12232
rect 3142 12180 3148 12232
rect 3200 12180 3206 12232
rect 3804 12220 3832 12396
rect 3878 12384 3884 12436
rect 3936 12424 3942 12436
rect 3973 12427 4031 12433
rect 3973 12424 3985 12427
rect 3936 12396 3985 12424
rect 3936 12384 3942 12396
rect 3973 12393 3985 12396
rect 4019 12393 4031 12427
rect 3973 12387 4031 12393
rect 4433 12427 4491 12433
rect 4433 12393 4445 12427
rect 4479 12424 4491 12427
rect 4614 12424 4620 12436
rect 4479 12396 4620 12424
rect 4479 12393 4491 12396
rect 4433 12387 4491 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 6730 12384 6736 12436
rect 6788 12424 6794 12436
rect 6788 12396 8524 12424
rect 6788 12384 6794 12396
rect 8496 12365 8524 12396
rect 10686 12384 10692 12436
rect 10744 12424 10750 12436
rect 12621 12427 12679 12433
rect 12621 12424 12633 12427
rect 10744 12396 12633 12424
rect 10744 12384 10750 12396
rect 12621 12393 12633 12396
rect 12667 12393 12679 12427
rect 12621 12387 12679 12393
rect 13173 12427 13231 12433
rect 13173 12393 13185 12427
rect 13219 12424 13231 12427
rect 13446 12424 13452 12436
rect 13219 12396 13452 12424
rect 13219 12393 13231 12396
rect 13173 12387 13231 12393
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 16574 12384 16580 12436
rect 16632 12384 16638 12436
rect 17313 12427 17371 12433
rect 17313 12393 17325 12427
rect 17359 12424 17371 12427
rect 17402 12424 17408 12436
rect 17359 12396 17408 12424
rect 17359 12393 17371 12396
rect 17313 12387 17371 12393
rect 17402 12384 17408 12396
rect 17460 12384 17466 12436
rect 8481 12359 8539 12365
rect 8481 12325 8493 12359
rect 8527 12325 8539 12359
rect 8481 12319 8539 12325
rect 5902 12288 5908 12300
rect 4264 12260 5908 12288
rect 4264 12229 4292 12260
rect 5902 12248 5908 12260
rect 5960 12248 5966 12300
rect 6178 12248 6184 12300
rect 6236 12248 6242 12300
rect 9766 12288 9772 12300
rect 8128 12260 9772 12288
rect 4249 12223 4307 12229
rect 3804 12192 4200 12220
rect 2038 12112 2044 12164
rect 2096 12112 2102 12164
rect 3786 12112 3792 12164
rect 3844 12112 3850 12164
rect 3513 12087 3571 12093
rect 3513 12053 3525 12087
rect 3559 12084 3571 12087
rect 3602 12084 3608 12096
rect 3559 12056 3608 12084
rect 3559 12053 3571 12056
rect 3513 12047 3571 12053
rect 3602 12044 3608 12056
rect 3660 12044 3666 12096
rect 3970 12044 3976 12096
rect 4028 12044 4034 12096
rect 4172 12084 4200 12192
rect 4249 12189 4261 12223
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 6270 12180 6276 12232
rect 6328 12180 6334 12232
rect 8128 12164 8156 12260
rect 9766 12248 9772 12260
rect 9824 12248 9830 12300
rect 10502 12248 10508 12300
rect 10560 12248 10566 12300
rect 10781 12291 10839 12297
rect 10781 12257 10793 12291
rect 10827 12288 10839 12291
rect 11882 12288 11888 12300
rect 10827 12260 11888 12288
rect 10827 12257 10839 12260
rect 10781 12251 10839 12257
rect 11882 12248 11888 12260
rect 11940 12248 11946 12300
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 15841 12291 15899 12297
rect 15841 12288 15853 12291
rect 15804 12260 15853 12288
rect 15804 12248 15810 12260
rect 15841 12257 15853 12260
rect 15887 12288 15899 12291
rect 17773 12291 17831 12297
rect 15887 12260 16068 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 10870 12180 10876 12232
rect 10928 12180 10934 12232
rect 13722 12180 13728 12232
rect 13780 12220 13786 12232
rect 16040 12229 16068 12260
rect 17773 12257 17785 12291
rect 17819 12288 17831 12291
rect 17819 12260 18460 12288
rect 17819 12257 17831 12260
rect 17773 12251 17831 12257
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13780 12192 14105 12220
rect 13780 12180 13786 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 14093 12183 14151 12189
rect 16025 12223 16083 12229
rect 16025 12189 16037 12223
rect 16071 12189 16083 12223
rect 16025 12183 16083 12189
rect 16758 12180 16764 12232
rect 16816 12180 16822 12232
rect 18322 12180 18328 12232
rect 18380 12180 18386 12232
rect 18432 12229 18460 12260
rect 20070 12248 20076 12300
rect 20128 12248 20134 12300
rect 20533 12291 20591 12297
rect 20533 12257 20545 12291
rect 20579 12288 20591 12291
rect 20622 12288 20628 12300
rect 20579 12260 20628 12288
rect 20579 12257 20591 12260
rect 20533 12251 20591 12257
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 22278 12248 22284 12300
rect 22336 12248 22342 12300
rect 18417 12223 18475 12229
rect 18417 12189 18429 12223
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 19245 12223 19303 12229
rect 19245 12189 19257 12223
rect 19291 12220 19303 12223
rect 19794 12220 19800 12232
rect 19291 12192 19800 12220
rect 19291 12189 19303 12192
rect 19245 12183 19303 12189
rect 19794 12180 19800 12192
rect 19852 12180 19858 12232
rect 19978 12180 19984 12232
rect 20036 12220 20042 12232
rect 20257 12223 20315 12229
rect 20257 12220 20269 12223
rect 20036 12192 20269 12220
rect 20036 12180 20042 12192
rect 20257 12189 20269 12192
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 5442 12112 5448 12164
rect 5500 12112 5506 12164
rect 5626 12112 5632 12164
rect 5684 12152 5690 12164
rect 5905 12155 5963 12161
rect 5905 12152 5917 12155
rect 5684 12124 5917 12152
rect 5684 12112 5690 12124
rect 5905 12121 5917 12124
rect 5951 12121 5963 12155
rect 5905 12115 5963 12121
rect 6546 12112 6552 12164
rect 6604 12112 6610 12164
rect 8110 12152 8116 12164
rect 7774 12124 8116 12152
rect 8110 12112 8116 12124
rect 8168 12112 8174 12164
rect 8205 12155 8263 12161
rect 8205 12121 8217 12155
rect 8251 12121 8263 12155
rect 8205 12115 8263 12121
rect 6730 12084 6736 12096
rect 4172 12056 6736 12084
rect 6730 12044 6736 12056
rect 6788 12044 6794 12096
rect 6822 12044 6828 12096
rect 6880 12084 6886 12096
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 6880 12056 8033 12084
rect 6880 12044 6886 12056
rect 8021 12053 8033 12056
rect 8067 12084 8079 12087
rect 8220 12084 8248 12115
rect 9490 12112 9496 12164
rect 9548 12112 9554 12164
rect 11149 12155 11207 12161
rect 11149 12121 11161 12155
rect 11195 12121 11207 12155
rect 12618 12152 12624 12164
rect 12374 12124 12624 12152
rect 11149 12115 11207 12121
rect 8067 12056 8248 12084
rect 8067 12053 8079 12056
rect 8021 12047 8079 12053
rect 8662 12044 8668 12096
rect 8720 12044 8726 12096
rect 9033 12087 9091 12093
rect 9033 12053 9045 12087
rect 9079 12084 9091 12087
rect 11164 12084 11192 12115
rect 12618 12112 12624 12124
rect 12676 12112 12682 12164
rect 14366 12112 14372 12164
rect 14424 12112 14430 12164
rect 22094 12152 22100 12164
rect 15594 12124 19104 12152
rect 21758 12124 22100 12152
rect 9079 12056 11192 12084
rect 9079 12053 9091 12056
rect 9033 12047 9091 12053
rect 14734 12044 14740 12096
rect 14792 12084 14798 12096
rect 15672 12084 15700 12124
rect 14792 12056 15700 12084
rect 14792 12044 14798 12056
rect 18874 12044 18880 12096
rect 18932 12084 18938 12096
rect 18969 12087 19027 12093
rect 18969 12084 18981 12087
rect 18932 12056 18981 12084
rect 18932 12044 18938 12056
rect 18969 12053 18981 12056
rect 19015 12053 19027 12087
rect 19076 12084 19104 12124
rect 21836 12084 21864 12124
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 19076 12056 21864 12084
rect 18969 12047 19027 12053
rect 1104 11994 22816 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 22816 11994
rect 1104 11920 22816 11942
rect 2869 11883 2927 11889
rect 2869 11849 2881 11883
rect 2915 11880 2927 11883
rect 2958 11880 2964 11892
rect 2915 11852 2964 11880
rect 2915 11849 2927 11852
rect 2869 11843 2927 11849
rect 2958 11840 2964 11852
rect 3016 11840 3022 11892
rect 3694 11880 3700 11892
rect 3160 11852 3700 11880
rect 2774 11812 2780 11824
rect 2332 11784 2780 11812
rect 1670 11704 1676 11756
rect 1728 11704 1734 11756
rect 2332 11730 2360 11784
rect 2774 11772 2780 11784
rect 2832 11772 2838 11824
rect 3160 11753 3188 11852
rect 3694 11840 3700 11852
rect 3752 11880 3758 11892
rect 5077 11883 5135 11889
rect 5077 11880 5089 11883
rect 3752 11852 5089 11880
rect 3752 11840 3758 11852
rect 5077 11849 5089 11852
rect 5123 11849 5135 11883
rect 5077 11843 5135 11849
rect 5353 11883 5411 11889
rect 5353 11849 5365 11883
rect 5399 11880 5411 11883
rect 6270 11880 6276 11892
rect 5399 11852 6276 11880
rect 5399 11849 5411 11852
rect 5353 11843 5411 11849
rect 6270 11840 6276 11852
rect 6328 11840 6334 11892
rect 7116 11852 10364 11880
rect 3602 11772 3608 11824
rect 3660 11772 3666 11824
rect 5166 11812 5172 11824
rect 4830 11784 5172 11812
rect 5166 11772 5172 11784
rect 5224 11812 5230 11824
rect 5442 11812 5448 11824
rect 5224 11784 5448 11812
rect 5224 11772 5230 11784
rect 5442 11772 5448 11784
rect 5500 11772 5506 11824
rect 5905 11815 5963 11821
rect 5905 11781 5917 11815
rect 5951 11812 5963 11815
rect 6822 11812 6828 11824
rect 5951 11784 6828 11812
rect 5951 11781 5963 11784
rect 5905 11775 5963 11781
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 7116 11756 7144 11852
rect 7193 11815 7251 11821
rect 7193 11781 7205 11815
rect 7239 11812 7251 11815
rect 8018 11812 8024 11824
rect 7239 11784 8024 11812
rect 7239 11781 7251 11784
rect 7193 11775 7251 11781
rect 8018 11772 8024 11784
rect 8076 11772 8082 11824
rect 8202 11772 8208 11824
rect 8260 11812 8266 11824
rect 9876 11821 9904 11852
rect 10336 11824 10364 11852
rect 10870 11840 10876 11892
rect 10928 11880 10934 11892
rect 11238 11880 11244 11892
rect 10928 11852 11244 11880
rect 10928 11840 10934 11852
rect 11238 11840 11244 11852
rect 11296 11840 11302 11892
rect 14366 11840 14372 11892
rect 14424 11880 14430 11892
rect 15657 11883 15715 11889
rect 15657 11880 15669 11883
rect 14424 11852 15669 11880
rect 14424 11840 14430 11852
rect 15657 11849 15669 11852
rect 15703 11849 15715 11883
rect 15657 11843 15715 11849
rect 18322 11840 18328 11892
rect 18380 11880 18386 11892
rect 18693 11883 18751 11889
rect 18693 11880 18705 11883
rect 18380 11852 18705 11880
rect 18380 11840 18386 11852
rect 18693 11849 18705 11852
rect 18739 11849 18751 11883
rect 18693 11843 18751 11849
rect 19429 11883 19487 11889
rect 19429 11849 19441 11883
rect 19475 11880 19487 11883
rect 19610 11880 19616 11892
rect 19475 11852 19616 11880
rect 19475 11849 19487 11852
rect 19429 11843 19487 11849
rect 19610 11840 19616 11852
rect 19668 11840 19674 11892
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20864 11852 20913 11880
rect 20864 11840 20870 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 9861 11815 9919 11821
rect 8260 11784 8418 11812
rect 8260 11772 8266 11784
rect 9861 11781 9873 11815
rect 9907 11781 9919 11815
rect 9861 11775 9919 11781
rect 10318 11772 10324 11824
rect 10376 11812 10382 11824
rect 12066 11812 12072 11824
rect 10376 11784 10916 11812
rect 10376 11772 10382 11784
rect 2869 11747 2927 11753
rect 2869 11744 2881 11747
rect 2608 11716 2881 11744
rect 1854 11636 1860 11688
rect 1912 11676 1918 11688
rect 2406 11676 2412 11688
rect 1912 11648 2412 11676
rect 1912 11636 1918 11648
rect 2406 11636 2412 11648
rect 2464 11676 2470 11688
rect 2608 11676 2636 11716
rect 2869 11713 2881 11716
rect 2915 11713 2927 11747
rect 2869 11707 2927 11713
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11713 3203 11747
rect 3145 11707 3203 11713
rect 3326 11704 3332 11756
rect 3384 11704 3390 11756
rect 5810 11753 5816 11756
rect 5261 11747 5319 11753
rect 5261 11713 5273 11747
rect 5307 11744 5319 11747
rect 5761 11747 5816 11753
rect 5761 11744 5773 11747
rect 5307 11716 5773 11744
rect 5307 11713 5319 11716
rect 5261 11707 5319 11713
rect 5761 11713 5773 11716
rect 5807 11713 5816 11747
rect 5761 11707 5816 11713
rect 2464 11648 2636 11676
rect 2464 11636 2470 11648
rect 2682 11636 2688 11688
rect 2740 11636 2746 11688
rect 3970 11636 3976 11688
rect 4028 11676 4034 11688
rect 5276 11676 5304 11707
rect 5810 11704 5816 11707
rect 5868 11704 5874 11756
rect 5997 11747 6055 11753
rect 5997 11713 6009 11747
rect 6043 11713 6055 11747
rect 5997 11707 6055 11713
rect 6181 11747 6239 11753
rect 6181 11713 6193 11747
rect 6227 11744 6239 11747
rect 6270 11744 6276 11756
rect 6227 11716 6276 11744
rect 6227 11713 6239 11716
rect 6181 11707 6239 11713
rect 4028 11648 5304 11676
rect 6012 11676 6040 11707
rect 6270 11704 6276 11716
rect 6328 11744 6334 11756
rect 6457 11747 6515 11753
rect 6457 11744 6469 11747
rect 6328 11716 6469 11744
rect 6328 11704 6334 11716
rect 6457 11713 6469 11716
rect 6503 11713 6515 11747
rect 6457 11707 6515 11713
rect 6730 11704 6736 11756
rect 6788 11704 6794 11756
rect 6917 11747 6975 11753
rect 6917 11713 6929 11747
rect 6963 11744 6975 11747
rect 7006 11744 7012 11756
rect 6963 11716 7012 11744
rect 6963 11713 6975 11716
rect 6917 11707 6975 11713
rect 7006 11704 7012 11716
rect 7064 11704 7070 11756
rect 7098 11704 7104 11756
rect 7156 11704 7162 11756
rect 7337 11747 7395 11753
rect 7337 11713 7349 11747
rect 7383 11744 7395 11747
rect 7383 11713 7420 11744
rect 7337 11707 7420 11713
rect 6012 11648 6592 11676
rect 4028 11636 4034 11648
rect 5629 11611 5687 11617
rect 5629 11577 5641 11611
rect 5675 11608 5687 11611
rect 6362 11608 6368 11620
rect 5675 11580 6368 11608
rect 5675 11577 5687 11580
rect 5629 11571 5687 11577
rect 6362 11568 6368 11580
rect 6420 11568 6426 11620
rect 6454 11568 6460 11620
rect 6512 11568 6518 11620
rect 6564 11608 6592 11648
rect 6914 11608 6920 11620
rect 6564 11580 6920 11608
rect 6914 11568 6920 11580
rect 6972 11568 6978 11620
rect 7392 11540 7420 11707
rect 7650 11704 7656 11756
rect 7708 11704 7714 11756
rect 9582 11704 9588 11756
rect 9640 11744 9646 11756
rect 9677 11747 9735 11753
rect 9677 11744 9689 11747
rect 9640 11716 9689 11744
rect 9640 11704 9646 11716
rect 9677 11713 9689 11716
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 9953 11747 10011 11753
rect 9953 11713 9965 11747
rect 9999 11713 10011 11747
rect 9953 11707 10011 11713
rect 10097 11747 10155 11753
rect 10097 11713 10109 11747
rect 10143 11744 10155 11747
rect 10502 11744 10508 11756
rect 10143 11716 10508 11744
rect 10143 11713 10155 11716
rect 10097 11707 10155 11713
rect 7929 11679 7987 11685
rect 7929 11645 7941 11679
rect 7975 11676 7987 11679
rect 8570 11676 8576 11688
rect 7975 11648 8576 11676
rect 7975 11645 7987 11648
rect 7929 11639 7987 11645
rect 8570 11636 8576 11648
rect 8628 11636 8634 11688
rect 9398 11636 9404 11688
rect 9456 11636 9462 11688
rect 7466 11568 7472 11620
rect 7524 11568 7530 11620
rect 8018 11540 8024 11552
rect 7392 11512 8024 11540
rect 8018 11500 8024 11512
rect 8076 11540 8082 11552
rect 9674 11540 9680 11552
rect 8076 11512 9680 11540
rect 8076 11500 8082 11512
rect 9674 11500 9680 11512
rect 9732 11500 9738 11552
rect 9968 11540 9996 11707
rect 10502 11704 10508 11716
rect 10560 11744 10566 11756
rect 10637 11747 10695 11753
rect 10637 11744 10649 11747
rect 10560 11716 10649 11744
rect 10560 11704 10566 11716
rect 10637 11713 10649 11716
rect 10683 11713 10695 11747
rect 10637 11707 10695 11713
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 10888 11753 10916 11784
rect 11164 11784 12072 11812
rect 10873 11747 10931 11753
rect 10873 11713 10885 11747
rect 10919 11713 10931 11747
rect 10873 11707 10931 11713
rect 11054 11704 11060 11756
rect 11112 11704 11118 11756
rect 11164 11753 11192 11784
rect 12066 11772 12072 11784
rect 12124 11812 12130 11824
rect 12124 11784 13860 11812
rect 12124 11772 12130 11784
rect 11149 11747 11207 11753
rect 11149 11713 11161 11747
rect 11195 11713 11207 11747
rect 11149 11707 11207 11713
rect 11164 11676 11192 11707
rect 11606 11704 11612 11756
rect 11664 11704 11670 11756
rect 11885 11747 11943 11753
rect 11885 11713 11897 11747
rect 11931 11744 11943 11747
rect 13538 11744 13544 11756
rect 11931 11716 13544 11744
rect 11931 11713 11943 11716
rect 11885 11707 11943 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13832 11753 13860 11784
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11713 13875 11747
rect 14553 11747 14611 11753
rect 14553 11744 14565 11747
rect 13817 11707 13875 11713
rect 13924 11716 14565 11744
rect 10244 11648 11192 11676
rect 11624 11676 11652 11704
rect 11624 11648 12434 11676
rect 10244 11617 10272 11648
rect 10229 11611 10287 11617
rect 10229 11577 10241 11611
rect 10275 11577 10287 11611
rect 10778 11608 10784 11620
rect 10229 11571 10287 11577
rect 10336 11580 10784 11608
rect 10336 11540 10364 11580
rect 10778 11568 10784 11580
rect 10836 11568 10842 11620
rect 10870 11568 10876 11620
rect 10928 11608 10934 11620
rect 11609 11611 11667 11617
rect 11609 11608 11621 11611
rect 10928 11580 11621 11608
rect 10928 11568 10934 11580
rect 11609 11577 11621 11580
rect 11655 11577 11667 11611
rect 12406 11608 12434 11648
rect 12710 11636 12716 11688
rect 12768 11636 12774 11688
rect 13446 11636 13452 11688
rect 13504 11676 13510 11688
rect 13924 11676 13952 11716
rect 14553 11713 14565 11716
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 14829 11747 14887 11753
rect 14829 11713 14841 11747
rect 14875 11713 14887 11747
rect 14829 11707 14887 11713
rect 13504 11648 13952 11676
rect 14369 11679 14427 11685
rect 13504 11636 13510 11648
rect 14369 11645 14381 11679
rect 14415 11676 14427 11679
rect 14844 11676 14872 11707
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 16666 11704 16672 11756
rect 16724 11704 16730 11756
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11713 17463 11747
rect 17405 11707 17463 11713
rect 18141 11747 18199 11753
rect 18141 11713 18153 11747
rect 18187 11713 18199 11747
rect 18141 11707 18199 11713
rect 14415 11648 14872 11676
rect 17221 11679 17279 11685
rect 14415 11645 14427 11648
rect 14369 11639 14427 11645
rect 17221 11645 17233 11679
rect 17267 11676 17279 11679
rect 17420 11676 17448 11707
rect 17267 11648 17448 11676
rect 17957 11679 18015 11685
rect 17267 11645 17279 11648
rect 17221 11639 17279 11645
rect 17957 11645 17969 11679
rect 18003 11676 18015 11679
rect 18156 11676 18184 11707
rect 18874 11704 18880 11756
rect 18932 11704 18938 11756
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11744 21051 11747
rect 21818 11744 21824 11756
rect 21039 11716 21824 11744
rect 21039 11713 21051 11716
rect 20993 11707 21051 11713
rect 21818 11704 21824 11716
rect 21876 11704 21882 11756
rect 18003 11648 18184 11676
rect 18003 11645 18015 11648
rect 17957 11639 18015 11645
rect 12989 11611 13047 11617
rect 12989 11608 13001 11611
rect 12406 11580 13001 11608
rect 11609 11571 11667 11577
rect 12989 11577 13001 11580
rect 13035 11577 13047 11611
rect 12989 11571 13047 11577
rect 14645 11611 14703 11617
rect 14645 11577 14657 11611
rect 14691 11608 14703 11611
rect 16022 11608 16028 11620
rect 14691 11580 16028 11608
rect 14691 11577 14703 11580
rect 14645 11571 14703 11577
rect 16022 11568 16028 11580
rect 16080 11568 16086 11620
rect 9968 11512 10364 11540
rect 10505 11543 10563 11549
rect 10505 11509 10517 11543
rect 10551 11540 10563 11543
rect 11146 11540 11152 11552
rect 10551 11512 11152 11540
rect 10551 11509 10563 11512
rect 10505 11503 10563 11509
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 13173 11543 13231 11549
rect 13173 11509 13185 11543
rect 13219 11540 13231 11543
rect 13354 11540 13360 11552
rect 13219 11512 13360 11540
rect 13219 11509 13231 11512
rect 13173 11503 13231 11509
rect 13354 11500 13360 11512
rect 13412 11500 13418 11552
rect 15378 11500 15384 11552
rect 15436 11500 15442 11552
rect 1104 11450 22816 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 20214 11450
rect 20266 11398 20278 11450
rect 20330 11398 20342 11450
rect 20394 11398 20406 11450
rect 20458 11398 20470 11450
rect 20522 11398 22816 11450
rect 1104 11376 22816 11398
rect 1857 11339 1915 11345
rect 1857 11305 1869 11339
rect 1903 11336 1915 11339
rect 2774 11336 2780 11348
rect 1903 11308 2780 11336
rect 1903 11305 1915 11308
rect 1857 11299 1915 11305
rect 2774 11296 2780 11308
rect 2832 11336 2838 11348
rect 3878 11336 3884 11348
rect 2832 11308 3884 11336
rect 2832 11296 2838 11308
rect 3878 11296 3884 11308
rect 3936 11296 3942 11348
rect 5442 11296 5448 11348
rect 5500 11336 5506 11348
rect 5500 11308 6316 11336
rect 5500 11296 5506 11308
rect 6288 11268 6316 11308
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 6733 11339 6791 11345
rect 6733 11336 6745 11339
rect 6604 11308 6745 11336
rect 6604 11296 6610 11308
rect 6733 11305 6745 11308
rect 6779 11305 6791 11339
rect 6733 11299 6791 11305
rect 7180 11339 7238 11345
rect 7180 11305 7192 11339
rect 7226 11336 7238 11339
rect 8662 11336 8668 11348
rect 7226 11308 8668 11336
rect 7226 11305 7238 11308
rect 7180 11299 7238 11305
rect 8662 11296 8668 11308
rect 8720 11296 8726 11348
rect 9401 11339 9459 11345
rect 9401 11305 9413 11339
rect 9447 11336 9459 11339
rect 9447 11308 11100 11336
rect 9447 11305 9459 11308
rect 9401 11299 9459 11305
rect 11072 11268 11100 11308
rect 12710 11296 12716 11348
rect 12768 11336 12774 11348
rect 12989 11339 13047 11345
rect 12989 11336 13001 11339
rect 12768 11308 13001 11336
rect 12768 11296 12774 11308
rect 12989 11305 13001 11308
rect 13035 11305 13047 11339
rect 12989 11299 13047 11305
rect 4264 11240 5028 11268
rect 6288 11240 6592 11268
rect 11072 11240 11376 11268
rect 2682 11160 2688 11212
rect 2740 11200 2746 11212
rect 3329 11203 3387 11209
rect 3329 11200 3341 11203
rect 2740 11172 3341 11200
rect 2740 11160 2746 11172
rect 3329 11169 3341 11172
rect 3375 11169 3387 11203
rect 3329 11163 3387 11169
rect 3878 11160 3884 11212
rect 3936 11160 3942 11212
rect 3970 11160 3976 11212
rect 4028 11200 4034 11212
rect 4264 11200 4292 11240
rect 5000 11209 5028 11240
rect 4028 11172 4292 11200
rect 4028 11160 4034 11172
rect 3602 11092 3608 11144
rect 3660 11092 3666 11144
rect 3786 11092 3792 11144
rect 3844 11132 3850 11144
rect 4065 11135 4123 11141
rect 4065 11132 4077 11135
rect 3844 11104 4077 11132
rect 3844 11092 3850 11104
rect 4065 11101 4077 11104
rect 4111 11101 4123 11135
rect 4264 11132 4292 11172
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 4985 11203 5043 11209
rect 4387 11172 4660 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 4632 11141 4660 11172
rect 4985 11169 4997 11203
rect 5031 11169 5043 11203
rect 4985 11163 5043 11169
rect 5261 11203 5319 11209
rect 5261 11169 5273 11203
rect 5307 11200 5319 11203
rect 6454 11200 6460 11212
rect 5307 11172 6460 11200
rect 5307 11169 5319 11172
rect 5261 11163 5319 11169
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 4433 11135 4491 11141
rect 4433 11132 4445 11135
rect 4264 11104 4445 11132
rect 4065 11095 4123 11101
rect 4433 11101 4445 11104
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 4617 11135 4675 11141
rect 4617 11101 4629 11135
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 4893 11135 4951 11141
rect 4893 11101 4905 11135
rect 4939 11101 4951 11135
rect 4893 11095 4951 11101
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 2924 11036 4476 11064
rect 2924 11024 2930 11036
rect 4448 10996 4476 11036
rect 4522 11024 4528 11076
rect 4580 11024 4586 11076
rect 4908 11064 4936 11095
rect 6564 11064 6592 11240
rect 6914 11160 6920 11212
rect 6972 11200 6978 11212
rect 6972 11172 8984 11200
rect 6972 11160 6978 11172
rect 8956 11141 8984 11172
rect 10870 11160 10876 11212
rect 10928 11160 10934 11212
rect 11146 11160 11152 11212
rect 11204 11160 11210 11212
rect 11238 11160 11244 11212
rect 11296 11160 11302 11212
rect 11348 11200 11376 11240
rect 11517 11203 11575 11209
rect 11517 11200 11529 11203
rect 11348 11172 11529 11200
rect 11517 11169 11529 11172
rect 11563 11169 11575 11203
rect 11517 11163 11575 11169
rect 12066 11160 12072 11212
rect 12124 11200 12130 11212
rect 12124 11172 12940 11200
rect 12124 11160 12130 11172
rect 8941 11135 8999 11141
rect 8941 11101 8953 11135
rect 8987 11101 8999 11135
rect 8941 11095 8999 11101
rect 9398 11092 9404 11144
rect 9456 11132 9462 11144
rect 9456 11104 9798 11132
rect 9456 11092 9462 11104
rect 12618 11092 12624 11144
rect 12676 11092 12682 11144
rect 8846 11064 8852 11076
rect 4908 11036 5212 11064
rect 6486 11036 6592 11064
rect 8418 11036 8852 11064
rect 4890 10996 4896 11008
rect 4448 10968 4896 10996
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 5184 10996 5212 11036
rect 5902 10996 5908 11008
rect 5184 10968 5908 10996
rect 5902 10956 5908 10968
rect 5960 10956 5966 11008
rect 6564 10996 6592 11036
rect 7558 10996 7564 11008
rect 6564 10968 7564 10996
rect 7558 10956 7564 10968
rect 7616 10996 7622 11008
rect 8496 10996 8524 11036
rect 8846 11024 8852 11036
rect 8904 11024 8910 11076
rect 10962 11024 10968 11076
rect 11020 11064 11026 11076
rect 11020 11036 12434 11064
rect 11020 11024 11026 11036
rect 7616 10968 8524 10996
rect 7616 10956 7622 10968
rect 8662 10956 8668 11008
rect 8720 10956 8726 11008
rect 9030 10956 9036 11008
rect 9088 10956 9094 11008
rect 9582 10956 9588 11008
rect 9640 10996 9646 11008
rect 10594 10996 10600 11008
rect 9640 10968 10600 10996
rect 9640 10956 9646 10968
rect 10594 10956 10600 10968
rect 10652 10996 10658 11008
rect 11054 10996 11060 11008
rect 10652 10968 11060 10996
rect 10652 10956 10658 10968
rect 11054 10956 11060 10968
rect 11112 10996 11118 11008
rect 11330 10996 11336 11008
rect 11112 10968 11336 10996
rect 11112 10956 11118 10968
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 12406 10996 12434 11036
rect 12636 10996 12664 11092
rect 12912 11064 12940 11172
rect 13004 11132 13032 11299
rect 13722 11296 13728 11348
rect 13780 11296 13786 11348
rect 16666 11296 16672 11348
rect 16724 11296 16730 11348
rect 14277 11203 14335 11209
rect 14277 11169 14289 11203
rect 14323 11169 14335 11203
rect 14277 11163 14335 11169
rect 13173 11135 13231 11141
rect 13173 11132 13185 11135
rect 13004 11104 13185 11132
rect 13173 11101 13185 11104
rect 13219 11101 13231 11135
rect 13173 11095 13231 11101
rect 13446 11092 13452 11144
rect 13504 11092 13510 11144
rect 13538 11092 13544 11144
rect 13596 11141 13602 11144
rect 13596 11132 13604 11141
rect 14292 11132 14320 11163
rect 15378 11160 15384 11212
rect 15436 11200 15442 11212
rect 15436 11172 16160 11200
rect 15436 11160 15442 11172
rect 13596 11104 14320 11132
rect 13596 11095 13604 11104
rect 13596 11092 13602 11095
rect 16022 11092 16028 11144
rect 16080 11092 16086 11144
rect 16132 11141 16160 11172
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 13357 11067 13415 11073
rect 13357 11064 13369 11067
rect 12912 11036 13369 11064
rect 13357 11033 13369 11036
rect 13403 11033 13415 11067
rect 13357 11027 13415 11033
rect 13814 11024 13820 11076
rect 13872 11064 13878 11076
rect 13872 11036 14582 11064
rect 13872 11024 13878 11036
rect 12406 10968 12664 10996
rect 14476 10996 14504 11036
rect 15746 11024 15752 11076
rect 15804 11024 15810 11076
rect 15010 10996 15016 11008
rect 14476 10968 15016 10996
rect 15010 10956 15016 10968
rect 15068 10956 15074 11008
rect 1104 10906 22816 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 22816 10906
rect 1104 10832 22816 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 1728 10764 3709 10792
rect 1728 10752 1734 10764
rect 3697 10761 3709 10764
rect 3743 10792 3755 10795
rect 3786 10792 3792 10804
rect 3743 10764 3792 10792
rect 3743 10761 3755 10764
rect 3697 10755 3755 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 5810 10752 5816 10804
rect 5868 10792 5874 10804
rect 5905 10795 5963 10801
rect 5905 10792 5917 10795
rect 5868 10764 5917 10792
rect 5868 10752 5874 10764
rect 5905 10761 5917 10764
rect 5951 10761 5963 10795
rect 9030 10792 9036 10804
rect 5905 10755 5963 10761
rect 7208 10764 9036 10792
rect 1765 10727 1823 10733
rect 1765 10693 1777 10727
rect 1811 10724 1823 10727
rect 2225 10727 2283 10733
rect 2225 10724 2237 10727
rect 1811 10696 2237 10724
rect 1811 10693 1823 10696
rect 1765 10687 1823 10693
rect 2225 10693 2237 10696
rect 2271 10693 2283 10727
rect 2225 10687 2283 10693
rect 2866 10684 2872 10736
rect 2924 10684 2930 10736
rect 4433 10727 4491 10733
rect 4433 10693 4445 10727
rect 4479 10724 4491 10727
rect 4522 10724 4528 10736
rect 4479 10696 4528 10724
rect 4479 10693 4491 10696
rect 4433 10687 4491 10693
rect 4522 10684 4528 10696
rect 4580 10684 4586 10736
rect 4890 10684 4896 10736
rect 4948 10684 4954 10736
rect 1670 10616 1676 10668
rect 1728 10616 1734 10668
rect 5902 10616 5908 10668
rect 5960 10656 5966 10668
rect 7208 10665 7236 10764
rect 9030 10752 9036 10764
rect 9088 10752 9094 10804
rect 9674 10752 9680 10804
rect 9732 10792 9738 10804
rect 10502 10792 10508 10804
rect 9732 10764 10508 10792
rect 9732 10752 9738 10764
rect 8846 10684 8852 10736
rect 8904 10684 8910 10736
rect 9048 10724 9076 10752
rect 9048 10696 9628 10724
rect 9600 10665 9628 10696
rect 9950 10684 9956 10736
rect 10008 10684 10014 10736
rect 6733 10659 6791 10665
rect 6733 10656 6745 10659
rect 5960 10628 6745 10656
rect 5960 10616 5966 10628
rect 6733 10625 6745 10628
rect 6779 10625 6791 10659
rect 6733 10619 6791 10625
rect 7193 10659 7251 10665
rect 7193 10625 7205 10659
rect 7239 10625 7251 10659
rect 7193 10619 7251 10625
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10244 10665 10272 10764
rect 10502 10752 10508 10764
rect 10560 10792 10566 10804
rect 11054 10792 11060 10804
rect 10560 10764 11060 10792
rect 10560 10752 10566 10764
rect 11054 10752 11060 10764
rect 11112 10792 11118 10804
rect 14829 10795 14887 10801
rect 11112 10764 11980 10792
rect 11112 10752 11118 10764
rect 10318 10684 10324 10736
rect 10376 10724 10382 10736
rect 10689 10727 10747 10733
rect 10689 10724 10701 10727
rect 10376 10696 10701 10724
rect 10376 10684 10382 10696
rect 10689 10693 10701 10696
rect 10735 10724 10747 10727
rect 10735 10696 11744 10724
rect 10735 10693 10747 10696
rect 10689 10687 10747 10693
rect 11716 10668 11744 10696
rect 10594 10665 10600 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9732 10628 9781 10656
rect 9732 10616 9738 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 10042 10659 10100 10665
rect 10042 10656 10054 10659
rect 9769 10619 9827 10625
rect 9968 10628 10054 10656
rect 1946 10548 1952 10600
rect 2004 10548 2010 10600
rect 4154 10548 4160 10600
rect 4212 10548 4218 10600
rect 5810 10548 5816 10600
rect 5868 10588 5874 10600
rect 6365 10591 6423 10597
rect 6365 10588 6377 10591
rect 5868 10560 6377 10588
rect 5868 10548 5874 10560
rect 6365 10557 6377 10560
rect 6411 10557 6423 10591
rect 6365 10551 6423 10557
rect 6454 10548 6460 10600
rect 6512 10588 6518 10600
rect 7837 10591 7895 10597
rect 7837 10588 7849 10591
rect 6512 10560 7849 10588
rect 6512 10548 6518 10560
rect 7837 10557 7849 10560
rect 7883 10557 7895 10591
rect 7837 10551 7895 10557
rect 8662 10548 8668 10600
rect 8720 10588 8726 10600
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 8720 10560 9321 10588
rect 8720 10548 8726 10560
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 9968 10520 9996 10628
rect 10042 10625 10054 10628
rect 10088 10625 10100 10659
rect 10042 10619 10100 10625
rect 10189 10659 10272 10665
rect 10189 10625 10201 10659
rect 10235 10628 10272 10659
rect 10551 10659 10600 10665
rect 10235 10625 10247 10628
rect 10189 10619 10247 10625
rect 10551 10625 10563 10659
rect 10597 10625 10600 10659
rect 10551 10619 10600 10625
rect 10594 10616 10600 10619
rect 10652 10616 10658 10668
rect 10778 10616 10784 10668
rect 10836 10616 10842 10668
rect 10925 10659 10983 10665
rect 10925 10625 10937 10659
rect 10971 10656 10983 10659
rect 11054 10656 11060 10668
rect 10971 10628 11060 10656
rect 10971 10625 10983 10628
rect 10925 10619 10983 10625
rect 11054 10616 11060 10628
rect 11112 10616 11118 10668
rect 11330 10616 11336 10668
rect 11388 10656 11394 10668
rect 11517 10659 11575 10665
rect 11517 10656 11529 10659
rect 11388 10628 11529 10656
rect 11388 10616 11394 10628
rect 11517 10625 11529 10628
rect 11563 10625 11575 10659
rect 11517 10619 11575 10625
rect 11698 10616 11704 10668
rect 11756 10616 11762 10668
rect 11790 10616 11796 10668
rect 11848 10616 11854 10668
rect 11952 10665 11980 10764
rect 14829 10761 14841 10795
rect 14875 10792 14887 10795
rect 15746 10792 15752 10804
rect 14875 10764 15752 10792
rect 14875 10761 14887 10764
rect 14829 10755 14887 10761
rect 15746 10752 15752 10764
rect 15804 10752 15810 10804
rect 16761 10795 16819 10801
rect 16761 10761 16773 10795
rect 16807 10792 16819 10795
rect 16807 10764 18828 10792
rect 16807 10761 16819 10764
rect 16761 10755 16819 10761
rect 13354 10684 13360 10736
rect 13412 10684 13418 10736
rect 13814 10684 13820 10736
rect 13872 10684 13878 10736
rect 15473 10727 15531 10733
rect 15473 10693 15485 10727
rect 15519 10724 15531 10727
rect 15930 10724 15936 10736
rect 15519 10696 15936 10724
rect 15519 10693 15531 10696
rect 15473 10687 15531 10693
rect 15930 10684 15936 10696
rect 15988 10724 15994 10736
rect 15988 10696 16712 10724
rect 15988 10684 15994 10696
rect 11937 10659 11980 10665
rect 11937 10625 11949 10659
rect 11937 10619 11980 10625
rect 11974 10616 11980 10619
rect 12032 10616 12038 10668
rect 15286 10665 15292 10668
rect 15284 10619 15292 10665
rect 15286 10616 15292 10619
rect 15344 10616 15350 10668
rect 15381 10659 15439 10665
rect 15381 10625 15393 10659
rect 15427 10625 15439 10659
rect 15381 10619 15439 10625
rect 10796 10588 10824 10616
rect 11808 10588 11836 10616
rect 10796 10560 11836 10588
rect 13081 10591 13139 10597
rect 10796 10520 10824 10560
rect 13081 10557 13093 10591
rect 13127 10588 13139 10591
rect 13446 10588 13452 10600
rect 13127 10560 13452 10588
rect 13127 10557 13139 10560
rect 13081 10551 13139 10557
rect 13446 10548 13452 10560
rect 13504 10548 13510 10600
rect 15396 10588 15424 10619
rect 15654 10616 15660 10668
rect 15712 10656 15718 10668
rect 16684 10665 16712 10696
rect 18800 10665 18828 10764
rect 16669 10659 16727 10665
rect 15712 10628 15884 10656
rect 15712 10616 15718 10628
rect 15746 10588 15752 10600
rect 15396 10560 15752 10588
rect 15746 10548 15752 10560
rect 15804 10548 15810 10600
rect 15856 10588 15884 10628
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 18785 10659 18843 10665
rect 16669 10619 16727 10625
rect 17037 10591 17095 10597
rect 17037 10588 17049 10591
rect 15856 10560 17049 10588
rect 17037 10557 17049 10560
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 9646 10492 10824 10520
rect 11057 10523 11115 10529
rect 4890 10412 4896 10464
rect 4948 10452 4954 10464
rect 6270 10452 6276 10464
rect 4948 10424 6276 10452
rect 4948 10412 4954 10424
rect 6270 10412 6276 10424
rect 6328 10412 6334 10464
rect 8110 10412 8116 10464
rect 8168 10452 8174 10464
rect 9646 10452 9674 10492
rect 11057 10489 11069 10523
rect 11103 10520 11115 10523
rect 16025 10523 16083 10529
rect 16025 10520 16037 10523
rect 11103 10492 12434 10520
rect 11103 10489 11115 10492
rect 11057 10483 11115 10489
rect 8168 10424 9674 10452
rect 10321 10455 10379 10461
rect 8168 10412 8174 10424
rect 10321 10421 10333 10455
rect 10367 10452 10379 10455
rect 11514 10452 11520 10464
rect 10367 10424 11520 10452
rect 10367 10421 10379 10424
rect 10321 10415 10379 10421
rect 11514 10412 11520 10424
rect 11572 10412 11578 10464
rect 11882 10412 11888 10464
rect 11940 10452 11946 10464
rect 12069 10455 12127 10461
rect 12069 10452 12081 10455
rect 11940 10424 12081 10452
rect 11940 10412 11946 10424
rect 12069 10421 12081 10424
rect 12115 10421 12127 10455
rect 12406 10452 12434 10492
rect 14384 10492 16037 10520
rect 12986 10452 12992 10464
rect 12406 10424 12992 10452
rect 12069 10415 12127 10421
rect 12986 10412 12992 10424
rect 13044 10412 13050 10464
rect 13906 10412 13912 10464
rect 13964 10452 13970 10464
rect 14384 10452 14412 10492
rect 16025 10489 16037 10492
rect 16071 10489 16083 10523
rect 16025 10483 16083 10489
rect 16574 10480 16580 10532
rect 16632 10520 16638 10532
rect 17420 10520 17448 10642
rect 18785 10625 18797 10659
rect 18831 10625 18843 10659
rect 18785 10619 18843 10625
rect 17954 10548 17960 10600
rect 18012 10588 18018 10600
rect 18509 10591 18567 10597
rect 18509 10588 18521 10591
rect 18012 10560 18521 10588
rect 18012 10548 18018 10560
rect 18509 10557 18521 10560
rect 18555 10557 18567 10591
rect 18509 10551 18567 10557
rect 16632 10492 17448 10520
rect 16632 10480 16638 10492
rect 13964 10424 14412 10452
rect 13964 10412 13970 10424
rect 15102 10412 15108 10464
rect 15160 10412 15166 10464
rect 16209 10455 16267 10461
rect 16209 10421 16221 10455
rect 16255 10452 16267 10455
rect 16482 10452 16488 10464
rect 16255 10424 16488 10452
rect 16255 10421 16267 10424
rect 16209 10415 16267 10421
rect 16482 10412 16488 10424
rect 16540 10412 16546 10464
rect 1104 10362 22816 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 20214 10362
rect 20266 10310 20278 10362
rect 20330 10310 20342 10362
rect 20394 10310 20406 10362
rect 20458 10310 20470 10362
rect 20522 10310 22816 10362
rect 1104 10288 22816 10310
rect 1857 10251 1915 10257
rect 1857 10217 1869 10251
rect 1903 10248 1915 10251
rect 1946 10248 1952 10260
rect 1903 10220 1952 10248
rect 1903 10217 1915 10220
rect 1857 10211 1915 10217
rect 1946 10208 1952 10220
rect 2004 10208 2010 10260
rect 2866 10248 2872 10260
rect 2051 10220 2872 10248
rect 2051 10053 2079 10220
rect 2866 10208 2872 10220
rect 2924 10208 2930 10260
rect 3053 10251 3111 10257
rect 3053 10217 3065 10251
rect 3099 10248 3111 10251
rect 3602 10248 3608 10260
rect 3099 10220 3608 10248
rect 3099 10217 3111 10220
rect 3053 10211 3111 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 4062 10208 4068 10260
rect 4120 10248 4126 10260
rect 4341 10251 4399 10257
rect 4341 10248 4353 10251
rect 4120 10220 4353 10248
rect 4120 10208 4126 10220
rect 4341 10217 4353 10220
rect 4387 10217 4399 10251
rect 5994 10248 6000 10260
rect 4341 10211 4399 10217
rect 5276 10220 6000 10248
rect 2498 10140 2504 10192
rect 2556 10180 2562 10192
rect 3786 10180 3792 10192
rect 2556 10152 3792 10180
rect 2556 10140 2562 10152
rect 3786 10140 3792 10152
rect 3844 10180 3850 10192
rect 4798 10180 4804 10192
rect 3844 10152 4804 10180
rect 3844 10140 3850 10152
rect 4798 10140 4804 10152
rect 4856 10140 4862 10192
rect 2148 10084 2820 10112
rect 2148 10056 2176 10084
rect 2036 10047 2094 10053
rect 2036 10013 2048 10047
rect 2082 10013 2094 10047
rect 2036 10007 2094 10013
rect 2130 10004 2136 10056
rect 2188 10004 2194 10056
rect 2409 10047 2467 10053
rect 2409 10013 2421 10047
rect 2455 10044 2467 10047
rect 2498 10044 2504 10056
rect 2455 10016 2504 10044
rect 2455 10013 2467 10016
rect 2409 10007 2467 10013
rect 2498 10004 2504 10016
rect 2556 10004 2562 10056
rect 2792 9985 2820 10084
rect 3878 10072 3884 10124
rect 3936 10112 3942 10124
rect 5276 10112 5304 10220
rect 5994 10208 6000 10220
rect 6052 10248 6058 10260
rect 6052 10220 6868 10248
rect 6052 10208 6058 10220
rect 5353 10183 5411 10189
rect 5353 10149 5365 10183
rect 5399 10180 5411 10183
rect 6840 10180 6868 10220
rect 6914 10208 6920 10260
rect 6972 10248 6978 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 6972 10220 7297 10248
rect 6972 10208 6978 10220
rect 7285 10217 7297 10220
rect 7331 10217 7343 10251
rect 7285 10211 7343 10217
rect 11330 10208 11336 10260
rect 11388 10248 11394 10260
rect 11606 10248 11612 10260
rect 11388 10220 11612 10248
rect 11388 10208 11394 10220
rect 11606 10208 11612 10220
rect 11664 10208 11670 10260
rect 13265 10251 13323 10257
rect 13265 10217 13277 10251
rect 13311 10248 13323 10251
rect 13446 10248 13452 10260
rect 13311 10220 13452 10248
rect 13311 10217 13323 10220
rect 13265 10211 13323 10217
rect 13446 10208 13452 10220
rect 13504 10208 13510 10260
rect 15654 10248 15660 10260
rect 13740 10220 15660 10248
rect 8018 10180 8024 10192
rect 5399 10152 5580 10180
rect 6840 10152 8024 10180
rect 5399 10149 5411 10152
rect 5353 10143 5411 10149
rect 5552 10121 5580 10152
rect 8018 10140 8024 10152
rect 8076 10180 8082 10192
rect 8389 10183 8447 10189
rect 8076 10152 8253 10180
rect 8076 10140 8082 10152
rect 3936 10084 5304 10112
rect 3936 10072 3942 10084
rect 2866 10004 2872 10056
rect 2924 10053 2930 10056
rect 2924 10047 2979 10053
rect 2924 10013 2933 10047
rect 2967 10044 2979 10047
rect 3694 10044 3700 10056
rect 2967 10016 3700 10044
rect 2967 10013 2979 10016
rect 2924 10007 2979 10013
rect 2924 10004 2930 10007
rect 3694 10004 3700 10016
rect 3752 10004 3758 10056
rect 3786 10004 3792 10056
rect 3844 10004 3850 10056
rect 4177 10053 4205 10084
rect 4162 10047 4220 10053
rect 3896 10016 4108 10044
rect 2225 9979 2283 9985
rect 2225 9945 2237 9979
rect 2271 9976 2283 9979
rect 2685 9979 2743 9985
rect 2685 9976 2697 9979
rect 2271 9948 2697 9976
rect 2271 9945 2283 9948
rect 2225 9939 2283 9945
rect 2685 9945 2697 9948
rect 2731 9945 2743 9979
rect 2685 9939 2743 9945
rect 2777 9979 2835 9985
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 3896 9976 3924 10016
rect 4080 9985 4108 10016
rect 4162 10013 4174 10047
rect 4208 10013 4220 10047
rect 4162 10007 4220 10013
rect 4798 10004 4804 10056
rect 4856 10004 4862 10056
rect 5276 10053 5304 10084
rect 5537 10115 5595 10121
rect 5537 10081 5549 10115
rect 5583 10081 5595 10115
rect 5537 10075 5595 10081
rect 5810 10072 5816 10124
rect 5868 10072 5874 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 5960 10084 8156 10112
rect 5960 10072 5966 10084
rect 8128 10056 8156 10084
rect 5221 10047 5304 10053
rect 4908 10016 5120 10044
rect 2823 9948 3924 9976
rect 3973 9979 4031 9985
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 3973 9945 3985 9979
rect 4019 9945 4031 9979
rect 3973 9939 4031 9945
rect 4065 9979 4123 9985
rect 4065 9945 4077 9979
rect 4111 9976 4123 9979
rect 4246 9976 4252 9988
rect 4111 9948 4252 9976
rect 4111 9945 4123 9948
rect 4065 9939 4123 9945
rect 2038 9868 2044 9920
rect 2096 9908 2102 9920
rect 2240 9908 2268 9939
rect 2096 9880 2268 9908
rect 2700 9908 2728 9939
rect 3988 9908 4016 9939
rect 4246 9936 4252 9948
rect 4304 9976 4310 9988
rect 4614 9976 4620 9988
rect 4304 9948 4620 9976
rect 4304 9936 4310 9948
rect 4614 9936 4620 9948
rect 4672 9976 4678 9988
rect 4908 9976 4936 10016
rect 5092 9985 5120 10016
rect 5221 10013 5233 10047
rect 5267 10016 5304 10047
rect 5267 10013 5279 10016
rect 5221 10007 5279 10013
rect 7190 10004 7196 10056
rect 7248 10044 7254 10056
rect 7561 10047 7619 10053
rect 7561 10044 7573 10047
rect 7248 10016 7573 10044
rect 7248 10004 7254 10016
rect 7561 10013 7573 10016
rect 7607 10013 7619 10047
rect 7561 10007 7619 10013
rect 7650 10004 7656 10056
rect 7708 10004 7714 10056
rect 7834 10004 7840 10056
rect 7892 10004 7898 10056
rect 8110 10004 8116 10056
rect 8168 10004 8174 10056
rect 8225 10053 8253 10152
rect 8389 10149 8401 10183
rect 8435 10180 8447 10183
rect 8570 10180 8576 10192
rect 8435 10152 8576 10180
rect 8435 10149 8447 10152
rect 8389 10143 8447 10149
rect 8570 10140 8576 10152
rect 8628 10140 8634 10192
rect 9766 10072 9772 10124
rect 9824 10112 9830 10124
rect 9824 10084 10824 10112
rect 9824 10072 9830 10084
rect 8210 10047 8268 10053
rect 8210 10013 8222 10047
rect 8256 10013 8268 10047
rect 8210 10007 8268 10013
rect 4672 9948 4936 9976
rect 4985 9979 5043 9985
rect 4672 9936 4678 9948
rect 4985 9945 4997 9979
rect 5031 9945 5043 9979
rect 4985 9939 5043 9945
rect 5077 9979 5135 9985
rect 5077 9945 5089 9979
rect 5123 9976 5135 9979
rect 5902 9976 5908 9988
rect 5123 9948 5908 9976
rect 5123 9945 5135 9948
rect 5077 9939 5135 9945
rect 5000 9908 5028 9939
rect 5902 9936 5908 9948
rect 5960 9936 5966 9988
rect 6270 9936 6276 9988
rect 6328 9936 6334 9988
rect 8021 9979 8079 9985
rect 8021 9945 8033 9979
rect 8067 9945 8079 9979
rect 8021 9939 8079 9945
rect 6638 9908 6644 9920
rect 2700 9880 6644 9908
rect 2096 9868 2102 9880
rect 6638 9868 6644 9880
rect 6696 9908 6702 9920
rect 7098 9908 7104 9920
rect 6696 9880 7104 9908
rect 6696 9868 6702 9880
rect 7098 9868 7104 9880
rect 7156 9908 7162 9920
rect 8036 9908 8064 9939
rect 8754 9936 8760 9988
rect 8812 9976 8818 9988
rect 8941 9979 8999 9985
rect 8941 9976 8953 9979
rect 8812 9948 8953 9976
rect 8812 9936 8818 9948
rect 8941 9945 8953 9948
rect 8987 9945 8999 9979
rect 8941 9939 8999 9945
rect 9490 9936 9496 9988
rect 9548 9976 9554 9988
rect 9876 9976 9904 10030
rect 10502 10004 10508 10056
rect 10560 10004 10566 10056
rect 10796 9988 10824 10084
rect 11514 10072 11520 10124
rect 11572 10072 11578 10124
rect 11793 10115 11851 10121
rect 11793 10081 11805 10115
rect 11839 10112 11851 10115
rect 11839 10084 13676 10112
rect 11839 10081 11851 10084
rect 11793 10075 11851 10081
rect 10870 10004 10876 10056
rect 10928 10053 10934 10056
rect 10928 10044 10936 10053
rect 10928 10016 10973 10044
rect 10928 10007 10936 10016
rect 10928 10004 10934 10007
rect 10226 9976 10232 9988
rect 9548 9948 10232 9976
rect 9548 9936 9554 9948
rect 10226 9936 10232 9948
rect 10284 9976 10290 9988
rect 10689 9979 10747 9985
rect 10689 9976 10701 9979
rect 10284 9948 10701 9976
rect 10284 9936 10290 9948
rect 10689 9945 10701 9948
rect 10735 9945 10747 9979
rect 10689 9939 10747 9945
rect 10778 9936 10784 9988
rect 10836 9936 10842 9988
rect 13078 9976 13084 9988
rect 13018 9948 13084 9976
rect 13078 9936 13084 9948
rect 13136 9976 13142 9988
rect 13262 9976 13268 9988
rect 13136 9948 13268 9976
rect 13136 9936 13142 9948
rect 13262 9936 13268 9948
rect 13320 9936 13326 9988
rect 13538 9936 13544 9988
rect 13596 9936 13602 9988
rect 13648 9976 13676 10084
rect 13740 10053 13768 10220
rect 15654 10208 15660 10220
rect 15712 10208 15718 10260
rect 15746 10208 15752 10260
rect 15804 10248 15810 10260
rect 16025 10251 16083 10257
rect 16025 10248 16037 10251
rect 15804 10220 16037 10248
rect 15804 10208 15810 10220
rect 16025 10217 16037 10220
rect 16071 10217 16083 10251
rect 16025 10211 16083 10217
rect 17954 10208 17960 10260
rect 18012 10208 18018 10260
rect 15102 10112 15108 10124
rect 13832 10084 15108 10112
rect 13725 10047 13783 10053
rect 13725 10013 13737 10047
rect 13771 10013 13783 10047
rect 13725 10007 13783 10013
rect 13832 9976 13860 10084
rect 15102 10072 15108 10084
rect 15160 10072 15166 10124
rect 16482 10072 16488 10124
rect 16540 10072 16546 10124
rect 13906 10004 13912 10056
rect 13964 10004 13970 10056
rect 14277 10047 14335 10053
rect 14277 10013 14289 10047
rect 14323 10013 14335 10047
rect 14277 10007 14335 10013
rect 13648 9948 13860 9976
rect 7156 9880 8064 9908
rect 11074 9911 11132 9917
rect 7156 9868 7162 9880
rect 11074 9877 11086 9911
rect 11120 9908 11132 9911
rect 13170 9908 13176 9920
rect 11120 9880 13176 9908
rect 11120 9877 11132 9880
rect 11074 9871 11132 9877
rect 13170 9868 13176 9880
rect 13228 9868 13234 9920
rect 14292 9908 14320 10007
rect 15930 10004 15936 10056
rect 15988 10044 15994 10056
rect 16209 10047 16267 10053
rect 16209 10044 16221 10047
rect 15988 10016 16221 10044
rect 15988 10004 15994 10016
rect 16209 10013 16221 10016
rect 16255 10013 16267 10047
rect 16209 10007 16267 10013
rect 14553 9979 14611 9985
rect 14553 9945 14565 9979
rect 14599 9976 14611 9979
rect 14826 9976 14832 9988
rect 14599 9948 14832 9976
rect 14599 9945 14611 9948
rect 14553 9939 14611 9945
rect 14826 9936 14832 9948
rect 14884 9936 14890 9988
rect 15010 9936 15016 9988
rect 15068 9936 15074 9988
rect 16574 9936 16580 9988
rect 16632 9976 16638 9988
rect 16632 9948 16974 9976
rect 16632 9936 16638 9948
rect 15470 9908 15476 9920
rect 14292 9880 15476 9908
rect 15470 9868 15476 9880
rect 15528 9868 15534 9920
rect 1104 9818 22816 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 22816 9818
rect 1104 9744 22816 9766
rect 2498 9704 2504 9716
rect 1964 9676 2504 9704
rect 1964 9645 1992 9676
rect 2498 9664 2504 9676
rect 2556 9664 2562 9716
rect 6270 9664 6276 9716
rect 6328 9704 6334 9716
rect 9398 9704 9404 9716
rect 6328 9676 9404 9704
rect 6328 9664 6334 9676
rect 1949 9639 2007 9645
rect 1949 9605 1961 9639
rect 1995 9605 2007 9639
rect 5721 9639 5779 9645
rect 5721 9636 5733 9639
rect 1949 9599 2007 9605
rect 4448 9608 5733 9636
rect 2038 9528 2044 9580
rect 2096 9528 2102 9580
rect 3418 9528 3424 9580
rect 3476 9528 3482 9580
rect 4157 9571 4215 9577
rect 4157 9537 4169 9571
rect 4203 9568 4215 9571
rect 4246 9568 4252 9580
rect 4203 9540 4252 9568
rect 4203 9537 4215 9540
rect 4157 9531 4215 9537
rect 4246 9528 4252 9540
rect 4304 9528 4310 9580
rect 4448 9577 4476 9608
rect 5721 9605 5733 9608
rect 5767 9636 5779 9639
rect 6638 9636 6644 9648
rect 5767 9608 6644 9636
rect 5767 9605 5779 9608
rect 5721 9599 5779 9605
rect 6638 9596 6644 9608
rect 6696 9596 6702 9648
rect 7944 9636 7972 9676
rect 9398 9664 9404 9676
rect 9456 9704 9462 9716
rect 13078 9704 13084 9716
rect 9456 9676 13084 9704
rect 9456 9664 9462 9676
rect 7866 9608 7972 9636
rect 8754 9596 8760 9648
rect 8812 9596 8818 9648
rect 10152 9636 10180 9676
rect 13078 9664 13084 9676
rect 13136 9664 13142 9716
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 15286 9704 15292 9716
rect 13228 9676 15292 9704
rect 13228 9664 13234 9676
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 9982 9608 10180 9636
rect 10226 9596 10232 9648
rect 10284 9636 10290 9648
rect 12066 9636 12072 9648
rect 10284 9608 12072 9636
rect 10284 9596 10290 9608
rect 12066 9596 12072 9608
rect 12124 9636 12130 9648
rect 12124 9608 12296 9636
rect 12124 9596 12130 9608
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9537 4491 9571
rect 4433 9531 4491 9537
rect 4798 9528 4804 9580
rect 4856 9568 4862 9580
rect 5442 9568 5448 9580
rect 4856 9540 5448 9568
rect 4856 9528 4862 9540
rect 5442 9528 5448 9540
rect 5500 9568 5506 9580
rect 5537 9571 5595 9577
rect 5537 9568 5549 9571
rect 5500 9540 5549 9568
rect 5500 9528 5506 9540
rect 5537 9537 5549 9540
rect 5583 9537 5595 9571
rect 5537 9531 5595 9537
rect 5810 9528 5816 9580
rect 5868 9528 5874 9580
rect 5994 9577 6000 9580
rect 5957 9571 6000 9577
rect 5957 9537 5969 9571
rect 5957 9531 6000 9537
rect 5994 9528 6000 9531
rect 6052 9528 6058 9580
rect 8478 9528 8484 9580
rect 8536 9528 8542 9580
rect 10042 9528 10048 9580
rect 10100 9568 10106 9580
rect 10413 9571 10471 9577
rect 10413 9568 10425 9571
rect 10100 9540 10425 9568
rect 10100 9528 10106 9540
rect 10413 9537 10425 9540
rect 10459 9568 10471 9571
rect 10594 9568 10600 9580
rect 10459 9540 10600 9568
rect 10459 9537 10471 9540
rect 10413 9531 10471 9537
rect 10594 9528 10600 9540
rect 10652 9528 10658 9580
rect 10778 9528 10784 9580
rect 10836 9568 10842 9580
rect 11517 9571 11575 9577
rect 10836 9540 11284 9568
rect 10836 9528 10842 9540
rect 2314 9460 2320 9512
rect 2372 9460 2378 9512
rect 6365 9503 6423 9509
rect 6365 9500 6377 9503
rect 6104 9472 6377 9500
rect 1302 9392 1308 9444
rect 1360 9432 1366 9444
rect 1581 9435 1639 9441
rect 1581 9432 1593 9435
rect 1360 9404 1593 9432
rect 1360 9392 1366 9404
rect 1581 9401 1593 9404
rect 1627 9401 1639 9435
rect 1581 9395 1639 9401
rect 3694 9392 3700 9444
rect 3752 9432 3758 9444
rect 6104 9441 6132 9472
rect 6365 9469 6377 9472
rect 6411 9469 6423 9503
rect 6365 9463 6423 9469
rect 6641 9503 6699 9509
rect 6641 9469 6653 9503
rect 6687 9500 6699 9503
rect 7190 9500 7196 9512
rect 6687 9472 7196 9500
rect 6687 9469 6699 9472
rect 6641 9463 6699 9469
rect 7190 9460 7196 9472
rect 7248 9460 7254 9512
rect 7650 9460 7656 9512
rect 7708 9500 7714 9512
rect 8113 9503 8171 9509
rect 8113 9500 8125 9503
rect 7708 9472 8125 9500
rect 7708 9460 7714 9472
rect 8113 9469 8125 9472
rect 8159 9500 8171 9503
rect 9766 9500 9772 9512
rect 8159 9472 9772 9500
rect 8159 9469 8171 9472
rect 8113 9463 8171 9469
rect 9766 9460 9772 9472
rect 9824 9460 9830 9512
rect 10226 9460 10232 9512
rect 10284 9460 10290 9512
rect 10962 9460 10968 9512
rect 11020 9500 11026 9512
rect 11149 9503 11207 9509
rect 11149 9500 11161 9503
rect 11020 9472 11161 9500
rect 11020 9460 11026 9472
rect 11149 9469 11161 9472
rect 11195 9469 11207 9503
rect 11256 9500 11284 9540
rect 11517 9537 11529 9571
rect 11563 9568 11575 9571
rect 11606 9568 11612 9580
rect 11563 9540 11612 9568
rect 11563 9537 11575 9540
rect 11517 9531 11575 9537
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 11698 9528 11704 9580
rect 11756 9528 11762 9580
rect 11790 9528 11796 9580
rect 11848 9528 11854 9580
rect 11974 9577 11980 9580
rect 11937 9571 11980 9577
rect 11937 9537 11949 9571
rect 11937 9531 11980 9537
rect 11974 9528 11980 9531
rect 12032 9528 12038 9580
rect 12268 9577 12296 9608
rect 13188 9577 13216 9664
rect 13449 9639 13507 9645
rect 13449 9605 13461 9639
rect 13495 9636 13507 9639
rect 13538 9636 13544 9648
rect 13495 9608 13544 9636
rect 13495 9605 13507 9608
rect 13449 9599 13507 9605
rect 13538 9596 13544 9608
rect 13596 9596 13602 9648
rect 13906 9596 13912 9648
rect 13964 9596 13970 9648
rect 15470 9596 15476 9648
rect 15528 9596 15534 9648
rect 16574 9596 16580 9648
rect 16632 9636 16638 9648
rect 17402 9636 17408 9648
rect 16632 9608 17408 9636
rect 16632 9596 16638 9608
rect 17402 9596 17408 9608
rect 17460 9636 17466 9648
rect 17460 9608 17986 9636
rect 17460 9596 17466 9608
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9537 12311 9571
rect 12253 9531 12311 9537
rect 12437 9571 12495 9577
rect 12437 9537 12449 9571
rect 12483 9568 12495 9571
rect 13173 9571 13231 9577
rect 12483 9540 12517 9568
rect 12483 9537 12495 9540
rect 12437 9531 12495 9537
rect 13173 9537 13185 9571
rect 13219 9537 13231 9571
rect 15105 9571 15163 9577
rect 15105 9568 15117 9571
rect 13173 9531 13231 9537
rect 14660 9540 15117 9568
rect 12452 9500 12480 9531
rect 12618 9500 12624 9512
rect 11256 9472 12624 9500
rect 11149 9463 11207 9469
rect 12618 9460 12624 9472
rect 12676 9460 12682 9512
rect 12805 9503 12863 9509
rect 12805 9469 12817 9503
rect 12851 9500 12863 9503
rect 13078 9500 13084 9512
rect 12851 9472 13084 9500
rect 12851 9469 12863 9472
rect 12805 9463 12863 9469
rect 13078 9460 13084 9472
rect 13136 9460 13142 9512
rect 13814 9460 13820 9512
rect 13872 9500 13878 9512
rect 14660 9500 14688 9540
rect 15105 9537 15117 9540
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 15286 9528 15292 9580
rect 15344 9568 15350 9580
rect 15381 9571 15439 9577
rect 15381 9568 15393 9571
rect 15344 9540 15393 9568
rect 15344 9528 15350 9540
rect 15381 9537 15393 9540
rect 15427 9537 15439 9571
rect 16669 9571 16727 9577
rect 16669 9568 16681 9571
rect 15381 9531 15439 9537
rect 15948 9540 16681 9568
rect 13872 9472 14688 9500
rect 13872 9460 13878 9472
rect 14826 9460 14832 9512
rect 14884 9500 14890 9512
rect 14921 9503 14979 9509
rect 14921 9500 14933 9503
rect 14884 9472 14933 9500
rect 14884 9460 14890 9472
rect 14921 9469 14933 9472
rect 14967 9469 14979 9503
rect 14921 9463 14979 9469
rect 4341 9435 4399 9441
rect 4341 9432 4353 9435
rect 3752 9404 4353 9432
rect 3752 9392 3758 9404
rect 4341 9401 4353 9404
rect 4387 9401 4399 9435
rect 4341 9395 4399 9401
rect 6089 9435 6147 9441
rect 6089 9401 6101 9435
rect 6135 9401 6147 9435
rect 6089 9395 6147 9401
rect 11054 9392 11060 9444
rect 11112 9432 11118 9444
rect 12713 9435 12771 9441
rect 12713 9432 12725 9435
rect 11112 9404 12725 9432
rect 11112 9392 11118 9404
rect 12713 9401 12725 9404
rect 12759 9401 12771 9435
rect 12713 9395 12771 9401
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 15289 9435 15347 9441
rect 15289 9432 15301 9435
rect 15068 9404 15301 9432
rect 15068 9392 15074 9404
rect 15289 9401 15301 9404
rect 15335 9401 15347 9435
rect 15289 9395 15347 9401
rect 15562 9392 15568 9444
rect 15620 9432 15626 9444
rect 15948 9441 15976 9540
rect 16669 9537 16681 9540
rect 16715 9537 16727 9571
rect 16669 9531 16727 9537
rect 16853 9571 16911 9577
rect 16853 9537 16865 9571
rect 16899 9537 16911 9571
rect 16853 9531 16911 9537
rect 16301 9503 16359 9509
rect 16301 9469 16313 9503
rect 16347 9469 16359 9503
rect 16301 9463 16359 9469
rect 15933 9435 15991 9441
rect 15933 9432 15945 9435
rect 15620 9404 15945 9432
rect 15620 9392 15626 9404
rect 15933 9401 15945 9404
rect 15979 9401 15991 9435
rect 15933 9395 15991 9401
rect 1486 9324 1492 9376
rect 1544 9324 1550 9376
rect 3789 9367 3847 9373
rect 3789 9333 3801 9367
rect 3835 9364 3847 9367
rect 3878 9364 3884 9376
rect 3835 9336 3884 9364
rect 3835 9333 3847 9336
rect 3789 9327 3847 9333
rect 3878 9324 3884 9336
rect 3936 9324 3942 9376
rect 3970 9324 3976 9376
rect 4028 9364 4034 9376
rect 4065 9367 4123 9373
rect 4065 9364 4077 9367
rect 4028 9336 4077 9364
rect 4028 9324 4034 9336
rect 4065 9333 4077 9336
rect 4111 9333 4123 9367
rect 4065 9327 4123 9333
rect 6822 9324 6828 9376
rect 6880 9364 6886 9376
rect 10502 9364 10508 9376
rect 6880 9336 10508 9364
rect 6880 9324 6886 9336
rect 10502 9324 10508 9336
rect 10560 9364 10566 9376
rect 11146 9364 11152 9376
rect 10560 9336 11152 9364
rect 10560 9324 10566 9336
rect 11146 9324 11152 9336
rect 11204 9324 11210 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 12069 9367 12127 9373
rect 12069 9364 12081 9367
rect 11388 9336 12081 9364
rect 11388 9324 11394 9336
rect 12069 9333 12081 9336
rect 12115 9333 12127 9367
rect 12069 9327 12127 9333
rect 15838 9324 15844 9376
rect 15896 9324 15902 9376
rect 16022 9324 16028 9376
rect 16080 9364 16086 9376
rect 16316 9364 16344 9463
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 16868 9500 16896 9531
rect 16540 9472 16896 9500
rect 16540 9460 16546 9472
rect 18414 9460 18420 9512
rect 18472 9500 18478 9512
rect 19153 9503 19211 9509
rect 19153 9500 19165 9503
rect 18472 9472 19165 9500
rect 18472 9460 18478 9472
rect 19153 9469 19165 9472
rect 19199 9469 19211 9503
rect 19153 9463 19211 9469
rect 19426 9460 19432 9512
rect 19484 9460 19490 9512
rect 16942 9392 16948 9444
rect 17000 9392 17006 9444
rect 17681 9367 17739 9373
rect 17681 9364 17693 9367
rect 16080 9336 17693 9364
rect 16080 9324 16086 9336
rect 17681 9333 17693 9336
rect 17727 9333 17739 9367
rect 17681 9327 17739 9333
rect 1104 9274 22816 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 20214 9274
rect 20266 9222 20278 9274
rect 20330 9222 20342 9274
rect 20394 9222 20406 9274
rect 20458 9222 20470 9274
rect 20522 9222 22816 9274
rect 1104 9200 22816 9222
rect 1486 9120 1492 9172
rect 1544 9160 1550 9172
rect 2022 9163 2080 9169
rect 2022 9160 2034 9163
rect 1544 9132 2034 9160
rect 1544 9120 1550 9132
rect 2022 9129 2034 9132
rect 2068 9129 2080 9163
rect 2022 9123 2080 9129
rect 5721 9163 5779 9169
rect 5721 9129 5733 9163
rect 5767 9160 5779 9163
rect 5994 9160 6000 9172
rect 5767 9132 6000 9160
rect 5767 9129 5779 9132
rect 5721 9123 5779 9129
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 11606 9160 11612 9172
rect 6512 9132 11612 9160
rect 6512 9120 6518 9132
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 11698 9120 11704 9172
rect 11756 9160 11762 9172
rect 13814 9160 13820 9172
rect 11756 9132 13820 9160
rect 11756 9120 11762 9132
rect 13814 9120 13820 9132
rect 13872 9120 13878 9172
rect 15010 9120 15016 9172
rect 15068 9160 15074 9172
rect 16390 9160 16396 9172
rect 15068 9132 16396 9160
rect 15068 9120 15074 9132
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 17681 9163 17739 9169
rect 17681 9129 17693 9163
rect 17727 9160 17739 9163
rect 19426 9160 19432 9172
rect 17727 9132 19432 9160
rect 17727 9129 17739 9132
rect 17681 9123 17739 9129
rect 19426 9120 19432 9132
rect 19484 9120 19490 9172
rect 3418 9092 3424 9104
rect 3160 9064 3424 9092
rect 1765 9027 1823 9033
rect 1765 8993 1777 9027
rect 1811 9024 1823 9027
rect 2130 9024 2136 9036
rect 1811 8996 2136 9024
rect 1811 8993 1823 8996
rect 1765 8987 1823 8993
rect 2130 8984 2136 8996
rect 2188 8984 2194 9036
rect 3160 8942 3188 9064
rect 3418 9052 3424 9064
rect 3476 9092 3482 9104
rect 6549 9095 6607 9101
rect 3476 9064 4108 9092
rect 3476 9052 3482 9064
rect 3970 8984 3976 9036
rect 4028 8984 4034 9036
rect 4080 9024 4108 9064
rect 6549 9061 6561 9095
rect 6595 9092 6607 9095
rect 6595 9064 6684 9092
rect 6595 9061 6607 9064
rect 6549 9055 6607 9061
rect 4080 8996 5488 9024
rect 4249 8891 4307 8897
rect 4249 8888 4261 8891
rect 3528 8860 4261 8888
rect 3528 8829 3556 8860
rect 4249 8857 4261 8860
rect 4295 8857 4307 8891
rect 5460 8888 5488 8996
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 6549 8959 6607 8965
rect 6549 8956 6561 8959
rect 6512 8928 6561 8956
rect 6512 8916 6518 8928
rect 6549 8925 6561 8928
rect 6595 8925 6607 8959
rect 6549 8919 6607 8925
rect 5534 8888 5540 8900
rect 5460 8874 5540 8888
rect 5474 8860 5540 8874
rect 4249 8851 4307 8857
rect 5534 8848 5540 8860
rect 5592 8888 5598 8900
rect 6656 8888 6684 9064
rect 11256 9064 11468 9092
rect 6917 9027 6975 9033
rect 6917 8993 6929 9027
rect 6963 9024 6975 9027
rect 7650 9024 7656 9036
rect 6963 8996 7656 9024
rect 6963 8993 6975 8996
rect 6917 8987 6975 8993
rect 7650 8984 7656 8996
rect 7708 8984 7714 9036
rect 8665 9027 8723 9033
rect 8665 8993 8677 9027
rect 8711 9024 8723 9027
rect 9217 9027 9275 9033
rect 9217 9024 9229 9027
rect 8711 8996 9229 9024
rect 8711 8993 8723 8996
rect 8665 8987 8723 8993
rect 9217 8993 9229 8996
rect 9263 8993 9275 9027
rect 9217 8987 9275 8993
rect 6822 8916 6828 8968
rect 6880 8916 6886 8968
rect 8938 8916 8944 8968
rect 8996 8916 9002 8968
rect 10962 8956 10968 8968
rect 10350 8942 10968 8956
rect 10336 8928 10968 8942
rect 7193 8891 7251 8897
rect 7193 8888 7205 8891
rect 5592 8860 6316 8888
rect 6656 8860 7205 8888
rect 5592 8848 5598 8860
rect 3513 8823 3571 8829
rect 3513 8789 3525 8823
rect 3559 8789 3571 8823
rect 6288 8820 6316 8860
rect 7193 8857 7205 8860
rect 7239 8857 7251 8891
rect 8418 8860 8524 8888
rect 7193 8851 7251 8857
rect 8496 8820 8524 8860
rect 8846 8820 8852 8832
rect 6288 8792 8852 8820
rect 3513 8783 3571 8789
rect 8846 8780 8852 8792
rect 8904 8820 8910 8832
rect 10336 8820 10364 8928
rect 10962 8916 10968 8928
rect 11020 8916 11026 8968
rect 11054 8916 11060 8968
rect 11112 8916 11118 8968
rect 11256 8965 11284 9064
rect 11330 8984 11336 9036
rect 11388 8984 11394 9036
rect 11440 9024 11468 9064
rect 13078 9052 13084 9104
rect 13136 9092 13142 9104
rect 13136 9064 14780 9092
rect 13136 9052 13142 9064
rect 12802 9024 12808 9036
rect 11440 8996 12808 9024
rect 12802 8984 12808 8996
rect 12860 9024 12866 9036
rect 14645 9027 14703 9033
rect 14645 9024 14657 9027
rect 12860 8996 14657 9024
rect 12860 8984 12866 8996
rect 14645 8993 14657 8996
rect 14691 8993 14703 9027
rect 14752 9024 14780 9064
rect 14752 8996 17264 9024
rect 14645 8987 14703 8993
rect 17236 8968 17264 8996
rect 11241 8959 11299 8965
rect 11241 8925 11253 8959
rect 11287 8925 11299 8959
rect 13262 8956 13268 8968
rect 12742 8928 13268 8956
rect 11241 8919 11299 8925
rect 13262 8916 13268 8928
rect 13320 8956 13326 8968
rect 13538 8956 13544 8968
rect 13320 8928 13544 8956
rect 13320 8916 13326 8928
rect 13538 8916 13544 8928
rect 13596 8916 13602 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15381 8959 15439 8965
rect 15381 8956 15393 8959
rect 14976 8928 15393 8956
rect 14976 8916 14982 8928
rect 15381 8925 15393 8928
rect 15427 8925 15439 8959
rect 15381 8919 15439 8925
rect 15470 8916 15476 8968
rect 15528 8956 15534 8968
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 15528 8928 15669 8956
rect 15528 8916 15534 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17589 8959 17647 8965
rect 17589 8956 17601 8959
rect 17276 8928 17601 8956
rect 17276 8916 17282 8928
rect 17589 8925 17601 8928
rect 17635 8925 17647 8959
rect 17589 8919 17647 8925
rect 11609 8891 11667 8897
rect 11609 8888 11621 8891
rect 11164 8860 11621 8888
rect 8904 8792 10364 8820
rect 8904 8780 8910 8792
rect 10686 8780 10692 8832
rect 10744 8780 10750 8832
rect 11164 8829 11192 8860
rect 11609 8857 11621 8860
rect 11655 8857 11667 8891
rect 15562 8888 15568 8900
rect 11609 8851 11667 8857
rect 13188 8860 15568 8888
rect 11149 8823 11207 8829
rect 11149 8789 11161 8823
rect 11195 8789 11207 8823
rect 11149 8783 11207 8789
rect 11698 8780 11704 8832
rect 11756 8820 11762 8832
rect 13188 8820 13216 8860
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 15838 8848 15844 8900
rect 15896 8888 15902 8900
rect 15933 8891 15991 8897
rect 15933 8888 15945 8891
rect 15896 8860 15945 8888
rect 15896 8848 15902 8860
rect 15933 8857 15945 8860
rect 15979 8857 15991 8891
rect 15933 8851 15991 8857
rect 16390 8848 16396 8900
rect 16448 8848 16454 8900
rect 11756 8792 13216 8820
rect 11756 8780 11762 8792
rect 13262 8780 13268 8832
rect 13320 8820 13326 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13320 8792 14105 8820
rect 13320 8780 13326 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14093 8783 14151 8789
rect 15194 8780 15200 8832
rect 15252 8820 15258 8832
rect 17405 8823 17463 8829
rect 17405 8820 17417 8823
rect 15252 8792 17417 8820
rect 15252 8780 15258 8792
rect 17405 8789 17417 8792
rect 17451 8789 17463 8823
rect 17405 8783 17463 8789
rect 1104 8730 22816 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 22816 8730
rect 1104 8656 22816 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 2593 8619 2651 8625
rect 2593 8616 2605 8619
rect 2372 8588 2605 8616
rect 2372 8576 2378 8588
rect 2593 8585 2605 8588
rect 2639 8585 2651 8619
rect 2593 8579 2651 8585
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 9858 8616 9864 8628
rect 9048 8588 9864 8616
rect 1486 8508 1492 8560
rect 1544 8548 1550 8560
rect 3145 8551 3203 8557
rect 3145 8548 3157 8551
rect 1544 8520 3157 8548
rect 1544 8508 1550 8520
rect 3145 8517 3157 8520
rect 3191 8517 3203 8551
rect 3145 8511 3203 8517
rect 3878 8508 3884 8560
rect 3936 8548 3942 8560
rect 3973 8551 4031 8557
rect 3973 8548 3985 8551
rect 3936 8520 3985 8548
rect 3936 8508 3942 8520
rect 3973 8517 3985 8520
rect 4019 8517 4031 8551
rect 5534 8548 5540 8560
rect 5198 8520 5540 8548
rect 3973 8511 4031 8517
rect 5534 8508 5540 8520
rect 5592 8508 5598 8560
rect 9048 8548 9076 8588
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10686 8576 10692 8628
rect 10744 8616 10750 8628
rect 11977 8619 12035 8625
rect 10744 8588 11560 8616
rect 10744 8576 10750 8588
rect 9766 8548 9772 8560
rect 7866 8520 9076 8548
rect 9140 8520 9772 8548
rect 1946 8440 1952 8492
rect 2004 8489 2010 8492
rect 2004 8483 2047 8489
rect 2035 8449 2047 8483
rect 2004 8443 2047 8449
rect 2004 8440 2010 8443
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 2225 8483 2283 8489
rect 2225 8449 2237 8483
rect 2271 8480 2283 8483
rect 2314 8480 2320 8492
rect 2271 8452 2320 8480
rect 2271 8449 2283 8452
rect 2225 8443 2283 8449
rect 2314 8440 2320 8452
rect 2372 8440 2378 8492
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 2501 8483 2559 8489
rect 2501 8449 2513 8483
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 1118 8372 1124 8424
rect 1176 8412 1182 8424
rect 2424 8412 2452 8443
rect 1176 8384 2452 8412
rect 1176 8372 1182 8384
rect 1302 8304 1308 8356
rect 1360 8344 1366 8356
rect 1360 8316 1716 8344
rect 1360 8304 1366 8316
rect 1688 8276 1716 8316
rect 1762 8304 1768 8356
rect 1820 8344 1826 8356
rect 1857 8347 1915 8353
rect 1857 8344 1869 8347
rect 1820 8316 1869 8344
rect 1820 8304 1826 8316
rect 1857 8313 1869 8316
rect 1903 8313 1915 8347
rect 2516 8344 2544 8443
rect 2682 8440 2688 8492
rect 2740 8440 2746 8492
rect 2961 8483 3019 8489
rect 2961 8449 2973 8483
rect 3007 8480 3019 8483
rect 3050 8480 3056 8492
rect 3007 8452 3056 8480
rect 3007 8449 3019 8452
rect 2961 8443 3019 8449
rect 3050 8440 3056 8452
rect 3108 8440 3114 8492
rect 3234 8440 3240 8492
rect 3292 8440 3298 8492
rect 3381 8483 3439 8489
rect 3381 8449 3393 8483
rect 3427 8480 3439 8483
rect 3602 8480 3608 8492
rect 3427 8452 3608 8480
rect 3427 8449 3439 8452
rect 3381 8443 3439 8449
rect 3602 8440 3608 8452
rect 3660 8440 3666 8492
rect 3694 8440 3700 8492
rect 3752 8440 3758 8492
rect 8938 8440 8944 8492
rect 8996 8480 9002 8492
rect 9140 8489 9168 8520
rect 9766 8508 9772 8520
rect 9824 8508 9830 8560
rect 9876 8548 9904 8576
rect 11532 8557 11560 8588
rect 11977 8585 11989 8619
rect 12023 8585 12035 8619
rect 12618 8616 12624 8628
rect 11977 8579 12035 8585
rect 12176 8588 12624 8616
rect 11517 8551 11575 8557
rect 9876 8520 10258 8548
rect 11517 8517 11529 8551
rect 11563 8517 11575 8551
rect 11517 8511 11575 8517
rect 9033 8483 9091 8489
rect 9033 8480 9045 8483
rect 8996 8452 9045 8480
rect 8996 8440 9002 8452
rect 9033 8449 9045 8452
rect 9079 8449 9091 8483
rect 9033 8443 9091 8449
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 11992 8480 12020 8579
rect 12176 8557 12204 8588
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13078 8576 13084 8628
rect 13136 8576 13142 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 15470 8616 15476 8628
rect 14783 8588 15476 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 15470 8576 15476 8588
rect 15528 8616 15534 8628
rect 15528 8588 16344 8616
rect 15528 8576 15534 8588
rect 12161 8551 12219 8557
rect 12161 8517 12173 8551
rect 12207 8517 12219 8551
rect 12161 8511 12219 8517
rect 12345 8551 12403 8557
rect 12345 8517 12357 8551
rect 12391 8548 12403 8551
rect 13096 8548 13124 8576
rect 12391 8520 13124 8548
rect 12391 8517 12403 8520
rect 12345 8511 12403 8517
rect 13262 8508 13268 8560
rect 13320 8508 13326 8560
rect 13538 8508 13544 8560
rect 13596 8548 13602 8560
rect 13596 8520 13754 8548
rect 13596 8508 13602 8520
rect 16022 8508 16028 8560
rect 16080 8548 16086 8560
rect 16316 8557 16344 8588
rect 18414 8576 18420 8628
rect 18472 8576 18478 8628
rect 16209 8551 16267 8557
rect 16209 8548 16221 8551
rect 16080 8520 16221 8548
rect 16080 8508 16086 8520
rect 16209 8517 16221 8520
rect 16255 8517 16267 8551
rect 16209 8511 16267 8517
rect 16301 8551 16359 8557
rect 16301 8517 16313 8551
rect 16347 8517 16359 8551
rect 17218 8548 17224 8560
rect 16301 8511 16359 8517
rect 16684 8520 17224 8548
rect 10980 8452 12020 8480
rect 6362 8372 6368 8424
rect 6420 8372 6426 8424
rect 6641 8415 6699 8421
rect 6641 8381 6653 8415
rect 6687 8412 6699 8415
rect 6730 8412 6736 8424
rect 6687 8384 6736 8412
rect 6687 8381 6699 8384
rect 6641 8375 6699 8381
rect 6730 8372 6736 8384
rect 6788 8372 6794 8424
rect 8294 8372 8300 8424
rect 8352 8372 8358 8424
rect 9769 8415 9827 8421
rect 9769 8381 9781 8415
rect 9815 8412 9827 8415
rect 10980 8412 11008 8452
rect 12066 8440 12072 8492
rect 12124 8480 12130 8492
rect 12713 8483 12771 8489
rect 12713 8480 12725 8483
rect 12124 8452 12725 8480
rect 12124 8440 12130 8452
rect 9815 8384 11008 8412
rect 9815 8381 9827 8384
rect 9769 8375 9827 8381
rect 11606 8372 11612 8424
rect 11664 8412 11670 8424
rect 11664 8384 11836 8412
rect 11664 8372 11670 8384
rect 1857 8307 1915 8313
rect 1964 8316 2544 8344
rect 3513 8347 3571 8353
rect 1964 8276 1992 8316
rect 3513 8313 3525 8347
rect 3559 8344 3571 8347
rect 3694 8344 3700 8356
rect 3559 8316 3700 8344
rect 3559 8313 3571 8316
rect 3513 8307 3571 8313
rect 3694 8304 3700 8316
rect 3752 8304 3758 8356
rect 8573 8347 8631 8353
rect 8573 8344 8585 8347
rect 8036 8316 8585 8344
rect 1688 8248 1992 8276
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 8036 8276 8064 8316
rect 8573 8313 8585 8316
rect 8619 8313 8631 8347
rect 8573 8307 8631 8313
rect 11241 8347 11299 8353
rect 11241 8313 11253 8347
rect 11287 8344 11299 8347
rect 11698 8344 11704 8356
rect 11287 8316 11704 8344
rect 11287 8313 11299 8316
rect 11241 8307 11299 8313
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 11808 8353 11836 8384
rect 11793 8347 11851 8353
rect 11793 8313 11805 8347
rect 11839 8313 11851 8347
rect 11793 8307 11851 8313
rect 7064 8248 8064 8276
rect 7064 8236 7070 8248
rect 8110 8236 8116 8288
rect 8168 8236 8174 8288
rect 8754 8236 8760 8288
rect 8812 8236 8818 8288
rect 12360 8285 12388 8452
rect 12713 8449 12725 8452
rect 12759 8449 12771 8483
rect 12713 8443 12771 8449
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 16112 8483 16170 8489
rect 16112 8449 16124 8483
rect 16158 8449 16170 8483
rect 16112 8443 16170 8449
rect 16485 8483 16543 8489
rect 16485 8449 16497 8483
rect 16531 8480 16543 8483
rect 16574 8480 16580 8492
rect 16531 8452 16580 8480
rect 16531 8449 16543 8452
rect 16485 8443 16543 8449
rect 12802 8412 12808 8424
rect 12544 8384 12808 8412
rect 12544 8353 12572 8384
rect 12802 8372 12808 8384
rect 12860 8372 12866 8424
rect 16132 8412 16160 8443
rect 16574 8440 16580 8452
rect 16632 8440 16638 8492
rect 16684 8489 16712 8520
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 17402 8508 17408 8560
rect 17460 8508 17466 8560
rect 16669 8483 16727 8489
rect 16669 8449 16681 8483
rect 16715 8449 16727 8483
rect 16669 8443 16727 8449
rect 16684 8412 16712 8443
rect 16132 8384 16712 8412
rect 16942 8372 16948 8424
rect 17000 8372 17006 8424
rect 12529 8347 12587 8353
rect 12529 8313 12541 8347
rect 12575 8313 12587 8347
rect 12529 8307 12587 8313
rect 15930 8304 15936 8356
rect 15988 8304 15994 8356
rect 12345 8279 12403 8285
rect 12345 8245 12357 8279
rect 12391 8245 12403 8279
rect 12345 8239 12403 8245
rect 12805 8279 12863 8285
rect 12805 8245 12817 8279
rect 12851 8276 12863 8279
rect 13354 8276 13360 8288
rect 12851 8248 13360 8276
rect 12851 8245 12863 8248
rect 12805 8239 12863 8245
rect 13354 8236 13360 8248
rect 13412 8236 13418 8288
rect 1104 8186 22816 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 20214 8186
rect 20266 8134 20278 8186
rect 20330 8134 20342 8186
rect 20394 8134 20406 8186
rect 20458 8134 20470 8186
rect 20522 8134 22816 8186
rect 1104 8112 22816 8134
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 3513 8075 3571 8081
rect 3513 8072 3525 8075
rect 3108 8044 3525 8072
rect 3108 8032 3114 8044
rect 3436 7936 3464 8044
rect 3513 8041 3525 8044
rect 3559 8041 3571 8075
rect 3513 8035 3571 8041
rect 3602 8032 3608 8084
rect 3660 8072 3666 8084
rect 6181 8075 6239 8081
rect 6181 8072 6193 8075
rect 3660 8044 6193 8072
rect 3660 8032 3666 8044
rect 6181 8041 6193 8044
rect 6227 8041 6239 8075
rect 6181 8035 6239 8041
rect 8205 8075 8263 8081
rect 8205 8041 8217 8075
rect 8251 8072 8263 8075
rect 8294 8072 8300 8084
rect 8251 8044 8300 8072
rect 8251 8041 8263 8044
rect 8205 8035 8263 8041
rect 8294 8032 8300 8044
rect 8352 8032 8358 8084
rect 11146 8032 11152 8084
rect 11204 8072 11210 8084
rect 11609 8075 11667 8081
rect 11609 8072 11621 8075
rect 11204 8044 11621 8072
rect 11204 8032 11210 8044
rect 11609 8041 11621 8044
rect 11655 8041 11667 8075
rect 11609 8035 11667 8041
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 16301 8075 16359 8081
rect 12952 8044 13492 8072
rect 12952 8032 12958 8044
rect 4065 8007 4123 8013
rect 4065 7973 4077 8007
rect 4111 7973 4123 8007
rect 4065 7967 4123 7973
rect 3789 7939 3847 7945
rect 3789 7936 3801 7939
rect 3436 7908 3801 7936
rect 3789 7905 3801 7908
rect 3835 7905 3847 7939
rect 3789 7899 3847 7905
rect 1486 7828 1492 7880
rect 1544 7828 1550 7880
rect 1581 7871 1639 7877
rect 1581 7837 1593 7871
rect 1627 7868 1639 7871
rect 1765 7871 1823 7877
rect 1765 7868 1777 7871
rect 1627 7840 1777 7868
rect 1627 7837 1639 7840
rect 1581 7831 1639 7837
rect 1765 7837 1777 7840
rect 1811 7837 1823 7871
rect 3418 7868 3424 7880
rect 3174 7840 3424 7868
rect 1765 7831 1823 7837
rect 3418 7828 3424 7840
rect 3476 7828 3482 7880
rect 2038 7760 2044 7812
rect 2096 7760 2102 7812
rect 4080 7800 4108 7967
rect 6733 7939 6791 7945
rect 6733 7905 6745 7939
rect 6779 7936 6791 7939
rect 8110 7936 8116 7948
rect 6779 7908 8116 7936
rect 6779 7905 6791 7908
rect 6733 7899 6791 7905
rect 8110 7896 8116 7908
rect 8168 7896 8174 7948
rect 10778 7936 10784 7948
rect 10060 7908 10784 7936
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4433 7871 4491 7877
rect 4433 7868 4445 7871
rect 4212 7840 4445 7868
rect 4212 7828 4218 7840
rect 4433 7837 4445 7840
rect 4479 7837 4491 7871
rect 4433 7831 4491 7837
rect 5810 7828 5816 7880
rect 5868 7868 5874 7880
rect 5868 7840 6000 7868
rect 5868 7828 5874 7840
rect 3436 7772 4108 7800
rect 1578 7692 1584 7744
rect 1636 7732 1642 7744
rect 3436 7732 3464 7772
rect 4706 7760 4712 7812
rect 4764 7760 4770 7812
rect 5972 7800 6000 7840
rect 6454 7828 6460 7880
rect 6512 7828 6518 7880
rect 10060 7854 10088 7908
rect 10778 7896 10784 7908
rect 10836 7936 10842 7948
rect 10836 7908 11560 7936
rect 10836 7896 10842 7908
rect 11422 7828 11428 7880
rect 11480 7828 11486 7880
rect 11532 7868 11560 7908
rect 11698 7896 11704 7948
rect 11756 7936 11762 7948
rect 13081 7939 13139 7945
rect 13081 7936 13093 7939
rect 11756 7908 13093 7936
rect 11756 7896 11762 7908
rect 13081 7905 13093 7908
rect 13127 7905 13139 7939
rect 13081 7899 13139 7905
rect 13354 7896 13360 7948
rect 13412 7896 13418 7948
rect 13464 7877 13492 8044
rect 16301 8041 16313 8075
rect 16347 8072 16359 8075
rect 16482 8072 16488 8084
rect 16347 8044 16488 8072
rect 16347 8041 16359 8044
rect 16301 8035 16359 8041
rect 16482 8032 16488 8044
rect 16540 8032 16546 8084
rect 14553 7939 14611 7945
rect 14553 7905 14565 7939
rect 14599 7936 14611 7939
rect 14918 7936 14924 7948
rect 14599 7908 14924 7936
rect 14599 7905 14611 7908
rect 14553 7899 14611 7905
rect 14918 7896 14924 7908
rect 14976 7896 14982 7948
rect 13449 7871 13507 7877
rect 11532 7840 12006 7868
rect 13449 7837 13461 7871
rect 13495 7837 13507 7871
rect 13449 7831 13507 7837
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 11149 7803 11207 7809
rect 5972 7772 7222 7800
rect 11149 7769 11161 7803
rect 11195 7769 11207 7803
rect 13740 7800 13768 7831
rect 14274 7828 14280 7880
rect 14332 7828 14338 7880
rect 14829 7803 14887 7809
rect 13740 7772 14780 7800
rect 11149 7763 11207 7769
rect 1636 7704 3464 7732
rect 1636 7692 1642 7704
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4249 7735 4307 7741
rect 4249 7732 4261 7735
rect 3936 7704 4261 7732
rect 3936 7692 3942 7704
rect 4249 7701 4261 7704
rect 4295 7701 4307 7735
rect 4249 7695 4307 7701
rect 8018 7692 8024 7744
rect 8076 7732 8082 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 8076 7704 9689 7732
rect 8076 7692 8082 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 9677 7695 9735 7701
rect 10134 7692 10140 7744
rect 10192 7732 10198 7744
rect 11164 7732 11192 7763
rect 10192 7704 11192 7732
rect 10192 7692 10198 7704
rect 13722 7692 13728 7744
rect 13780 7692 13786 7744
rect 14090 7692 14096 7744
rect 14148 7732 14154 7744
rect 14185 7735 14243 7741
rect 14185 7732 14197 7735
rect 14148 7704 14197 7732
rect 14148 7692 14154 7704
rect 14185 7701 14197 7704
rect 14231 7701 14243 7735
rect 14752 7732 14780 7772
rect 14829 7769 14841 7803
rect 14875 7800 14887 7803
rect 15102 7800 15108 7812
rect 14875 7772 15108 7800
rect 14875 7769 14887 7772
rect 14829 7763 14887 7769
rect 15102 7760 15108 7772
rect 15160 7760 15166 7812
rect 15286 7760 15292 7812
rect 15344 7760 15350 7812
rect 15654 7732 15660 7744
rect 14752 7704 15660 7732
rect 14185 7695 14243 7701
rect 15654 7692 15660 7704
rect 15712 7692 15718 7744
rect 1104 7642 22816 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 22816 7642
rect 1104 7568 22816 7590
rect 2038 7488 2044 7540
rect 2096 7528 2102 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 2096 7500 3157 7528
rect 2096 7488 2102 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 3421 7531 3479 7537
rect 3421 7497 3433 7531
rect 3467 7528 3479 7531
rect 4154 7528 4160 7540
rect 3467 7500 4160 7528
rect 3467 7497 3479 7500
rect 3421 7491 3479 7497
rect 4154 7488 4160 7500
rect 4212 7488 4218 7540
rect 4706 7488 4712 7540
rect 4764 7528 4770 7540
rect 5353 7531 5411 7537
rect 5353 7528 5365 7531
rect 4764 7500 5365 7528
rect 4764 7488 4770 7500
rect 5353 7497 5365 7500
rect 5399 7497 5411 7531
rect 5353 7491 5411 7497
rect 6454 7488 6460 7540
rect 6512 7528 6518 7540
rect 6549 7531 6607 7537
rect 6549 7528 6561 7531
rect 6512 7500 6561 7528
rect 6512 7488 6518 7500
rect 6549 7497 6561 7500
rect 6595 7497 6607 7531
rect 6549 7491 6607 7497
rect 6730 7488 6736 7540
rect 6788 7528 6794 7540
rect 6825 7531 6883 7537
rect 6825 7528 6837 7531
rect 6788 7500 6837 7528
rect 6788 7488 6794 7500
rect 6825 7497 6837 7500
rect 6871 7497 6883 7531
rect 6825 7491 6883 7497
rect 9953 7531 10011 7537
rect 9953 7497 9965 7531
rect 9999 7528 10011 7531
rect 10134 7528 10140 7540
rect 9999 7500 10140 7528
rect 9999 7497 10011 7500
rect 9953 7491 10011 7497
rect 10134 7488 10140 7500
rect 10192 7488 10198 7540
rect 10689 7531 10747 7537
rect 10689 7497 10701 7531
rect 10735 7528 10747 7531
rect 11422 7528 11428 7540
rect 10735 7500 11428 7528
rect 10735 7497 10747 7500
rect 10689 7491 10747 7497
rect 11422 7488 11428 7500
rect 11480 7488 11486 7540
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 13504 7500 15608 7528
rect 13504 7488 13510 7500
rect 3878 7420 3884 7472
rect 3936 7420 3942 7472
rect 6362 7420 6368 7472
rect 6420 7460 6426 7472
rect 7745 7463 7803 7469
rect 6420 7432 7144 7460
rect 6420 7420 6426 7432
rect 1394 7352 1400 7404
rect 1452 7352 1458 7404
rect 1670 7284 1676 7336
rect 1728 7284 1734 7336
rect 2792 7324 2820 7378
rect 3234 7352 3240 7404
rect 3292 7392 3298 7404
rect 3329 7395 3387 7401
rect 3329 7392 3341 7395
rect 3292 7364 3341 7392
rect 3292 7352 3298 7364
rect 3329 7361 3341 7364
rect 3375 7392 3387 7395
rect 3605 7395 3663 7401
rect 3605 7392 3617 7395
rect 3375 7364 3617 7392
rect 3375 7361 3387 7364
rect 3329 7355 3387 7361
rect 3605 7361 3617 7364
rect 3651 7361 3663 7395
rect 5718 7392 5724 7404
rect 5014 7378 5724 7392
rect 3605 7355 3663 7361
rect 5000 7364 5724 7378
rect 3142 7324 3148 7336
rect 2792 7296 3148 7324
rect 3142 7284 3148 7296
rect 3200 7324 3206 7336
rect 5000 7324 5028 7364
rect 5718 7352 5724 7364
rect 5776 7352 5782 7404
rect 6656 7401 6684 7432
rect 6641 7395 6699 7401
rect 6641 7361 6653 7395
rect 6687 7361 6699 7395
rect 6641 7355 6699 7361
rect 6917 7395 6975 7401
rect 6917 7361 6929 7395
rect 6963 7361 6975 7395
rect 6917 7355 6975 7361
rect 3200 7296 5028 7324
rect 6932 7324 6960 7355
rect 7006 7352 7012 7404
rect 7064 7352 7070 7404
rect 7116 7392 7144 7432
rect 7745 7429 7757 7463
rect 7791 7460 7803 7463
rect 8110 7460 8116 7472
rect 7791 7432 8116 7460
rect 7791 7429 7803 7432
rect 7745 7423 7803 7429
rect 8110 7420 8116 7432
rect 8168 7420 8174 7472
rect 8481 7463 8539 7469
rect 8481 7429 8493 7463
rect 8527 7460 8539 7463
rect 8754 7460 8760 7472
rect 8527 7432 8760 7460
rect 8527 7429 8539 7432
rect 8481 7423 8539 7429
rect 8754 7420 8760 7432
rect 8812 7420 8818 7472
rect 9214 7420 9220 7472
rect 9272 7420 9278 7472
rect 10042 7420 10048 7472
rect 10100 7460 10106 7472
rect 10100 7432 10364 7460
rect 10100 7420 10106 7432
rect 7650 7401 7656 7404
rect 7648 7392 7656 7401
rect 7116 7364 7656 7392
rect 7648 7355 7656 7364
rect 7650 7352 7656 7355
rect 7708 7352 7714 7404
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7361 7895 7395
rect 7837 7355 7895 7361
rect 7852 7324 7880 7355
rect 8018 7352 8024 7404
rect 8076 7352 8082 7404
rect 10134 7352 10140 7404
rect 10192 7352 10198 7404
rect 10336 7401 10364 7432
rect 13722 7420 13728 7472
rect 13780 7420 13786 7472
rect 15580 7469 15608 7500
rect 15565 7463 15623 7469
rect 15565 7429 15577 7463
rect 15611 7460 15623 7463
rect 15611 7432 16160 7460
rect 15611 7429 15623 7432
rect 15565 7423 15623 7429
rect 10321 7395 10379 7401
rect 10321 7361 10333 7395
rect 10367 7361 10379 7395
rect 10321 7355 10379 7361
rect 10597 7395 10655 7401
rect 10597 7361 10609 7395
rect 10643 7361 10655 7395
rect 10597 7355 10655 7361
rect 8205 7327 8263 7333
rect 8205 7324 8217 7327
rect 6932 7296 7052 7324
rect 7852 7296 8217 7324
rect 3200 7284 3206 7296
rect 7024 7256 7052 7296
rect 8205 7293 8217 7296
rect 8251 7293 8263 7327
rect 8205 7287 8263 7293
rect 8018 7256 8024 7268
rect 7024 7228 8024 7256
rect 8018 7216 8024 7228
rect 8076 7216 8082 7268
rect 7466 7148 7472 7200
rect 7524 7148 7530 7200
rect 8220 7188 8248 7287
rect 9490 7284 9496 7336
rect 9548 7324 9554 7336
rect 10612 7324 10640 7355
rect 11054 7352 11060 7404
rect 11112 7352 11118 7404
rect 14826 7352 14832 7404
rect 14884 7392 14890 7404
rect 15286 7392 15292 7404
rect 14884 7364 15292 7392
rect 14884 7352 14890 7364
rect 15286 7352 15292 7364
rect 15344 7352 15350 7404
rect 15378 7352 15384 7404
rect 15436 7352 15442 7404
rect 15654 7352 15660 7404
rect 15712 7352 15718 7404
rect 16132 7401 16160 7432
rect 15795 7395 15853 7401
rect 15795 7361 15807 7395
rect 15841 7392 15853 7395
rect 16117 7395 16175 7401
rect 15841 7364 16068 7392
rect 15841 7361 15853 7364
rect 15795 7355 15853 7361
rect 9548 7296 10640 7324
rect 9548 7284 9554 7296
rect 12894 7284 12900 7336
rect 12952 7324 12958 7336
rect 13357 7327 13415 7333
rect 12952 7296 13032 7324
rect 12952 7284 12958 7296
rect 10413 7259 10471 7265
rect 10413 7225 10425 7259
rect 10459 7256 10471 7259
rect 10686 7256 10692 7268
rect 10459 7228 10692 7256
rect 10459 7225 10471 7228
rect 10413 7219 10471 7225
rect 10686 7216 10692 7228
rect 10744 7216 10750 7268
rect 13004 7265 13032 7296
rect 13357 7293 13369 7327
rect 13403 7293 13415 7327
rect 13357 7287 13415 7293
rect 12989 7259 13047 7265
rect 12989 7225 13001 7259
rect 13035 7225 13047 7259
rect 12989 7219 13047 7225
rect 9490 7188 9496 7200
rect 8220 7160 9496 7188
rect 9490 7148 9496 7160
rect 9548 7148 9554 7200
rect 11146 7148 11152 7200
rect 11204 7148 11210 7200
rect 12894 7148 12900 7200
rect 12952 7148 12958 7200
rect 13372 7188 13400 7287
rect 13446 7284 13452 7336
rect 13504 7284 13510 7336
rect 13814 7284 13820 7336
rect 13872 7324 13878 7336
rect 14274 7324 14280 7336
rect 13872 7296 14280 7324
rect 13872 7284 13878 7296
rect 14274 7284 14280 7296
rect 14332 7324 14338 7336
rect 16040 7324 16068 7364
rect 16117 7361 16129 7395
rect 16163 7361 16175 7395
rect 16117 7355 16175 7361
rect 22094 7324 22100 7336
rect 14332 7296 22100 7324
rect 14332 7284 14338 7296
rect 22094 7284 22100 7296
rect 22152 7284 22158 7336
rect 15378 7256 15384 7268
rect 14752 7228 15384 7256
rect 14752 7188 14780 7228
rect 15378 7216 15384 7228
rect 15436 7216 15442 7268
rect 15933 7259 15991 7265
rect 15933 7225 15945 7259
rect 15979 7256 15991 7259
rect 19978 7256 19984 7268
rect 15979 7228 19984 7256
rect 15979 7225 15991 7228
rect 15933 7219 15991 7225
rect 19978 7216 19984 7228
rect 20036 7216 20042 7268
rect 13372 7160 14780 7188
rect 15197 7191 15255 7197
rect 15197 7157 15209 7191
rect 15243 7188 15255 7191
rect 15838 7188 15844 7200
rect 15243 7160 15844 7188
rect 15243 7157 15255 7160
rect 15197 7151 15255 7157
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 16022 7148 16028 7200
rect 16080 7188 16086 7200
rect 16209 7191 16267 7197
rect 16209 7188 16221 7191
rect 16080 7160 16221 7188
rect 16080 7148 16086 7160
rect 16209 7157 16221 7160
rect 16255 7157 16267 7191
rect 16209 7151 16267 7157
rect 1104 7098 22816 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 20214 7098
rect 20266 7046 20278 7098
rect 20330 7046 20342 7098
rect 20394 7046 20406 7098
rect 20458 7046 20470 7098
rect 20522 7046 22816 7098
rect 1104 7024 22816 7046
rect 2028 6987 2086 6993
rect 2028 6953 2040 6987
rect 2074 6984 2086 6987
rect 7466 6984 7472 6996
rect 2074 6956 7472 6984
rect 2074 6953 2086 6956
rect 2028 6947 2086 6953
rect 7466 6944 7472 6956
rect 7524 6944 7530 6996
rect 9398 6984 9404 6996
rect 8036 6956 9404 6984
rect 3234 6876 3240 6928
rect 3292 6916 3298 6928
rect 3513 6919 3571 6925
rect 3513 6916 3525 6919
rect 3292 6888 3525 6916
rect 3292 6876 3298 6888
rect 3513 6885 3525 6888
rect 3559 6885 3571 6919
rect 7101 6919 7159 6925
rect 3513 6879 3571 6885
rect 4816 6888 5488 6916
rect 1762 6808 1768 6860
rect 1820 6808 1826 6860
rect 3878 6808 3884 6860
rect 3936 6848 3942 6860
rect 4816 6848 4844 6888
rect 5353 6851 5411 6857
rect 5353 6848 5365 6851
rect 3936 6820 4568 6848
rect 3936 6808 3942 6820
rect 3142 6740 3148 6792
rect 3200 6740 3206 6792
rect 3326 6740 3332 6792
rect 3384 6780 3390 6792
rect 4540 6789 4568 6820
rect 4632 6820 4844 6848
rect 5000 6820 5365 6848
rect 4157 6783 4215 6789
rect 4157 6780 4169 6783
rect 3384 6752 4169 6780
rect 3384 6740 3390 6752
rect 4157 6749 4169 6752
rect 4203 6749 4215 6783
rect 4530 6783 4588 6789
rect 4157 6743 4215 6749
rect 4264 6752 4476 6780
rect 3970 6672 3976 6724
rect 4028 6712 4034 6724
rect 4264 6712 4292 6752
rect 4028 6684 4292 6712
rect 4028 6672 4034 6684
rect 4338 6672 4344 6724
rect 4396 6672 4402 6724
rect 4448 6721 4476 6752
rect 4530 6749 4542 6783
rect 4576 6749 4588 6783
rect 4530 6743 4588 6749
rect 4433 6715 4491 6721
rect 4433 6681 4445 6715
rect 4479 6712 4491 6715
rect 4632 6712 4660 6820
rect 4726 6783 4784 6789
rect 4726 6749 4738 6783
rect 4772 6780 4784 6783
rect 5000 6780 5028 6820
rect 5353 6817 5365 6820
rect 5399 6817 5411 6851
rect 5460 6848 5488 6888
rect 7101 6885 7113 6919
rect 7147 6916 7159 6919
rect 7190 6916 7196 6928
rect 7147 6888 7196 6916
rect 7147 6885 7159 6888
rect 7101 6879 7159 6885
rect 7190 6876 7196 6888
rect 7248 6916 7254 6928
rect 8036 6916 8064 6956
rect 9398 6944 9404 6956
rect 9456 6944 9462 6996
rect 9490 6944 9496 6996
rect 9548 6944 9554 6996
rect 10400 6987 10458 6993
rect 10400 6953 10412 6987
rect 10446 6984 10458 6987
rect 11422 6984 11428 6996
rect 10446 6956 11428 6984
rect 10446 6953 10458 6956
rect 10400 6947 10458 6953
rect 11422 6944 11428 6956
rect 11480 6944 11486 6996
rect 12332 6987 12390 6993
rect 12332 6953 12344 6987
rect 12378 6984 12390 6987
rect 12894 6984 12900 6996
rect 12378 6956 12900 6984
rect 12378 6953 12390 6956
rect 12332 6947 12390 6953
rect 12894 6944 12900 6956
rect 12952 6944 12958 6996
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 16282 6987 16340 6993
rect 16282 6984 16294 6987
rect 15896 6956 16294 6984
rect 15896 6944 15902 6956
rect 16282 6953 16294 6956
rect 16328 6953 16340 6987
rect 16282 6947 16340 6953
rect 7248 6888 8064 6916
rect 9048 6888 10272 6916
rect 7248 6876 7254 6888
rect 9048 6848 9076 6888
rect 10137 6851 10195 6857
rect 10137 6848 10149 6851
rect 5460 6820 9076 6848
rect 9232 6820 10149 6848
rect 5353 6811 5411 6817
rect 4772 6752 5028 6780
rect 5077 6783 5135 6789
rect 4772 6749 4784 6752
rect 4726 6743 4784 6749
rect 5077 6749 5089 6783
rect 5123 6749 5135 6783
rect 5077 6743 5135 6749
rect 4479 6684 4660 6712
rect 5092 6712 5120 6743
rect 6914 6740 6920 6792
rect 6972 6780 6978 6792
rect 9232 6789 9260 6820
rect 10137 6817 10149 6820
rect 10183 6817 10195 6851
rect 10244 6848 10272 6888
rect 15378 6876 15384 6928
rect 15436 6916 15442 6928
rect 15436 6888 16160 6916
rect 15436 6876 15442 6888
rect 12069 6851 12127 6857
rect 12069 6848 12081 6851
rect 10244 6820 12081 6848
rect 10137 6811 10195 6817
rect 12069 6817 12081 6820
rect 12115 6848 12127 6851
rect 13814 6848 13820 6860
rect 12115 6820 13820 6848
rect 12115 6817 12127 6820
rect 12069 6811 12127 6817
rect 13814 6808 13820 6820
rect 13872 6808 13878 6860
rect 14090 6808 14096 6860
rect 14148 6808 14154 6860
rect 15654 6808 15660 6860
rect 15712 6848 15718 6860
rect 15841 6851 15899 6857
rect 15841 6848 15853 6851
rect 15712 6820 15853 6848
rect 15712 6808 15718 6820
rect 15841 6817 15853 6820
rect 15887 6817 15899 6851
rect 15841 6811 15899 6817
rect 16022 6808 16028 6860
rect 16080 6808 16086 6860
rect 16132 6848 16160 6888
rect 17773 6851 17831 6857
rect 17773 6848 17785 6851
rect 16132 6820 17785 6848
rect 17773 6817 17785 6820
rect 17819 6817 17831 6851
rect 17773 6811 17831 6817
rect 7653 6783 7711 6789
rect 7653 6780 7665 6783
rect 6972 6752 7665 6780
rect 6972 6740 6978 6752
rect 7653 6749 7665 6752
rect 7699 6749 7711 6783
rect 7653 6743 7711 6749
rect 8113 6783 8171 6789
rect 8113 6749 8125 6783
rect 8159 6780 8171 6783
rect 9217 6783 9275 6789
rect 9217 6780 9229 6783
rect 8159 6752 9229 6780
rect 8159 6749 8171 6752
rect 8113 6743 8171 6749
rect 9217 6749 9229 6752
rect 9263 6749 9275 6783
rect 9217 6743 9275 6749
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9364 6752 9449 6780
rect 9364 6740 9370 6752
rect 5534 6712 5540 6724
rect 5092 6684 5540 6712
rect 4479 6681 4491 6684
rect 4433 6675 4491 6681
rect 5534 6672 5540 6684
rect 5592 6672 5598 6724
rect 5626 6672 5632 6724
rect 5684 6672 5690 6724
rect 5718 6672 5724 6724
rect 5776 6712 5782 6724
rect 5776 6684 6118 6712
rect 5776 6672 5782 6684
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4985 6647 5043 6653
rect 4985 6644 4997 6647
rect 4120 6616 4997 6644
rect 4120 6604 4126 6616
rect 4985 6613 4997 6616
rect 5031 6613 5043 6647
rect 4985 6607 5043 6613
rect 7285 6647 7343 6653
rect 7285 6613 7297 6647
rect 7331 6644 7343 6647
rect 7742 6644 7748 6656
rect 7331 6616 7748 6644
rect 7331 6613 7343 6616
rect 7285 6607 7343 6613
rect 7742 6604 7748 6616
rect 7800 6604 7806 6656
rect 9421 6644 9449 6752
rect 9490 6740 9496 6792
rect 9548 6780 9554 6792
rect 9672 6783 9730 6789
rect 9672 6780 9684 6783
rect 9548 6752 9684 6780
rect 9548 6740 9554 6752
rect 9672 6749 9684 6752
rect 9718 6780 9730 6783
rect 9718 6752 9996 6780
rect 9718 6749 9730 6752
rect 9672 6743 9730 6749
rect 9766 6672 9772 6724
rect 9824 6672 9830 6724
rect 9861 6715 9919 6721
rect 9861 6681 9873 6715
rect 9907 6681 9919 6715
rect 9861 6675 9919 6681
rect 9876 6644 9904 6675
rect 9421 6616 9904 6644
rect 9968 6644 9996 6752
rect 10042 6740 10048 6792
rect 10100 6740 10106 6792
rect 11790 6712 11796 6724
rect 11638 6684 11796 6712
rect 11790 6672 11796 6684
rect 11848 6672 11854 6724
rect 13354 6672 13360 6724
rect 13412 6672 13418 6724
rect 14369 6715 14427 6721
rect 14369 6681 14381 6715
rect 14415 6681 14427 6715
rect 14369 6675 14427 6681
rect 11054 6644 11060 6656
rect 9968 6616 11060 6644
rect 11054 6604 11060 6616
rect 11112 6604 11118 6656
rect 11238 6604 11244 6656
rect 11296 6644 11302 6656
rect 11885 6647 11943 6653
rect 11885 6644 11897 6647
rect 11296 6616 11897 6644
rect 11296 6604 11302 6616
rect 11885 6613 11897 6616
rect 11931 6613 11943 6647
rect 11885 6607 11943 6613
rect 13817 6647 13875 6653
rect 13817 6613 13829 6647
rect 13863 6644 13875 6647
rect 14384 6644 14412 6675
rect 14918 6672 14924 6724
rect 14976 6672 14982 6724
rect 15672 6684 16790 6712
rect 13863 6616 14412 6644
rect 13863 6613 13875 6616
rect 13817 6607 13875 6613
rect 15102 6604 15108 6656
rect 15160 6644 15166 6656
rect 15672 6644 15700 6684
rect 15160 6616 15700 6644
rect 15160 6604 15166 6616
rect 1104 6554 22816 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 22816 6554
rect 1104 6480 22816 6502
rect 1670 6400 1676 6452
rect 1728 6400 1734 6452
rect 3142 6400 3148 6452
rect 3200 6440 3206 6452
rect 3970 6440 3976 6452
rect 3200 6412 3976 6440
rect 3200 6400 3206 6412
rect 3970 6400 3976 6412
rect 4028 6400 4034 6452
rect 5534 6400 5540 6452
rect 5592 6440 5598 6452
rect 6730 6440 6736 6452
rect 5592 6412 6736 6440
rect 5592 6400 5598 6412
rect 6730 6400 6736 6412
rect 6788 6400 6794 6452
rect 6825 6443 6883 6449
rect 6825 6409 6837 6443
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 9217 6443 9275 6449
rect 9217 6409 9229 6443
rect 9263 6440 9275 6443
rect 9306 6440 9312 6452
rect 9263 6412 9312 6440
rect 9263 6409 9275 6412
rect 9217 6403 9275 6409
rect 3602 6372 3608 6384
rect 1780 6344 3608 6372
rect 1578 6264 1584 6316
rect 1636 6264 1642 6316
rect 1780 6313 1808 6344
rect 3602 6332 3608 6344
rect 3660 6332 3666 6384
rect 3786 6332 3792 6384
rect 3844 6332 3850 6384
rect 4062 6332 4068 6384
rect 4120 6332 4126 6384
rect 5626 6332 5632 6384
rect 5684 6372 5690 6384
rect 5813 6375 5871 6381
rect 5813 6372 5825 6375
rect 5684 6344 5825 6372
rect 5684 6332 5690 6344
rect 5813 6341 5825 6344
rect 5859 6341 5871 6375
rect 6840 6372 6868 6403
rect 9306 6400 9312 6412
rect 9364 6400 9370 6452
rect 10042 6400 10048 6452
rect 10100 6440 10106 6452
rect 11149 6443 11207 6449
rect 10100 6412 11008 6440
rect 10100 6400 10106 6412
rect 5813 6335 5871 6341
rect 6012 6344 6868 6372
rect 1765 6307 1823 6313
rect 1765 6273 1777 6307
rect 1811 6273 1823 6307
rect 1765 6267 1823 6273
rect 1946 6264 1952 6316
rect 2004 6304 2010 6316
rect 2130 6313 2136 6316
rect 2128 6304 2136 6313
rect 2004 6276 2136 6304
rect 2004 6264 2010 6276
rect 2128 6267 2136 6276
rect 2130 6264 2136 6267
rect 2188 6264 2194 6316
rect 2222 6264 2228 6316
rect 2280 6264 2286 6316
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2501 6307 2559 6313
rect 2501 6273 2513 6307
rect 2547 6273 2559 6307
rect 2501 6267 2559 6273
rect 1026 6196 1032 6248
rect 1084 6236 1090 6248
rect 2516 6236 2544 6267
rect 2774 6264 2780 6316
rect 2832 6264 2838 6316
rect 2869 6307 2927 6313
rect 2869 6273 2881 6307
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 2884 6236 2912 6267
rect 3050 6264 3056 6316
rect 3108 6264 3114 6316
rect 3142 6264 3148 6316
rect 3200 6264 3206 6316
rect 3289 6307 3347 6313
rect 3289 6273 3301 6307
rect 3335 6304 3347 6307
rect 3804 6304 3832 6332
rect 5718 6304 5724 6316
rect 3335 6276 3832 6304
rect 5198 6276 5724 6304
rect 3335 6273 3347 6276
rect 3289 6267 3347 6273
rect 5718 6264 5724 6276
rect 5776 6264 5782 6316
rect 6012 6313 6040 6344
rect 7742 6332 7748 6384
rect 7800 6332 7806 6384
rect 5997 6307 6055 6313
rect 5997 6273 6009 6307
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6181 6307 6239 6313
rect 6181 6273 6193 6307
rect 6227 6304 6239 6307
rect 6227 6276 6776 6304
rect 6227 6273 6239 6276
rect 6181 6267 6239 6273
rect 3789 6239 3847 6245
rect 1084 6208 3372 6236
rect 1084 6196 1090 6208
rect 3344 6180 3372 6208
rect 3789 6205 3801 6239
rect 3835 6205 3847 6239
rect 3789 6199 3847 6205
rect 1486 6128 1492 6180
rect 1544 6168 1550 6180
rect 1949 6171 2007 6177
rect 1949 6168 1961 6171
rect 1544 6140 1961 6168
rect 1544 6128 1550 6140
rect 1949 6137 1961 6140
rect 1995 6137 2007 6171
rect 1949 6131 2007 6137
rect 2222 6128 2228 6180
rect 2280 6168 2286 6180
rect 2774 6168 2780 6180
rect 2280 6140 2780 6168
rect 2280 6128 2286 6140
rect 2774 6128 2780 6140
rect 2832 6168 2838 6180
rect 3142 6168 3148 6180
rect 2832 6140 3148 6168
rect 2832 6128 2838 6140
rect 3142 6128 3148 6140
rect 3200 6128 3206 6180
rect 3326 6128 3332 6180
rect 3384 6128 3390 6180
rect 3421 6171 3479 6177
rect 3421 6137 3433 6171
rect 3467 6168 3479 6171
rect 3804 6168 3832 6199
rect 6546 6196 6552 6248
rect 6604 6236 6610 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6604 6208 6653 6236
rect 6604 6196 6610 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6748 6236 6776 6276
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 7190 6264 7196 6316
rect 7248 6264 7254 6316
rect 8754 6264 8760 6316
rect 8812 6304 8818 6316
rect 9324 6304 9352 6400
rect 10980 6372 11008 6412
rect 11149 6409 11161 6443
rect 11195 6440 11207 6443
rect 11422 6440 11428 6452
rect 11195 6412 11428 6440
rect 11195 6409 11207 6412
rect 11149 6403 11207 6409
rect 11422 6400 11428 6412
rect 11480 6400 11486 6452
rect 11238 6372 11244 6384
rect 10980 6344 11244 6372
rect 11238 6332 11244 6344
rect 11296 6332 11302 6384
rect 13354 6372 13360 6384
rect 13110 6344 13360 6372
rect 13354 6332 13360 6344
rect 13412 6372 13418 6384
rect 14918 6372 14924 6384
rect 13412 6344 14924 6372
rect 13412 6332 13418 6344
rect 14918 6332 14924 6344
rect 14976 6332 14982 6384
rect 9401 6307 9459 6313
rect 9401 6304 9413 6307
rect 8812 6276 8878 6304
rect 9324 6276 9413 6304
rect 8812 6264 8818 6276
rect 9401 6273 9413 6276
rect 9447 6273 9459 6307
rect 9401 6267 9459 6273
rect 10778 6264 10784 6316
rect 10836 6264 10842 6316
rect 11146 6264 11152 6316
rect 11204 6304 11210 6316
rect 11609 6307 11667 6313
rect 11609 6304 11621 6307
rect 11204 6276 11621 6304
rect 11204 6264 11210 6276
rect 11609 6273 11621 6276
rect 11655 6273 11667 6307
rect 11609 6267 11667 6273
rect 6914 6236 6920 6248
rect 6748 6208 6920 6236
rect 6641 6199 6699 6205
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7469 6239 7527 6245
rect 7469 6205 7481 6239
rect 7515 6205 7527 6239
rect 7469 6199 7527 6205
rect 9677 6239 9735 6245
rect 9677 6205 9689 6239
rect 9723 6236 9735 6239
rect 9766 6236 9772 6248
rect 9723 6208 9772 6236
rect 9723 6205 9735 6208
rect 9677 6199 9735 6205
rect 3467 6140 3832 6168
rect 3467 6137 3479 6140
rect 3421 6131 3479 6137
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 7484 6168 7512 6199
rect 9766 6196 9772 6208
rect 9824 6196 9830 6248
rect 11885 6239 11943 6245
rect 11885 6205 11897 6239
rect 11931 6236 11943 6239
rect 11974 6236 11980 6248
rect 11931 6208 11980 6236
rect 11931 6205 11943 6208
rect 11885 6199 11943 6205
rect 11974 6196 11980 6208
rect 12032 6196 12038 6248
rect 5500 6140 7512 6168
rect 5500 6128 5506 6140
rect 2682 6060 2688 6112
rect 2740 6060 2746 6112
rect 3050 6060 3056 6112
rect 3108 6100 3114 6112
rect 4246 6100 4252 6112
rect 3108 6072 4252 6100
rect 3108 6060 3114 6072
rect 4246 6060 4252 6072
rect 4304 6060 4310 6112
rect 7098 6060 7104 6112
rect 7156 6100 7162 6112
rect 9674 6100 9680 6112
rect 7156 6072 9680 6100
rect 7156 6060 7162 6072
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 10042 6060 10048 6112
rect 10100 6100 10106 6112
rect 13357 6103 13415 6109
rect 13357 6100 13369 6103
rect 10100 6072 13369 6100
rect 10100 6060 10106 6072
rect 13357 6069 13369 6072
rect 13403 6069 13415 6103
rect 13357 6063 13415 6069
rect 1104 6010 22816 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 20214 6010
rect 20266 5958 20278 6010
rect 20330 5958 20342 6010
rect 20394 5958 20406 6010
rect 20458 5958 20470 6010
rect 20522 5958 22816 6010
rect 1104 5936 22816 5958
rect 2130 5856 2136 5908
rect 2188 5896 2194 5908
rect 4525 5899 4583 5905
rect 2188 5868 3556 5896
rect 2188 5856 2194 5868
rect 1765 5763 1823 5769
rect 1765 5729 1777 5763
rect 1811 5760 1823 5763
rect 2682 5760 2688 5772
rect 1811 5732 2688 5760
rect 1811 5729 1823 5732
rect 1765 5723 1823 5729
rect 2682 5720 2688 5732
rect 2740 5720 2746 5772
rect 3528 5769 3556 5868
rect 4525 5865 4537 5899
rect 4571 5896 4583 5899
rect 5442 5896 5448 5908
rect 4571 5868 5448 5896
rect 4571 5865 4583 5868
rect 4525 5859 4583 5865
rect 5442 5856 5448 5868
rect 5500 5856 5506 5908
rect 6546 5856 6552 5908
rect 6604 5896 6610 5908
rect 6825 5899 6883 5905
rect 6825 5896 6837 5899
rect 6604 5868 6837 5896
rect 6604 5856 6610 5868
rect 6825 5865 6837 5868
rect 6871 5896 6883 5899
rect 6871 5868 7328 5896
rect 6871 5865 6883 5868
rect 6825 5859 6883 5865
rect 3602 5788 3608 5840
rect 3660 5828 3666 5840
rect 5718 5828 5724 5840
rect 3660 5800 5724 5828
rect 3660 5788 3666 5800
rect 5718 5788 5724 5800
rect 5776 5788 5782 5840
rect 6641 5831 6699 5837
rect 6641 5797 6653 5831
rect 6687 5828 6699 5831
rect 6914 5828 6920 5840
rect 6687 5800 6920 5828
rect 6687 5797 6699 5800
rect 6641 5791 6699 5797
rect 6914 5788 6920 5800
rect 6972 5788 6978 5840
rect 3513 5763 3571 5769
rect 3513 5729 3525 5763
rect 3559 5760 3571 5763
rect 3878 5760 3884 5772
rect 3559 5732 3884 5760
rect 3559 5729 3571 5732
rect 3513 5723 3571 5729
rect 3878 5720 3884 5732
rect 3936 5760 3942 5772
rect 3936 5732 4384 5760
rect 3936 5720 3942 5732
rect 3326 5652 3332 5704
rect 3384 5692 3390 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3384 5664 3985 5692
rect 3384 5652 3390 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4356 5701 4384 5732
rect 5534 5720 5540 5772
rect 5592 5720 5598 5772
rect 7300 5760 7328 5868
rect 7650 5856 7656 5908
rect 7708 5856 7714 5908
rect 9585 5899 9643 5905
rect 9585 5865 9597 5899
rect 9631 5896 9643 5899
rect 9766 5896 9772 5908
rect 9631 5868 9772 5896
rect 9631 5865 9643 5868
rect 9585 5859 9643 5865
rect 9766 5856 9772 5868
rect 9824 5856 9830 5908
rect 11974 5856 11980 5908
rect 12032 5896 12038 5908
rect 12161 5899 12219 5905
rect 12161 5896 12173 5899
rect 12032 5868 12173 5896
rect 12032 5856 12038 5868
rect 12161 5865 12173 5868
rect 12207 5865 12219 5899
rect 12161 5859 12219 5865
rect 13538 5856 13544 5908
rect 13596 5896 13602 5908
rect 14093 5899 14151 5905
rect 14093 5896 14105 5899
rect 13596 5868 14105 5896
rect 13596 5856 13602 5868
rect 14093 5865 14105 5868
rect 14139 5865 14151 5899
rect 14093 5859 14151 5865
rect 7374 5788 7380 5840
rect 7432 5828 7438 5840
rect 8481 5831 8539 5837
rect 8481 5828 8493 5831
rect 7432 5800 8493 5828
rect 7432 5788 7438 5800
rect 8481 5797 8493 5800
rect 8527 5828 8539 5831
rect 9677 5831 9735 5837
rect 9677 5828 9689 5831
rect 8527 5800 9689 5828
rect 8527 5797 8539 5800
rect 8481 5791 8539 5797
rect 9677 5797 9689 5800
rect 9723 5828 9735 5831
rect 10134 5828 10140 5840
rect 9723 5800 10140 5828
rect 9723 5797 9735 5800
rect 9677 5791 9735 5797
rect 10134 5788 10140 5800
rect 10192 5788 10198 5840
rect 7300 5732 8616 5760
rect 4249 5695 4307 5701
rect 4249 5692 4261 5695
rect 4120 5664 4261 5692
rect 4120 5652 4126 5664
rect 4249 5661 4261 5664
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4346 5695 4404 5701
rect 4346 5661 4358 5695
rect 4392 5661 4404 5695
rect 4346 5655 4404 5661
rect 2038 5584 2044 5636
rect 2096 5584 2102 5636
rect 3418 5624 3424 5636
rect 3266 5596 3424 5624
rect 3418 5584 3424 5596
rect 3476 5624 3482 5636
rect 3602 5624 3608 5636
rect 3476 5596 3608 5624
rect 3476 5584 3482 5596
rect 3602 5584 3608 5596
rect 3660 5584 3666 5636
rect 3786 5584 3792 5636
rect 3844 5624 3850 5636
rect 4157 5627 4215 5633
rect 4157 5624 4169 5627
rect 3844 5596 4169 5624
rect 3844 5584 3850 5596
rect 4157 5593 4169 5596
rect 4203 5593 4215 5627
rect 4157 5587 4215 5593
rect 4706 5584 4712 5636
rect 4764 5584 4770 5636
rect 5644 5624 5672 5678
rect 6178 5652 6184 5704
rect 6236 5652 6242 5704
rect 6457 5695 6515 5701
rect 6457 5661 6469 5695
rect 6503 5692 6515 5695
rect 7098 5692 7104 5704
rect 6503 5664 7104 5692
rect 6503 5661 6515 5664
rect 6457 5655 6515 5661
rect 7098 5652 7104 5664
rect 7156 5652 7162 5704
rect 7300 5701 7328 5732
rect 8588 5704 8616 5732
rect 10042 5720 10048 5772
rect 10100 5720 10106 5772
rect 10413 5763 10471 5769
rect 10413 5729 10425 5763
rect 10459 5760 10471 5763
rect 11054 5760 11060 5772
rect 10459 5732 11060 5760
rect 10459 5729 10471 5732
rect 10413 5723 10471 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 11330 5720 11336 5772
rect 11388 5760 11394 5772
rect 11698 5760 11704 5772
rect 11388 5732 11704 5760
rect 11388 5720 11394 5732
rect 11698 5720 11704 5732
rect 11756 5760 11762 5772
rect 11756 5732 12480 5760
rect 11756 5720 11762 5732
rect 7558 5701 7564 5704
rect 7285 5695 7343 5701
rect 7285 5661 7297 5695
rect 7331 5661 7343 5695
rect 7285 5655 7343 5661
rect 7521 5695 7564 5701
rect 7521 5661 7533 5695
rect 7521 5655 7564 5661
rect 7558 5652 7564 5655
rect 7616 5652 7622 5704
rect 7837 5695 7895 5701
rect 7837 5692 7849 5695
rect 7663 5664 7849 5692
rect 6546 5624 6552 5636
rect 5644 5596 6552 5624
rect 6546 5584 6552 5596
rect 6604 5584 6610 5636
rect 6730 5584 6736 5636
rect 6788 5624 6794 5636
rect 7009 5627 7067 5633
rect 7009 5624 7021 5627
rect 6788 5596 7021 5624
rect 6788 5584 6794 5596
rect 7009 5593 7021 5596
rect 7055 5624 7067 5627
rect 7377 5627 7435 5633
rect 7377 5624 7389 5627
rect 7055 5596 7389 5624
rect 7055 5593 7067 5596
rect 7009 5587 7067 5593
rect 7377 5593 7389 5596
rect 7423 5624 7435 5627
rect 7663 5624 7691 5664
rect 7837 5661 7849 5664
rect 7883 5661 7895 5695
rect 7837 5655 7895 5661
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 8941 5695 8999 5701
rect 8941 5692 8953 5695
rect 8628 5664 8953 5692
rect 8628 5652 8634 5664
rect 8941 5661 8953 5664
rect 8987 5661 8999 5695
rect 8941 5655 8999 5661
rect 11790 5652 11796 5704
rect 11848 5652 11854 5704
rect 12452 5701 12480 5732
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12526 5652 12532 5704
rect 12584 5692 12590 5704
rect 12621 5695 12679 5701
rect 12621 5692 12633 5695
rect 12584 5664 12633 5692
rect 12584 5652 12590 5664
rect 12621 5661 12633 5664
rect 12667 5661 12679 5695
rect 12621 5655 12679 5661
rect 12710 5652 12716 5704
rect 12768 5692 12774 5704
rect 12989 5695 13047 5701
rect 12989 5692 13001 5695
rect 12768 5664 13001 5692
rect 12768 5652 12774 5664
rect 12989 5661 13001 5664
rect 13035 5661 13047 5695
rect 12989 5655 13047 5661
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 14918 5692 14924 5704
rect 14783 5664 14924 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 14918 5652 14924 5664
rect 14976 5652 14982 5704
rect 7423 5596 7691 5624
rect 8205 5627 8263 5633
rect 7423 5593 7435 5596
rect 7377 5587 7435 5593
rect 8205 5593 8217 5627
rect 8251 5624 8263 5627
rect 8846 5624 8852 5636
rect 8251 5596 8852 5624
rect 8251 5593 8263 5596
rect 8205 5587 8263 5593
rect 8846 5584 8852 5596
rect 8904 5584 8910 5636
rect 10686 5584 10692 5636
rect 10744 5584 10750 5636
rect 2314 5516 2320 5568
rect 2372 5556 2378 5568
rect 3050 5556 3056 5568
rect 2372 5528 3056 5556
rect 2372 5516 2378 5528
rect 3050 5516 3056 5528
rect 3108 5556 3114 5568
rect 3804 5556 3832 5584
rect 3108 5528 3832 5556
rect 6181 5559 6239 5565
rect 3108 5516 3114 5528
rect 6181 5525 6193 5559
rect 6227 5556 6239 5559
rect 6270 5556 6276 5568
rect 6227 5528 6276 5556
rect 6227 5525 6239 5528
rect 6181 5519 6239 5525
rect 6270 5516 6276 5528
rect 6328 5516 6334 5568
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 6914 5556 6920 5568
rect 6871 5528 6920 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 6914 5516 6920 5528
rect 6972 5516 6978 5568
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 7156 5528 7941 5556
rect 7156 5516 7162 5528
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 7929 5519 7987 5525
rect 8662 5516 8668 5568
rect 8720 5516 8726 5568
rect 9030 5516 9036 5568
rect 9088 5516 9094 5568
rect 9306 5516 9312 5568
rect 9364 5556 9370 5568
rect 11808 5556 11836 5652
rect 9364 5528 11836 5556
rect 12621 5559 12679 5565
rect 9364 5516 9370 5528
rect 12621 5525 12633 5559
rect 12667 5556 12679 5559
rect 12710 5556 12716 5568
rect 12667 5528 12716 5556
rect 12667 5525 12679 5528
rect 12621 5519 12679 5525
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13078 5516 13084 5568
rect 13136 5516 13142 5568
rect 1104 5466 22816 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 22816 5466
rect 1104 5392 22816 5414
rect 1489 5355 1547 5361
rect 1489 5321 1501 5355
rect 1535 5352 1547 5355
rect 2038 5352 2044 5364
rect 1535 5324 2044 5352
rect 1535 5321 1547 5324
rect 1489 5315 1547 5321
rect 2038 5312 2044 5324
rect 2096 5312 2102 5364
rect 3418 5352 3424 5364
rect 3160 5324 3424 5352
rect 3160 5284 3188 5324
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 6089 5355 6147 5361
rect 6089 5321 6101 5355
rect 6135 5352 6147 5355
rect 6546 5352 6552 5364
rect 6135 5324 6552 5352
rect 6135 5321 6147 5324
rect 6089 5315 6147 5321
rect 6546 5312 6552 5324
rect 6604 5312 6610 5364
rect 7558 5312 7564 5364
rect 7616 5352 7622 5364
rect 8846 5352 8852 5364
rect 7616 5324 8852 5352
rect 7616 5312 7622 5324
rect 8846 5312 8852 5324
rect 8904 5312 8910 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 10965 5355 11023 5361
rect 10965 5352 10977 5355
rect 9732 5324 10977 5352
rect 9732 5312 9738 5324
rect 10965 5321 10977 5324
rect 11011 5321 11023 5355
rect 15105 5355 15163 5361
rect 15105 5352 15117 5355
rect 10965 5315 11023 5321
rect 12084 5324 15117 5352
rect 3881 5287 3939 5293
rect 3881 5284 3893 5287
rect 2530 5256 3188 5284
rect 3252 5256 3893 5284
rect 3252 5225 3280 5256
rect 3881 5253 3893 5256
rect 3927 5284 3939 5287
rect 4062 5284 4068 5296
rect 3927 5256 4068 5284
rect 3927 5253 3939 5256
rect 3881 5247 3939 5253
rect 4062 5244 4068 5256
rect 4120 5244 4126 5296
rect 4617 5287 4675 5293
rect 4617 5253 4629 5287
rect 4663 5284 4675 5287
rect 4706 5284 4712 5296
rect 4663 5256 4712 5284
rect 4663 5253 4675 5256
rect 4617 5247 4675 5253
rect 4706 5244 4712 5256
rect 4764 5244 4770 5296
rect 8754 5284 8760 5296
rect 8602 5256 8760 5284
rect 8754 5244 8760 5256
rect 8812 5284 8818 5296
rect 9950 5284 9956 5296
rect 8812 5256 9956 5284
rect 8812 5244 8818 5256
rect 9950 5244 9956 5256
rect 10008 5244 10014 5296
rect 10778 5284 10784 5296
rect 10718 5256 10784 5284
rect 10778 5244 10784 5256
rect 10836 5244 10842 5296
rect 12084 5293 12112 5324
rect 12069 5287 12127 5293
rect 12069 5253 12081 5287
rect 12115 5253 12127 5287
rect 12069 5247 12127 5253
rect 3237 5219 3295 5225
rect 3237 5185 3249 5219
rect 3283 5185 3295 5219
rect 3237 5179 3295 5185
rect 3326 5176 3332 5228
rect 3384 5216 3390 5228
rect 3605 5219 3663 5225
rect 3605 5216 3617 5219
rect 3384 5188 3617 5216
rect 3384 5176 3390 5188
rect 3605 5185 3617 5188
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 3789 5219 3847 5225
rect 3789 5185 3801 5219
rect 3835 5216 3847 5219
rect 3835 5188 3924 5216
rect 3835 5185 3847 5188
rect 3789 5179 3847 5185
rect 2958 5108 2964 5160
rect 3016 5108 3022 5160
rect 3896 5092 3924 5188
rect 3970 5176 3976 5228
rect 4028 5225 4034 5228
rect 4028 5216 4036 5225
rect 4028 5188 4073 5216
rect 4028 5179 4036 5188
rect 4028 5176 4034 5179
rect 5718 5176 5724 5228
rect 5776 5216 5782 5228
rect 5776 5188 6960 5216
rect 5776 5176 5782 5188
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 6365 5151 6423 5157
rect 6365 5148 6377 5151
rect 4341 5111 4399 5117
rect 4448 5120 6377 5148
rect 3878 5040 3884 5092
rect 3936 5040 3942 5092
rect 4157 5083 4215 5089
rect 4157 5049 4169 5083
rect 4203 5080 4215 5083
rect 4356 5080 4384 5111
rect 4203 5052 4384 5080
rect 4203 5049 4215 5052
rect 4157 5043 4215 5049
rect 3421 5015 3479 5021
rect 3421 4981 3433 5015
rect 3467 5012 3479 5015
rect 3786 5012 3792 5024
rect 3467 4984 3792 5012
rect 3467 4981 3479 4984
rect 3421 4975 3479 4981
rect 3786 4972 3792 4984
rect 3844 4972 3850 5024
rect 4062 4972 4068 5024
rect 4120 5012 4126 5024
rect 4448 5012 4476 5120
rect 6365 5117 6377 5120
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 6641 5083 6699 5089
rect 6641 5080 6653 5083
rect 6380 5052 6653 5080
rect 6380 5024 6408 5052
rect 6641 5049 6653 5052
rect 6687 5049 6699 5083
rect 6641 5043 6699 5049
rect 4120 4984 4476 5012
rect 4120 4972 4126 4984
rect 6362 4972 6368 5024
rect 6420 4972 6426 5024
rect 6730 4972 6736 5024
rect 6788 5012 6794 5024
rect 6825 5015 6883 5021
rect 6825 5012 6837 5015
rect 6788 4984 6837 5012
rect 6788 4972 6794 4984
rect 6825 4981 6837 4984
rect 6871 4981 6883 5015
rect 6932 5012 6960 5188
rect 7098 5176 7104 5228
rect 7156 5176 7162 5228
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 12452 5225 12480 5324
rect 15105 5321 15117 5324
rect 15151 5321 15163 5355
rect 15105 5315 15163 5321
rect 12526 5244 12532 5296
rect 12584 5284 12590 5296
rect 12713 5287 12771 5293
rect 12713 5284 12725 5287
rect 12584 5256 12725 5284
rect 12584 5244 12590 5256
rect 12713 5253 12725 5256
rect 12759 5284 12771 5287
rect 13538 5284 13544 5296
rect 12759 5256 13544 5284
rect 12759 5253 12771 5256
rect 12713 5247 12771 5253
rect 13538 5244 13544 5256
rect 13596 5244 13602 5296
rect 14918 5284 14924 5296
rect 14858 5256 14924 5284
rect 14918 5244 14924 5256
rect 14976 5244 14982 5296
rect 9217 5219 9275 5225
rect 9217 5216 9229 5219
rect 9088 5188 9229 5216
rect 9088 5176 9094 5188
rect 9217 5185 9229 5188
rect 9263 5185 9275 5219
rect 12345 5219 12403 5225
rect 12345 5216 12357 5219
rect 9217 5179 9275 5185
rect 11256 5188 12357 5216
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 7742 5148 7748 5160
rect 7423 5120 7748 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 7742 5108 7748 5120
rect 7800 5108 7806 5160
rect 9493 5151 9551 5157
rect 9493 5117 9505 5151
rect 9539 5148 9551 5151
rect 10042 5148 10048 5160
rect 9539 5120 10048 5148
rect 9539 5117 9551 5120
rect 9493 5111 9551 5117
rect 10042 5108 10048 5120
rect 10100 5108 10106 5160
rect 10134 5108 10140 5160
rect 10192 5148 10198 5160
rect 11256 5148 11284 5188
rect 12345 5185 12357 5188
rect 12391 5185 12403 5219
rect 12345 5179 12403 5185
rect 12437 5219 12495 5225
rect 12437 5185 12449 5219
rect 12483 5185 12495 5219
rect 12437 5179 12495 5185
rect 10192 5120 11284 5148
rect 12360 5148 12388 5179
rect 12618 5176 12624 5228
rect 12676 5176 12682 5228
rect 12810 5219 12868 5225
rect 12810 5185 12822 5219
rect 12856 5185 12868 5219
rect 12810 5179 12868 5185
rect 12820 5148 12848 5179
rect 13078 5176 13084 5228
rect 13136 5216 13142 5228
rect 13357 5219 13415 5225
rect 13357 5216 13369 5219
rect 13136 5188 13369 5216
rect 13136 5176 13142 5188
rect 13357 5185 13369 5188
rect 13403 5185 13415 5219
rect 13357 5179 13415 5185
rect 12360 5120 12848 5148
rect 10192 5108 10198 5120
rect 13630 5108 13636 5160
rect 13688 5108 13694 5160
rect 11698 5040 11704 5092
rect 11756 5040 11762 5092
rect 9306 5012 9312 5024
rect 6932 4984 9312 5012
rect 6825 4975 6883 4981
rect 9306 4972 9312 4984
rect 9364 4972 9370 5024
rect 11606 4972 11612 5024
rect 11664 4972 11670 5024
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 12253 5015 12311 5021
rect 12253 5012 12265 5015
rect 11848 4984 12265 5012
rect 11848 4972 11854 4984
rect 12253 4981 12265 4984
rect 12299 4981 12311 5015
rect 12253 4975 12311 4981
rect 12989 5015 13047 5021
rect 12989 4981 13001 5015
rect 13035 5012 13047 5015
rect 13446 5012 13452 5024
rect 13035 4984 13452 5012
rect 13035 4981 13047 4984
rect 12989 4975 13047 4981
rect 13446 4972 13452 4984
rect 13504 4972 13510 5024
rect 1104 4922 22816 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 20214 4922
rect 20266 4870 20278 4922
rect 20330 4870 20342 4922
rect 20394 4870 20406 4922
rect 20458 4870 20470 4922
rect 20522 4870 22816 4922
rect 1104 4848 22816 4870
rect 3878 4768 3884 4820
rect 3936 4808 3942 4820
rect 5537 4811 5595 4817
rect 5537 4808 5549 4811
rect 3936 4780 5549 4808
rect 3936 4768 3942 4780
rect 5537 4777 5549 4780
rect 5583 4808 5595 4811
rect 5994 4808 6000 4820
rect 5583 4780 6000 4808
rect 5583 4777 5595 4780
rect 5537 4771 5595 4777
rect 5994 4768 6000 4780
rect 6052 4768 6058 4820
rect 6638 4768 6644 4820
rect 6696 4808 6702 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 6696 4780 8125 4808
rect 6696 4768 6702 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 8113 4771 8171 4777
rect 12332 4811 12390 4817
rect 12332 4777 12344 4811
rect 12378 4808 12390 4811
rect 12710 4808 12716 4820
rect 12378 4780 12716 4808
rect 12378 4777 12390 4780
rect 12332 4771 12390 4777
rect 12710 4768 12716 4780
rect 12768 4768 12774 4820
rect 13630 4768 13636 4820
rect 13688 4808 13694 4820
rect 13817 4811 13875 4817
rect 13817 4808 13829 4811
rect 13688 4780 13829 4808
rect 13688 4768 13694 4780
rect 13817 4777 13829 4780
rect 13863 4777 13875 4811
rect 13817 4771 13875 4777
rect 3513 4743 3571 4749
rect 3513 4709 3525 4743
rect 3559 4740 3571 4743
rect 3559 4712 3924 4740
rect 3559 4709 3571 4712
rect 3513 4703 3571 4709
rect 1765 4675 1823 4681
rect 1765 4641 1777 4675
rect 1811 4672 1823 4675
rect 3326 4672 3332 4684
rect 1811 4644 3332 4672
rect 1811 4641 1823 4644
rect 1765 4635 1823 4641
rect 3326 4632 3332 4644
rect 3384 4632 3390 4684
rect 3786 4632 3792 4684
rect 3844 4632 3850 4684
rect 3896 4672 3924 4712
rect 7742 4700 7748 4752
rect 7800 4700 7806 4752
rect 9125 4743 9183 4749
rect 9125 4740 9137 4743
rect 7852 4712 9137 4740
rect 4065 4675 4123 4681
rect 4065 4672 4077 4675
rect 3896 4644 4077 4672
rect 4065 4641 4077 4644
rect 4111 4641 4123 4675
rect 4065 4635 4123 4641
rect 5534 4632 5540 4684
rect 5592 4672 5598 4684
rect 5997 4675 6055 4681
rect 5997 4672 6009 4675
rect 5592 4644 6009 4672
rect 5592 4632 5598 4644
rect 5997 4641 6009 4644
rect 6043 4641 6055 4675
rect 5997 4635 6055 4641
rect 6270 4632 6276 4684
rect 6328 4632 6334 4684
rect 3142 4564 3148 4616
rect 3200 4604 3206 4616
rect 3200 4576 3832 4604
rect 3200 4564 3206 4576
rect 2038 4496 2044 4548
rect 2096 4496 2102 4548
rect 3804 4536 3832 4576
rect 5902 4564 5908 4616
rect 5960 4564 5966 4616
rect 3804 4508 4554 4536
rect 5368 4508 5948 4536
rect 4448 4480 4476 4508
rect 4430 4428 4436 4480
rect 4488 4428 4494 4480
rect 4706 4428 4712 4480
rect 4764 4468 4770 4480
rect 5368 4468 5396 4508
rect 4764 4440 5396 4468
rect 4764 4428 4770 4440
rect 5810 4428 5816 4480
rect 5868 4428 5874 4480
rect 5920 4468 5948 4508
rect 6822 4496 6828 4548
rect 6880 4496 6886 4548
rect 7852 4468 7880 4712
rect 9125 4709 9137 4712
rect 9171 4709 9183 4743
rect 9125 4703 9183 4709
rect 10413 4675 10471 4681
rect 8404 4644 9628 4672
rect 8110 4564 8116 4616
rect 8168 4604 8174 4616
rect 8404 4613 8432 4644
rect 9600 4616 9628 4644
rect 10413 4641 10425 4675
rect 10459 4672 10471 4675
rect 11606 4672 11612 4684
rect 10459 4644 11612 4672
rect 10459 4641 10471 4644
rect 10413 4635 10471 4641
rect 11606 4632 11612 4644
rect 11664 4632 11670 4684
rect 12069 4675 12127 4681
rect 12069 4641 12081 4675
rect 12115 4672 12127 4675
rect 12710 4672 12716 4684
rect 12115 4644 12716 4672
rect 12115 4641 12127 4644
rect 12069 4635 12127 4641
rect 12710 4632 12716 4644
rect 12768 4672 12774 4684
rect 13354 4672 13360 4684
rect 12768 4644 13360 4672
rect 12768 4632 12774 4644
rect 13354 4632 13360 4644
rect 13412 4632 13418 4684
rect 8251 4607 8309 4613
rect 8251 4604 8263 4607
rect 8168 4576 8263 4604
rect 8168 4564 8174 4576
rect 8251 4573 8263 4576
rect 8297 4573 8309 4607
rect 8251 4567 8309 4573
rect 8389 4607 8447 4613
rect 8389 4573 8401 4607
rect 8435 4573 8447 4607
rect 8389 4567 8447 4573
rect 8665 4607 8723 4613
rect 8665 4573 8677 4607
rect 8711 4604 8723 4607
rect 9214 4604 9220 4616
rect 8711 4576 9220 4604
rect 8711 4573 8723 4576
rect 8665 4567 8723 4573
rect 9214 4564 9220 4576
rect 9272 4604 9278 4616
rect 9493 4607 9551 4613
rect 9493 4604 9505 4607
rect 9272 4576 9505 4604
rect 9272 4564 9278 4576
rect 9493 4573 9505 4576
rect 9539 4573 9551 4607
rect 9493 4567 9551 4573
rect 9582 4564 9588 4616
rect 9640 4604 9646 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 9640 4576 9781 4604
rect 9640 4564 9646 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 10134 4564 10140 4616
rect 10192 4564 10198 4616
rect 14274 4564 14280 4616
rect 14332 4564 14338 4616
rect 8481 4539 8539 4545
rect 8481 4505 8493 4539
rect 8527 4536 8539 4539
rect 8754 4536 8760 4548
rect 8527 4508 8760 4536
rect 8527 4505 8539 4508
rect 8481 4499 8539 4505
rect 8754 4496 8760 4508
rect 8812 4496 8818 4548
rect 10870 4496 10876 4548
rect 10928 4496 10934 4548
rect 13078 4496 13084 4548
rect 13136 4496 13142 4548
rect 5920 4440 7880 4468
rect 8846 4428 8852 4480
rect 8904 4468 8910 4480
rect 9033 4471 9091 4477
rect 9033 4468 9045 4471
rect 8904 4440 9045 4468
rect 8904 4428 8910 4440
rect 9033 4437 9045 4440
rect 9079 4437 9091 4471
rect 9033 4431 9091 4437
rect 9674 4428 9680 4480
rect 9732 4428 9738 4480
rect 11885 4471 11943 4477
rect 11885 4437 11897 4471
rect 11931 4468 11943 4471
rect 12066 4468 12072 4480
rect 11931 4440 12072 4468
rect 11931 4437 11943 4440
rect 11885 4431 11943 4437
rect 12066 4428 12072 4440
rect 12124 4428 12130 4480
rect 14090 4428 14096 4480
rect 14148 4468 14154 4480
rect 14185 4471 14243 4477
rect 14185 4468 14197 4471
rect 14148 4440 14197 4468
rect 14148 4428 14154 4440
rect 14185 4437 14197 4440
rect 14231 4437 14243 4471
rect 14185 4431 14243 4437
rect 1104 4378 22816 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 22816 4378
rect 1104 4304 22816 4326
rect 1581 4267 1639 4273
rect 1581 4233 1593 4267
rect 1627 4264 1639 4267
rect 2038 4264 2044 4276
rect 1627 4236 2044 4264
rect 1627 4233 1639 4236
rect 1581 4227 1639 4233
rect 2038 4224 2044 4236
rect 2096 4224 2102 4276
rect 2958 4224 2964 4276
rect 3016 4264 3022 4276
rect 5905 4267 5963 4273
rect 5905 4264 5917 4267
rect 3016 4236 5917 4264
rect 3016 4224 3022 4236
rect 5905 4233 5917 4236
rect 5951 4233 5963 4267
rect 5905 4227 5963 4233
rect 9048 4236 9996 4264
rect 4157 4199 4215 4205
rect 4157 4196 4169 4199
rect 2884 4168 4169 4196
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2130 4128 2136 4140
rect 2087 4100 2136 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2130 4088 2136 4100
rect 2188 4088 2194 4140
rect 2884 4128 2912 4168
rect 4157 4165 4169 4168
rect 4203 4165 4215 4199
rect 4157 4159 4215 4165
rect 4430 4156 4436 4208
rect 4488 4196 4494 4208
rect 4488 4168 4646 4196
rect 4488 4156 4494 4168
rect 5534 4156 5540 4208
rect 5592 4196 5598 4208
rect 6730 4196 6736 4208
rect 5592 4168 6736 4196
rect 5592 4156 5598 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 9048 4196 9076 4236
rect 9968 4208 9996 4236
rect 10042 4224 10048 4276
rect 10100 4264 10106 4276
rect 10137 4267 10195 4273
rect 10137 4264 10149 4267
rect 10100 4236 10149 4264
rect 10100 4224 10106 4236
rect 10137 4233 10149 4236
rect 10183 4233 10195 4267
rect 10137 4227 10195 4233
rect 13538 4224 13544 4276
rect 13596 4224 13602 4276
rect 9950 4196 9956 4208
rect 7958 4168 9076 4196
rect 9890 4168 9956 4196
rect 9950 4156 9956 4168
rect 10008 4196 10014 4208
rect 10778 4196 10784 4208
rect 10008 4168 10784 4196
rect 10008 4156 10014 4168
rect 10778 4156 10784 4168
rect 10836 4156 10842 4208
rect 12066 4156 12072 4208
rect 12124 4156 12130 4208
rect 3050 4137 3056 4140
rect 2240 4100 2912 4128
rect 2240 4001 2268 4100
rect 3048 4091 3056 4137
rect 3050 4088 3056 4091
rect 3108 4088 3114 4140
rect 3145 4131 3203 4137
rect 3145 4097 3157 4131
rect 3191 4097 3203 4131
rect 3145 4091 3203 4097
rect 3237 4131 3295 4137
rect 3237 4097 3249 4131
rect 3283 4097 3295 4131
rect 3237 4091 3295 4097
rect 3421 4131 3479 4137
rect 3421 4097 3433 4131
rect 3467 4126 3479 4131
rect 3510 4126 3516 4140
rect 3467 4098 3516 4126
rect 3467 4097 3479 4098
rect 3421 4091 3479 4097
rect 2685 4063 2743 4069
rect 2685 4029 2697 4063
rect 2731 4060 2743 4063
rect 2774 4060 2780 4072
rect 2731 4032 2780 4060
rect 2731 4029 2743 4032
rect 2685 4023 2743 4029
rect 2774 4020 2780 4032
rect 2832 4020 2838 4072
rect 2958 4020 2964 4072
rect 3016 4060 3022 4072
rect 3160 4060 3188 4091
rect 3016 4032 3188 4060
rect 3252 4060 3280 4091
rect 3510 4088 3516 4098
rect 3568 4088 3574 4140
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 3878 4128 3884 4140
rect 3752 4100 3884 4128
rect 3752 4088 3758 4100
rect 3878 4088 3884 4100
rect 3936 4088 3942 4140
rect 5813 4131 5871 4137
rect 5813 4097 5825 4131
rect 5859 4097 5871 4131
rect 5813 4091 5871 4097
rect 3602 4060 3608 4072
rect 3252 4032 3608 4060
rect 3016 4020 3022 4032
rect 3602 4020 3608 4032
rect 3660 4020 3666 4072
rect 5828 4060 5856 4091
rect 5994 4088 6000 4140
rect 6052 4088 6058 4140
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 10321 4131 10379 4137
rect 10321 4097 10333 4131
rect 10367 4097 10379 4131
rect 10321 4091 10379 4097
rect 3804 4032 5856 4060
rect 6457 4063 6515 4069
rect 1765 3995 1823 4001
rect 1765 3961 1777 3995
rect 1811 3961 1823 3995
rect 1765 3955 1823 3961
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3961 2283 3995
rect 2225 3955 2283 3961
rect 1302 3884 1308 3936
rect 1360 3924 1366 3936
rect 1780 3924 1808 3955
rect 2406 3952 2412 4004
rect 2464 3952 2470 4004
rect 2869 3995 2927 4001
rect 2869 3961 2881 3995
rect 2915 3992 2927 3995
rect 3234 3992 3240 4004
rect 2915 3964 3240 3992
rect 2915 3961 2927 3964
rect 2869 3955 2927 3961
rect 3234 3952 3240 3964
rect 3292 3952 3298 4004
rect 3804 3992 3832 4032
rect 6457 4029 6469 4063
rect 6503 4029 6515 4063
rect 6457 4023 6515 4029
rect 3528 3964 3832 3992
rect 3528 3924 3556 3964
rect 1360 3896 3556 3924
rect 1360 3884 1366 3896
rect 3602 3884 3608 3936
rect 3660 3884 3666 3936
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5316 3896 5641 3924
rect 5316 3884 5322 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 6472 3924 6500 4023
rect 6730 4020 6736 4072
rect 6788 4020 6794 4072
rect 8662 4020 8668 4072
rect 8720 4020 8726 4072
rect 8754 4020 8760 4072
rect 8812 4060 8818 4072
rect 10336 4060 10364 4091
rect 11790 4088 11796 4140
rect 11848 4088 11854 4140
rect 13078 4088 13084 4140
rect 13136 4128 13142 4140
rect 13136 4114 13202 4128
rect 13136 4100 13216 4114
rect 13136 4088 13142 4100
rect 8812 4032 10364 4060
rect 8812 4020 8818 4032
rect 10410 4020 10416 4072
rect 10468 4020 10474 4072
rect 13188 4060 13216 4100
rect 13906 4088 13912 4140
rect 13964 4088 13970 4140
rect 13262 4060 13268 4072
rect 13188 4032 13268 4060
rect 13262 4020 13268 4032
rect 13320 4060 13326 4072
rect 14918 4060 14924 4072
rect 13320 4032 14924 4060
rect 13320 4020 13326 4032
rect 14918 4020 14924 4032
rect 14976 4060 14982 4072
rect 15654 4060 15660 4072
rect 14976 4032 15660 4060
rect 14976 4020 14982 4032
rect 15654 4020 15660 4032
rect 15712 4020 15718 4072
rect 7760 3964 8340 3992
rect 6914 3924 6920 3936
rect 6472 3896 6920 3924
rect 5629 3887 5687 3893
rect 6914 3884 6920 3896
rect 6972 3924 6978 3936
rect 7760 3924 7788 3964
rect 6972 3896 7788 3924
rect 6972 3884 6978 3896
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8205 3927 8263 3933
rect 8205 3924 8217 3927
rect 8168 3896 8217 3924
rect 8168 3884 8174 3896
rect 8205 3893 8217 3896
rect 8251 3893 8263 3927
rect 8312 3924 8340 3964
rect 10042 3952 10048 4004
rect 10100 3992 10106 4004
rect 10428 3992 10456 4020
rect 10962 3992 10968 4004
rect 10100 3964 10968 3992
rect 10100 3952 10106 3964
rect 10962 3952 10968 3964
rect 11020 3952 11026 4004
rect 8754 3924 8760 3936
rect 8312 3896 8760 3924
rect 8205 3887 8263 3893
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 10410 3884 10416 3936
rect 10468 3884 10474 3936
rect 1104 3834 22816 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 20214 3834
rect 20266 3782 20278 3834
rect 20330 3782 20342 3834
rect 20394 3782 20406 3834
rect 20458 3782 20470 3834
rect 20522 3782 22816 3834
rect 1104 3760 22816 3782
rect 2774 3680 2780 3732
rect 2832 3720 2838 3732
rect 2832 3692 3280 3720
rect 2832 3680 2838 3692
rect 3252 3652 3280 3692
rect 3326 3680 3332 3732
rect 3384 3720 3390 3732
rect 3881 3723 3939 3729
rect 3881 3720 3893 3723
rect 3384 3692 3893 3720
rect 3384 3680 3390 3692
rect 3881 3689 3893 3692
rect 3927 3689 3939 3723
rect 6730 3720 6736 3732
rect 3881 3683 3939 3689
rect 4816 3692 6736 3720
rect 4522 3652 4528 3664
rect 3252 3624 4528 3652
rect 4522 3612 4528 3624
rect 4580 3612 4586 3664
rect 4816 3661 4844 3692
rect 6730 3680 6736 3692
rect 6788 3680 6794 3732
rect 9030 3720 9036 3732
rect 7024 3692 9036 3720
rect 4801 3655 4859 3661
rect 4801 3621 4813 3655
rect 4847 3621 4859 3655
rect 7024 3652 7052 3692
rect 9030 3680 9036 3692
rect 9088 3680 9094 3732
rect 9490 3680 9496 3732
rect 9548 3720 9554 3732
rect 11241 3723 11299 3729
rect 11241 3720 11253 3723
rect 9548 3692 11253 3720
rect 9548 3680 9554 3692
rect 11241 3689 11253 3692
rect 11287 3689 11299 3723
rect 11241 3683 11299 3689
rect 4801 3615 4859 3621
rect 6748 3624 7052 3652
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 1627 3556 1777 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1765 3553 1777 3556
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 3050 3544 3056 3596
rect 3108 3584 3114 3596
rect 3513 3587 3571 3593
rect 3513 3584 3525 3587
rect 3108 3556 3525 3584
rect 3108 3544 3114 3556
rect 3513 3553 3525 3556
rect 3559 3553 3571 3587
rect 3513 3547 3571 3553
rect 1673 3519 1731 3525
rect 1673 3485 1685 3519
rect 1719 3485 1731 3519
rect 1673 3479 1731 3485
rect 1688 3380 1716 3479
rect 3142 3476 3148 3528
rect 3200 3476 3206 3528
rect 3418 3476 3424 3528
rect 3476 3516 3482 3528
rect 3528 3516 3556 3547
rect 3878 3544 3884 3596
rect 3936 3584 3942 3596
rect 4706 3584 4712 3596
rect 3936 3556 4476 3584
rect 3936 3544 3942 3556
rect 4448 3525 4476 3556
rect 4540 3556 4712 3584
rect 4540 3525 4568 3556
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 4985 3587 5043 3593
rect 4985 3553 4997 3587
rect 5031 3584 5043 3587
rect 5810 3584 5816 3596
rect 5031 3556 5816 3584
rect 5031 3553 5043 3556
rect 4985 3547 5043 3553
rect 5810 3544 5816 3556
rect 5868 3544 5874 3596
rect 6546 3544 6552 3596
rect 6604 3584 6610 3596
rect 6748 3593 6776 3624
rect 10962 3612 10968 3664
rect 11020 3652 11026 3664
rect 11609 3655 11667 3661
rect 11609 3652 11621 3655
rect 11020 3624 11621 3652
rect 11020 3612 11026 3624
rect 11609 3621 11621 3624
rect 11655 3621 11667 3655
rect 11609 3615 11667 3621
rect 6733 3587 6791 3593
rect 6733 3584 6745 3587
rect 6604 3556 6745 3584
rect 6604 3544 6610 3556
rect 6733 3553 6745 3556
rect 6779 3553 6791 3587
rect 6733 3547 6791 3553
rect 6917 3587 6975 3593
rect 6917 3553 6929 3587
rect 6963 3584 6975 3587
rect 8570 3584 8576 3596
rect 6963 3556 8576 3584
rect 6963 3553 6975 3556
rect 6917 3547 6975 3553
rect 8570 3544 8576 3556
rect 8628 3544 8634 3596
rect 8665 3587 8723 3593
rect 8665 3553 8677 3587
rect 8711 3584 8723 3587
rect 9769 3587 9827 3593
rect 9769 3584 9781 3587
rect 8711 3556 9781 3584
rect 8711 3553 8723 3556
rect 8665 3547 8723 3553
rect 9769 3553 9781 3556
rect 9815 3553 9827 3587
rect 9769 3547 9827 3553
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 12069 3587 12127 3593
rect 12069 3584 12081 3587
rect 11940 3556 12081 3584
rect 11940 3544 11946 3556
rect 12069 3553 12081 3556
rect 12115 3584 12127 3587
rect 12115 3556 13952 3584
rect 12115 3553 12127 3556
rect 12069 3547 12127 3553
rect 4013 3519 4071 3525
rect 4013 3516 4025 3519
rect 3476 3488 4025 3516
rect 3476 3476 3482 3488
rect 4013 3485 4025 3488
rect 4059 3485 4071 3519
rect 4013 3479 4071 3485
rect 4157 3519 4215 3525
rect 4157 3485 4169 3519
rect 4203 3516 4215 3519
rect 4433 3519 4491 3525
rect 4203 3488 4384 3516
rect 4203 3485 4215 3488
rect 4157 3479 4215 3485
rect 2038 3408 2044 3460
rect 2096 3408 2102 3460
rect 4172 3448 4200 3479
rect 3344 3420 4200 3448
rect 4249 3451 4307 3457
rect 2958 3380 2964 3392
rect 1688 3352 2964 3380
rect 2958 3340 2964 3352
rect 3016 3380 3022 3392
rect 3344 3380 3372 3420
rect 4249 3417 4261 3451
rect 4295 3417 4307 3451
rect 4356 3448 4384 3488
rect 4433 3485 4445 3519
rect 4479 3485 4491 3519
rect 4433 3479 4491 3485
rect 4525 3519 4583 3525
rect 4525 3485 4537 3519
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4798 3476 4804 3528
rect 4856 3476 4862 3528
rect 8938 3476 8944 3528
rect 8996 3476 9002 3528
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 9088 3488 9137 3516
rect 9088 3476 9094 3488
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9493 3519 9551 3525
rect 9493 3485 9505 3519
rect 9539 3485 9551 3519
rect 9493 3479 9551 3485
rect 4614 3448 4620 3460
rect 4356 3420 4620 3448
rect 4249 3411 4307 3417
rect 3016 3352 3372 3380
rect 3016 3340 3022 3352
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 4264 3380 4292 3411
rect 4614 3408 4620 3420
rect 4672 3408 4678 3460
rect 5258 3408 5264 3460
rect 5316 3408 5322 3460
rect 6822 3448 6828 3460
rect 6486 3420 6828 3448
rect 5442 3380 5448 3392
rect 3752 3352 5448 3380
rect 3752 3340 3758 3352
rect 5442 3340 5448 3352
rect 5500 3340 5506 3392
rect 5626 3340 5632 3392
rect 5684 3380 5690 3392
rect 6564 3380 6592 3420
rect 6822 3408 6828 3420
rect 6880 3408 6886 3460
rect 7193 3451 7251 3457
rect 7193 3417 7205 3451
rect 7239 3417 7251 3451
rect 8662 3448 8668 3460
rect 8418 3420 8668 3448
rect 7193 3411 7251 3417
rect 5684 3352 6592 3380
rect 7208 3380 7236 3411
rect 8662 3408 8668 3420
rect 8720 3448 8726 3460
rect 9508 3448 9536 3479
rect 9674 3448 9680 3460
rect 8720 3420 9449 3448
rect 9508 3420 9680 3448
rect 8720 3408 8726 3420
rect 8846 3380 8852 3392
rect 7208 3352 8852 3380
rect 5684 3340 5690 3352
rect 8846 3340 8852 3352
rect 8904 3340 8910 3392
rect 8938 3340 8944 3392
rect 8996 3380 9002 3392
rect 9033 3383 9091 3389
rect 9033 3380 9045 3383
rect 8996 3352 9045 3380
rect 8996 3340 9002 3352
rect 9033 3349 9045 3352
rect 9079 3349 9091 3383
rect 9421 3380 9449 3420
rect 9674 3408 9680 3420
rect 9732 3408 9738 3460
rect 10778 3408 10784 3460
rect 10836 3408 10842 3460
rect 11974 3408 11980 3460
rect 12032 3408 12038 3460
rect 12345 3451 12403 3457
rect 12345 3417 12357 3451
rect 12391 3417 12403 3451
rect 12345 3411 12403 3417
rect 9950 3380 9956 3392
rect 9421 3352 9956 3380
rect 9033 3343 9091 3349
rect 9950 3340 9956 3352
rect 10008 3340 10014 3392
rect 11517 3383 11575 3389
rect 11517 3349 11529 3383
rect 11563 3380 11575 3383
rect 12360 3380 12388 3411
rect 13078 3408 13084 3460
rect 13136 3408 13142 3460
rect 13924 3448 13952 3556
rect 14090 3544 14096 3596
rect 14148 3544 14154 3596
rect 14274 3448 14280 3460
rect 13924 3420 14280 3448
rect 14274 3408 14280 3420
rect 14332 3408 14338 3460
rect 14369 3451 14427 3457
rect 14369 3417 14381 3451
rect 14415 3417 14427 3451
rect 15654 3448 15660 3460
rect 15594 3420 15660 3448
rect 14369 3411 14427 3417
rect 11563 3352 12388 3380
rect 13817 3383 13875 3389
rect 11563 3349 11575 3352
rect 11517 3343 11575 3349
rect 13817 3349 13829 3383
rect 13863 3380 13875 3383
rect 14384 3380 14412 3411
rect 15654 3408 15660 3420
rect 15712 3408 15718 3460
rect 13863 3352 14412 3380
rect 13863 3349 13875 3352
rect 13817 3343 13875 3349
rect 15838 3340 15844 3392
rect 15896 3340 15902 3392
rect 1104 3290 22816 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 22816 3290
rect 1104 3216 22816 3238
rect 1486 3136 1492 3188
rect 1544 3176 1550 3188
rect 6089 3179 6147 3185
rect 1544 3148 4016 3176
rect 1544 3136 1550 3148
rect 2774 3108 2780 3120
rect 2622 3080 2780 3108
rect 2774 3068 2780 3080
rect 2832 3108 2838 3120
rect 3142 3108 3148 3120
rect 2832 3080 3148 3108
rect 2832 3068 2838 3080
rect 3142 3068 3148 3080
rect 3200 3068 3206 3120
rect 3694 3049 3700 3052
rect 3692 3003 3700 3049
rect 3694 3000 3700 3003
rect 3752 3000 3758 3052
rect 3786 3000 3792 3052
rect 3844 3000 3850 3052
rect 3881 3043 3939 3049
rect 3881 3009 3893 3043
rect 3927 3040 3939 3043
rect 3988 3040 4016 3148
rect 6089 3145 6101 3179
rect 6135 3176 6147 3179
rect 6135 3148 6776 3176
rect 6135 3145 6147 3148
rect 6089 3139 6147 3145
rect 4706 3068 4712 3120
rect 4764 3108 4770 3120
rect 6748 3117 6776 3148
rect 6822 3136 6828 3188
rect 6880 3176 6886 3188
rect 8205 3179 8263 3185
rect 8205 3176 8217 3179
rect 6880 3148 8217 3176
rect 6880 3136 6886 3148
rect 8205 3145 8217 3148
rect 8251 3145 8263 3179
rect 8205 3139 8263 3145
rect 8570 3136 8576 3188
rect 8628 3176 8634 3188
rect 9582 3176 9588 3188
rect 8628 3148 9588 3176
rect 8628 3136 8634 3148
rect 9582 3136 9588 3148
rect 9640 3176 9646 3188
rect 15838 3176 15844 3188
rect 9640 3148 10548 3176
rect 9640 3136 9646 3148
rect 6733 3111 6791 3117
rect 4764 3080 5106 3108
rect 4764 3068 4770 3080
rect 6733 3077 6745 3111
rect 6779 3077 6791 3111
rect 8294 3108 8300 3120
rect 7958 3080 8300 3108
rect 6733 3071 6791 3077
rect 8294 3068 8300 3080
rect 8352 3108 8358 3120
rect 8662 3108 8668 3120
rect 8352 3080 8668 3108
rect 8352 3068 8358 3080
rect 8662 3068 8668 3080
rect 8720 3068 8726 3120
rect 9950 3108 9956 3120
rect 9522 3080 9956 3108
rect 9950 3068 9956 3080
rect 10008 3068 10014 3120
rect 10410 3108 10416 3120
rect 10244 3080 10416 3108
rect 3927 3012 4016 3040
rect 3927 3009 3939 3012
rect 3881 3003 3939 3009
rect 4062 3000 4068 3052
rect 4120 3000 4126 3052
rect 10244 3049 10272 3080
rect 10410 3068 10416 3080
rect 10468 3068 10474 3120
rect 10229 3043 10287 3049
rect 10229 3009 10241 3043
rect 10275 3009 10287 3043
rect 10229 3003 10287 3009
rect 10321 3043 10379 3049
rect 10321 3009 10333 3043
rect 10367 3040 10379 3043
rect 10520 3040 10548 3148
rect 12406 3148 15844 3176
rect 12406 3108 12434 3148
rect 11348 3080 12434 3108
rect 10367 3012 10548 3040
rect 10367 3009 10379 3012
rect 10321 3003 10379 3009
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11348 3049 11376 3080
rect 14274 3068 14280 3120
rect 14332 3108 14338 3120
rect 15013 3111 15071 3117
rect 15013 3108 15025 3111
rect 14332 3080 15025 3108
rect 14332 3068 14338 3080
rect 15013 3077 15025 3080
rect 15059 3077 15071 3111
rect 15013 3071 15071 3077
rect 11057 3043 11115 3049
rect 11057 3040 11069 3043
rect 11020 3012 11069 3040
rect 11020 3000 11026 3012
rect 11057 3009 11069 3012
rect 11103 3009 11115 3043
rect 11057 3003 11115 3009
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3009 11391 3043
rect 11333 3003 11391 3009
rect 11514 3000 11520 3052
rect 11572 3040 11578 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11572 3012 11621 3040
rect 11572 3000 11578 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11609 3003 11667 3009
rect 13262 3000 13268 3052
rect 13320 3000 13326 3052
rect 14777 3043 14835 3049
rect 14777 3040 14789 3043
rect 13464 3012 14789 3040
rect 1581 2975 1639 2981
rect 1581 2941 1593 2975
rect 1627 2972 1639 2975
rect 2038 2972 2044 2984
rect 1627 2944 2044 2972
rect 1627 2941 1639 2944
rect 1581 2935 1639 2941
rect 2038 2932 2044 2944
rect 2096 2932 2102 2984
rect 3050 2932 3056 2984
rect 3108 2932 3114 2984
rect 3329 2975 3387 2981
rect 3329 2941 3341 2975
rect 3375 2972 3387 2975
rect 3375 2944 4108 2972
rect 3375 2941 3387 2944
rect 3329 2935 3387 2941
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 3878 2836 3884 2848
rect 3568 2808 3884 2836
rect 3568 2796 3574 2808
rect 3878 2796 3884 2808
rect 3936 2796 3942 2848
rect 4080 2836 4108 2944
rect 4154 2932 4160 2984
rect 4212 2972 4218 2984
rect 4341 2975 4399 2981
rect 4341 2972 4353 2975
rect 4212 2944 4353 2972
rect 4212 2932 4218 2944
rect 4341 2941 4353 2944
rect 4387 2941 4399 2975
rect 4341 2935 4399 2941
rect 4617 2975 4675 2981
rect 4617 2941 4629 2975
rect 4663 2972 4675 2975
rect 4663 2944 6408 2972
rect 4663 2941 4675 2944
rect 4617 2935 4675 2941
rect 6380 2904 6408 2944
rect 6454 2932 6460 2984
rect 6512 2932 6518 2984
rect 8110 2932 8116 2984
rect 8168 2972 8174 2984
rect 9953 2975 10011 2981
rect 9953 2972 9965 2975
rect 8168 2944 9965 2972
rect 8168 2932 8174 2944
rect 9953 2941 9965 2944
rect 9999 2941 10011 2975
rect 9953 2935 10011 2941
rect 10502 2932 10508 2984
rect 10560 2972 10566 2984
rect 10597 2975 10655 2981
rect 10597 2972 10609 2975
rect 10560 2944 10609 2972
rect 10560 2932 10566 2944
rect 10597 2941 10609 2944
rect 10643 2941 10655 2975
rect 10597 2935 10655 2941
rect 11701 2975 11759 2981
rect 11701 2941 11713 2975
rect 11747 2972 11759 2975
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11747 2944 11897 2972
rect 11747 2941 11759 2944
rect 11701 2935 11759 2941
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11885 2935 11943 2941
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2972 12219 2975
rect 12618 2972 12624 2984
rect 12207 2944 12624 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12618 2932 12624 2944
rect 12676 2932 12682 2984
rect 13464 2972 13492 3012
rect 14777 3009 14789 3012
rect 14823 3009 14835 3043
rect 14777 3003 14835 3009
rect 14918 3000 14924 3052
rect 14976 3000 14982 3052
rect 15212 3049 15240 3148
rect 15838 3136 15844 3148
rect 15896 3136 15902 3188
rect 15197 3043 15255 3049
rect 15197 3009 15209 3043
rect 15243 3009 15255 3043
rect 15197 3003 15255 3009
rect 13280 2944 13492 2972
rect 8938 2904 8944 2916
rect 6380 2876 6592 2904
rect 4614 2836 4620 2848
rect 4080 2808 4620 2836
rect 4614 2796 4620 2808
rect 4672 2796 4678 2848
rect 6564 2836 6592 2876
rect 7760 2876 8944 2904
rect 7760 2836 7788 2876
rect 8938 2864 8944 2876
rect 8996 2864 9002 2916
rect 11054 2864 11060 2916
rect 11112 2864 11118 2916
rect 6564 2808 7788 2836
rect 8481 2839 8539 2845
rect 8481 2805 8493 2839
rect 8527 2836 8539 2839
rect 9214 2836 9220 2848
rect 8527 2808 9220 2836
rect 8527 2805 8539 2808
rect 8481 2799 8539 2805
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 10410 2796 10416 2848
rect 10468 2796 10474 2848
rect 11974 2796 11980 2848
rect 12032 2836 12038 2848
rect 13280 2836 13308 2944
rect 13538 2932 13544 2984
rect 13596 2972 13602 2984
rect 14369 2975 14427 2981
rect 14369 2972 14381 2975
rect 13596 2944 14381 2972
rect 13596 2932 13602 2944
rect 14369 2941 14381 2944
rect 14415 2941 14427 2975
rect 14369 2935 14427 2941
rect 13354 2864 13360 2916
rect 13412 2904 13418 2916
rect 14645 2907 14703 2913
rect 14645 2904 14657 2907
rect 13412 2876 14657 2904
rect 13412 2864 13418 2876
rect 14645 2873 14657 2876
rect 14691 2873 14703 2907
rect 14645 2867 14703 2873
rect 13633 2839 13691 2845
rect 13633 2836 13645 2839
rect 12032 2808 13645 2836
rect 12032 2796 12038 2808
rect 13633 2805 13645 2808
rect 13679 2805 13691 2839
rect 13633 2799 13691 2805
rect 13814 2796 13820 2848
rect 13872 2796 13878 2848
rect 15654 2796 15660 2848
rect 15712 2836 15718 2848
rect 22186 2836 22192 2848
rect 15712 2808 22192 2836
rect 15712 2796 15718 2808
rect 22186 2796 22192 2808
rect 22244 2796 22250 2848
rect 1104 2746 22816 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 20214 2746
rect 20266 2694 20278 2746
rect 20330 2694 20342 2746
rect 20394 2694 20406 2746
rect 20458 2694 20470 2746
rect 20522 2694 22816 2746
rect 1104 2672 22816 2694
rect 4522 2592 4528 2644
rect 4580 2632 4586 2644
rect 4706 2632 4712 2644
rect 4580 2604 4712 2632
rect 4580 2592 4586 2604
rect 4706 2592 4712 2604
rect 4764 2632 4770 2644
rect 5718 2632 5724 2644
rect 4764 2604 5724 2632
rect 4764 2592 4770 2604
rect 5718 2592 5724 2604
rect 5776 2592 5782 2644
rect 7180 2635 7238 2641
rect 7180 2601 7192 2635
rect 7226 2632 7238 2635
rect 9585 2635 9643 2641
rect 7226 2604 8800 2632
rect 7226 2601 7238 2604
rect 7180 2595 7238 2601
rect 3326 2524 3332 2576
rect 3384 2564 3390 2576
rect 8772 2564 8800 2604
rect 9585 2601 9597 2635
rect 9631 2632 9643 2635
rect 10134 2632 10140 2644
rect 9631 2604 10140 2632
rect 9631 2601 9643 2604
rect 9585 2595 9643 2601
rect 10134 2592 10140 2604
rect 10192 2592 10198 2644
rect 12342 2632 12348 2644
rect 10612 2604 12348 2632
rect 3384 2536 4016 2564
rect 8772 2536 9352 2564
rect 3384 2524 3390 2536
rect 1765 2499 1823 2505
rect 1765 2465 1777 2499
rect 1811 2496 1823 2499
rect 3510 2496 3516 2508
rect 1811 2468 3516 2496
rect 1811 2465 1823 2468
rect 1765 2459 1823 2465
rect 3510 2456 3516 2468
rect 3568 2456 3574 2508
rect 3602 2456 3608 2508
rect 3660 2496 3666 2508
rect 3881 2499 3939 2505
rect 3881 2496 3893 2499
rect 3660 2468 3893 2496
rect 3660 2456 3666 2468
rect 3881 2465 3893 2468
rect 3927 2465 3939 2499
rect 3988 2496 4016 2536
rect 6917 2499 6975 2505
rect 3988 2468 6224 2496
rect 3881 2459 3939 2465
rect 1486 2388 1492 2440
rect 1544 2388 1550 2440
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 5905 2431 5963 2437
rect 5905 2428 5917 2431
rect 5776 2400 5917 2428
rect 5776 2388 5782 2400
rect 5905 2397 5917 2400
rect 5951 2397 5963 2431
rect 5905 2391 5963 2397
rect 2038 2320 2044 2372
rect 2096 2320 2102 2372
rect 2774 2320 2780 2372
rect 2832 2320 2838 2372
rect 4157 2363 4215 2369
rect 4157 2329 4169 2363
rect 4203 2329 4215 2363
rect 4157 2323 4215 2329
rect 1581 2295 1639 2301
rect 1581 2261 1593 2295
rect 1627 2292 1639 2295
rect 2130 2292 2136 2304
rect 1627 2264 2136 2292
rect 1627 2261 1639 2264
rect 1581 2255 1639 2261
rect 2130 2252 2136 2264
rect 2188 2252 2194 2304
rect 3513 2295 3571 2301
rect 3513 2261 3525 2295
rect 3559 2292 3571 2295
rect 4172 2292 4200 2323
rect 4614 2320 4620 2372
rect 4672 2320 4678 2372
rect 3559 2264 4200 2292
rect 3559 2261 3571 2264
rect 3513 2255 3571 2261
rect 5534 2252 5540 2304
rect 5592 2292 5598 2304
rect 5629 2295 5687 2301
rect 5629 2292 5641 2295
rect 5592 2264 5641 2292
rect 5592 2252 5598 2264
rect 5629 2261 5641 2264
rect 5675 2292 5687 2295
rect 6086 2292 6092 2304
rect 5675 2264 6092 2292
rect 5675 2261 5687 2264
rect 5629 2255 5687 2261
rect 6086 2252 6092 2264
rect 6144 2252 6150 2304
rect 6196 2292 6224 2468
rect 6917 2465 6929 2499
rect 6963 2496 6975 2499
rect 8570 2496 8576 2508
rect 6963 2468 8576 2496
rect 6963 2465 6975 2468
rect 6917 2459 6975 2465
rect 8570 2456 8576 2468
rect 8628 2496 8634 2508
rect 9324 2496 9352 2536
rect 9766 2524 9772 2576
rect 9824 2564 9830 2576
rect 10042 2564 10048 2576
rect 9824 2536 10048 2564
rect 9824 2524 9830 2536
rect 10042 2524 10048 2536
rect 10100 2524 10106 2576
rect 10229 2567 10287 2573
rect 10229 2533 10241 2567
rect 10275 2533 10287 2567
rect 10229 2527 10287 2533
rect 10244 2496 10272 2527
rect 8628 2468 9260 2496
rect 9324 2468 10272 2496
rect 8628 2456 8634 2468
rect 8294 2388 8300 2440
rect 8352 2388 8358 2440
rect 9030 2388 9036 2440
rect 9088 2388 9094 2440
rect 9232 2437 9260 2468
rect 9217 2431 9275 2437
rect 9217 2397 9229 2431
rect 9263 2397 9275 2431
rect 9217 2391 9275 2397
rect 9398 2388 9404 2440
rect 9456 2437 9462 2440
rect 9456 2428 9464 2437
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9456 2400 9781 2428
rect 9456 2391 9464 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 10318 2428 10324 2440
rect 9769 2391 9827 2397
rect 9876 2400 10324 2428
rect 9456 2388 9462 2391
rect 6733 2363 6791 2369
rect 6733 2329 6745 2363
rect 6779 2360 6791 2363
rect 6822 2360 6828 2372
rect 6779 2332 6828 2360
rect 6779 2329 6791 2332
rect 6733 2323 6791 2329
rect 6822 2320 6828 2332
rect 6880 2320 6886 2372
rect 8496 2332 8800 2360
rect 8496 2292 8524 2332
rect 6196 2264 8524 2292
rect 8662 2252 8668 2304
rect 8720 2252 8726 2304
rect 8772 2292 8800 2332
rect 8938 2320 8944 2372
rect 8996 2360 9002 2372
rect 9309 2363 9367 2369
rect 9309 2360 9321 2363
rect 8996 2332 9321 2360
rect 8996 2320 9002 2332
rect 9309 2329 9321 2332
rect 9355 2329 9367 2363
rect 9876 2360 9904 2400
rect 10318 2388 10324 2400
rect 10376 2388 10382 2440
rect 10612 2437 10640 2604
rect 12342 2592 12348 2604
rect 12400 2592 12406 2644
rect 12437 2635 12495 2641
rect 12437 2601 12449 2635
rect 12483 2632 12495 2635
rect 12618 2632 12624 2644
rect 12483 2604 12624 2632
rect 12483 2601 12495 2604
rect 12437 2595 12495 2601
rect 12618 2592 12624 2604
rect 12676 2592 12682 2644
rect 12710 2592 12716 2644
rect 12768 2632 12774 2644
rect 13633 2635 13691 2641
rect 13633 2632 13645 2635
rect 12768 2604 13645 2632
rect 12768 2592 12774 2604
rect 13633 2601 13645 2604
rect 13679 2632 13691 2635
rect 13906 2632 13912 2644
rect 13679 2604 13912 2632
rect 13679 2601 13691 2604
rect 13633 2595 13691 2601
rect 13906 2592 13912 2604
rect 13964 2592 13970 2644
rect 13998 2592 14004 2644
rect 14056 2632 14062 2644
rect 14056 2604 18920 2632
rect 14056 2592 14062 2604
rect 11974 2524 11980 2576
rect 12032 2564 12038 2576
rect 14182 2564 14188 2576
rect 12032 2536 14188 2564
rect 12032 2524 12038 2536
rect 14182 2524 14188 2536
rect 14240 2524 14246 2576
rect 10965 2499 11023 2505
rect 10965 2465 10977 2499
rect 11011 2496 11023 2499
rect 11054 2496 11060 2508
rect 11011 2468 11060 2496
rect 11011 2465 11023 2468
rect 10965 2459 11023 2465
rect 11054 2456 11060 2468
rect 11112 2456 11118 2508
rect 11606 2456 11612 2508
rect 11664 2496 11670 2508
rect 13722 2496 13728 2508
rect 11664 2468 13728 2496
rect 11664 2456 11670 2468
rect 13722 2456 13728 2468
rect 13780 2456 13786 2508
rect 13906 2456 13912 2508
rect 13964 2496 13970 2508
rect 14553 2499 14611 2505
rect 14553 2496 14565 2499
rect 13964 2468 14565 2496
rect 13964 2456 13970 2468
rect 14553 2465 14565 2468
rect 14599 2465 14611 2499
rect 18892 2496 18920 2604
rect 18892 2468 21128 2496
rect 14553 2459 14611 2465
rect 10597 2431 10655 2437
rect 10597 2397 10609 2431
rect 10643 2397 10655 2431
rect 10597 2391 10655 2397
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2397 10747 2431
rect 13357 2431 13415 2437
rect 13357 2428 13369 2431
rect 12098 2400 13369 2428
rect 10689 2391 10747 2397
rect 13357 2397 13369 2400
rect 13403 2397 13415 2431
rect 13357 2391 13415 2397
rect 10704 2360 10732 2391
rect 13814 2388 13820 2440
rect 13872 2388 13878 2440
rect 14090 2388 14096 2440
rect 14148 2388 14154 2440
rect 21100 2437 21128 2468
rect 21085 2431 21143 2437
rect 21085 2397 21097 2431
rect 21131 2397 21143 2431
rect 21085 2391 21143 2397
rect 9309 2323 9367 2329
rect 9416 2332 9904 2360
rect 10336 2332 10732 2360
rect 9416 2292 9444 2332
rect 8772 2264 9444 2292
rect 9490 2252 9496 2304
rect 9548 2292 9554 2304
rect 10336 2292 10364 2332
rect 9548 2264 10364 2292
rect 10413 2295 10471 2301
rect 9548 2252 9554 2264
rect 10413 2261 10425 2295
rect 10459 2292 10471 2295
rect 10594 2292 10600 2304
rect 10459 2264 10600 2292
rect 10459 2261 10471 2264
rect 10413 2255 10471 2261
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 10704 2292 10732 2332
rect 10962 2320 10968 2372
rect 11020 2360 11026 2372
rect 11020 2332 11454 2360
rect 11020 2320 11026 2332
rect 12250 2320 12256 2372
rect 12308 2360 12314 2372
rect 12621 2363 12679 2369
rect 12621 2360 12633 2363
rect 12308 2332 12633 2360
rect 12308 2320 12314 2332
rect 12621 2329 12633 2332
rect 12667 2329 12679 2363
rect 22094 2360 22100 2372
rect 12621 2323 12679 2329
rect 13648 2332 22100 2360
rect 11054 2292 11060 2304
rect 10704 2264 11060 2292
rect 11054 2252 11060 2264
rect 11112 2252 11118 2304
rect 11882 2252 11888 2304
rect 11940 2292 11946 2304
rect 13648 2292 13676 2332
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 22281 2363 22339 2369
rect 22281 2329 22293 2363
rect 22327 2360 22339 2363
rect 23014 2360 23020 2372
rect 22327 2332 23020 2360
rect 22327 2329 22339 2332
rect 22281 2323 22339 2329
rect 23014 2320 23020 2332
rect 23072 2320 23078 2372
rect 11940 2264 13676 2292
rect 11940 2252 11946 2264
rect 13722 2252 13728 2304
rect 13780 2292 13786 2304
rect 15010 2292 15016 2304
rect 13780 2264 15016 2292
rect 13780 2252 13786 2264
rect 15010 2252 15016 2264
rect 15068 2252 15074 2304
rect 1104 2202 22816 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 22816 2202
rect 1104 2128 22816 2150
rect 1581 2091 1639 2097
rect 1581 2057 1593 2091
rect 1627 2088 1639 2091
rect 2038 2088 2044 2100
rect 1627 2060 2044 2088
rect 1627 2057 1639 2060
rect 1581 2051 1639 2057
rect 2038 2048 2044 2060
rect 2096 2048 2102 2100
rect 3418 2088 3424 2100
rect 2746 2060 3424 2088
rect 2746 2020 2774 2060
rect 3418 2048 3424 2060
rect 3476 2048 3482 2100
rect 3881 2091 3939 2097
rect 3881 2057 3893 2091
rect 3927 2088 3939 2091
rect 3970 2088 3976 2100
rect 3927 2060 3976 2088
rect 3927 2057 3939 2060
rect 3881 2051 3939 2057
rect 3970 2048 3976 2060
rect 4028 2048 4034 2100
rect 4157 2091 4215 2097
rect 4157 2057 4169 2091
rect 4203 2088 4215 2091
rect 6454 2088 6460 2100
rect 4203 2060 6460 2088
rect 4203 2057 4215 2060
rect 4157 2051 4215 2057
rect 6454 2048 6460 2060
rect 6512 2048 6518 2100
rect 6638 2048 6644 2100
rect 6696 2088 6702 2100
rect 9309 2091 9367 2097
rect 6696 2060 9168 2088
rect 6696 2048 6702 2060
rect 2056 1992 2774 2020
rect 2056 1961 2084 1992
rect 2866 1980 2872 2032
rect 2924 1980 2930 2032
rect 4614 2020 4620 2032
rect 3988 1992 4620 2020
rect 3988 1964 4016 1992
rect 4614 1980 4620 1992
rect 4672 2020 4678 2032
rect 4672 1992 5106 2020
rect 4672 1980 4678 1992
rect 6546 1980 6552 2032
rect 6604 1980 6610 2032
rect 8294 1980 8300 2032
rect 8352 1980 8358 2032
rect 9140 2020 9168 2060
rect 9309 2057 9321 2091
rect 9355 2088 9367 2091
rect 9398 2088 9404 2100
rect 9355 2060 9404 2088
rect 9355 2057 9367 2060
rect 9309 2051 9367 2057
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 9508 2060 11100 2088
rect 9508 2020 9536 2060
rect 9140 1992 9536 2020
rect 11072 2020 11100 2060
rect 11514 2048 11520 2100
rect 11572 2088 11578 2100
rect 14918 2088 14924 2100
rect 11572 2060 14924 2088
rect 11572 2048 11578 2060
rect 11606 2020 11612 2032
rect 11072 1992 11612 2020
rect 11606 1980 11612 1992
rect 11664 1980 11670 2032
rect 11793 2023 11851 2029
rect 11793 1989 11805 2023
rect 11839 2020 11851 2023
rect 11882 2020 11888 2032
rect 11839 1992 11888 2020
rect 11839 1989 11851 1992
rect 11793 1983 11851 1989
rect 11882 1980 11888 1992
rect 11940 1980 11946 2032
rect 11974 1980 11980 2032
rect 12032 1980 12038 2032
rect 2041 1955 2099 1961
rect 2041 1921 2053 1955
rect 2087 1921 2099 1955
rect 2041 1915 2099 1921
rect 2130 1912 2136 1964
rect 2188 1912 2194 1964
rect 3970 1912 3976 1964
rect 4028 1912 4034 1964
rect 4062 1912 4068 1964
rect 4120 1912 4126 1964
rect 5902 1912 5908 1964
rect 5960 1952 5966 1964
rect 6365 1955 6423 1961
rect 6365 1952 6377 1955
rect 5960 1924 6377 1952
rect 5960 1912 5966 1924
rect 6365 1921 6377 1924
rect 6411 1921 6423 1955
rect 6365 1915 6423 1921
rect 6641 1955 6699 1961
rect 6641 1921 6653 1955
rect 6687 1921 6699 1955
rect 6641 1915 6699 1921
rect 2406 1844 2412 1896
rect 2464 1844 2470 1896
rect 2774 1844 2780 1896
rect 2832 1884 2838 1896
rect 4080 1884 4108 1912
rect 2832 1856 4108 1884
rect 2832 1844 2838 1856
rect 1762 1776 1768 1828
rect 1820 1776 1826 1828
rect 4080 1748 4108 1856
rect 4154 1844 4160 1896
rect 4212 1884 4218 1896
rect 4341 1887 4399 1893
rect 4341 1884 4353 1887
rect 4212 1856 4353 1884
rect 4212 1844 4218 1856
rect 4341 1853 4353 1856
rect 4387 1853 4399 1887
rect 4341 1847 4399 1853
rect 4614 1844 4620 1896
rect 4672 1844 4678 1896
rect 5994 1844 6000 1896
rect 6052 1884 6058 1896
rect 6089 1887 6147 1893
rect 6089 1884 6101 1887
rect 6052 1856 6101 1884
rect 6052 1844 6058 1856
rect 6089 1853 6101 1856
rect 6135 1853 6147 1887
rect 6089 1847 6147 1853
rect 6656 1748 6684 1915
rect 6730 1912 6736 1964
rect 6788 1961 6794 1964
rect 6788 1915 6796 1961
rect 7285 1955 7343 1961
rect 7285 1921 7297 1955
rect 7331 1921 7343 1955
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 10902 1924 11529 1952
rect 7285 1915 7343 1921
rect 11517 1921 11529 1924
rect 11563 1952 11575 1955
rect 12618 1952 12624 1964
rect 11563 1924 12624 1952
rect 11563 1921 11575 1924
rect 11517 1915 11575 1921
rect 6788 1912 6794 1915
rect 7300 1884 7328 1915
rect 12618 1912 12624 1924
rect 12676 1912 12682 1964
rect 13924 1961 13952 2060
rect 14918 2048 14924 2060
rect 14976 2048 14982 2100
rect 15010 2048 15016 2100
rect 15068 2088 15074 2100
rect 15068 2060 18644 2088
rect 15068 2048 15074 2060
rect 13909 1955 13967 1961
rect 13909 1921 13921 1955
rect 13955 1921 13967 1955
rect 13909 1915 13967 1921
rect 14182 1912 14188 1964
rect 14240 1952 14246 1964
rect 14921 1955 14979 1961
rect 14921 1952 14933 1955
rect 14240 1924 14933 1952
rect 14240 1912 14246 1924
rect 14921 1921 14933 1924
rect 14967 1921 14979 1955
rect 14921 1915 14979 1921
rect 15010 1912 15016 1964
rect 15068 1952 15074 1964
rect 18616 1961 18644 2060
rect 16761 1955 16819 1961
rect 16761 1952 16773 1955
rect 15068 1924 16773 1952
rect 15068 1912 15074 1924
rect 16761 1921 16773 1924
rect 16807 1921 16819 1955
rect 16761 1915 16819 1921
rect 18601 1955 18659 1961
rect 18601 1921 18613 1955
rect 18647 1921 18659 1955
rect 18601 1915 18659 1921
rect 20254 1912 20260 1964
rect 20312 1912 20318 1964
rect 22097 1955 22155 1961
rect 22097 1921 22109 1955
rect 22143 1952 22155 1955
rect 22186 1952 22192 1964
rect 22143 1924 22192 1952
rect 22143 1921 22155 1924
rect 22097 1915 22155 1921
rect 22186 1912 22192 1924
rect 22244 1912 22250 1964
rect 6748 1856 7328 1884
rect 7377 1887 7435 1893
rect 6748 1828 6776 1856
rect 7377 1853 7389 1887
rect 7423 1884 7435 1887
rect 7561 1887 7619 1893
rect 7561 1884 7573 1887
rect 7423 1856 7573 1884
rect 7423 1853 7435 1856
rect 7377 1847 7435 1853
rect 7561 1853 7573 1856
rect 7607 1853 7619 1887
rect 7561 1847 7619 1853
rect 7834 1844 7840 1896
rect 7892 1844 7898 1896
rect 9490 1844 9496 1896
rect 9548 1844 9554 1896
rect 9769 1887 9827 1893
rect 9769 1853 9781 1887
rect 9815 1884 9827 1887
rect 10502 1884 10508 1896
rect 9815 1856 10508 1884
rect 9815 1853 9827 1856
rect 9769 1847 9827 1853
rect 10502 1844 10508 1856
rect 10560 1844 10566 1896
rect 10778 1844 10784 1896
rect 10836 1884 10842 1896
rect 12066 1884 12072 1896
rect 10836 1856 12072 1884
rect 10836 1844 10842 1856
rect 12066 1844 12072 1856
rect 12124 1844 12130 1896
rect 12161 1887 12219 1893
rect 12161 1853 12173 1887
rect 12207 1884 12219 1887
rect 13538 1884 13544 1896
rect 12207 1856 13544 1884
rect 12207 1853 12219 1856
rect 12161 1847 12219 1853
rect 13538 1844 13544 1856
rect 13596 1844 13602 1896
rect 13633 1887 13691 1893
rect 13633 1853 13645 1887
rect 13679 1884 13691 1887
rect 14001 1887 14059 1893
rect 14001 1884 14013 1887
rect 13679 1856 14013 1884
rect 13679 1853 13691 1856
rect 13633 1847 13691 1853
rect 14001 1853 14013 1856
rect 14047 1853 14059 1887
rect 14001 1847 14059 1853
rect 14550 1844 14556 1896
rect 14608 1844 14614 1896
rect 15654 1844 15660 1896
rect 15712 1844 15718 1896
rect 17494 1844 17500 1896
rect 17552 1844 17558 1896
rect 19334 1844 19340 1896
rect 19392 1844 19398 1896
rect 21174 1844 21180 1896
rect 21232 1844 21238 1896
rect 6730 1776 6736 1828
rect 6788 1776 6794 1828
rect 6914 1776 6920 1828
rect 6972 1776 6978 1828
rect 9508 1748 9536 1844
rect 11241 1819 11299 1825
rect 11241 1785 11253 1819
rect 11287 1816 11299 1819
rect 11287 1788 12664 1816
rect 11287 1785 11299 1788
rect 11241 1779 11299 1785
rect 4080 1720 9536 1748
rect 10134 1708 10140 1760
rect 10192 1748 10198 1760
rect 11793 1751 11851 1757
rect 11793 1748 11805 1751
rect 10192 1720 11805 1748
rect 10192 1708 10198 1720
rect 11793 1717 11805 1720
rect 11839 1717 11851 1751
rect 12636 1748 12664 1788
rect 14642 1748 14648 1760
rect 12636 1720 14648 1748
rect 11793 1711 11851 1717
rect 14642 1708 14648 1720
rect 14700 1708 14706 1760
rect 1104 1658 22816 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 20214 1658
rect 20266 1606 20278 1658
rect 20330 1606 20342 1658
rect 20394 1606 20406 1658
rect 20458 1606 20470 1658
rect 20522 1606 22816 1658
rect 1104 1584 22816 1606
rect 1489 1547 1547 1553
rect 1489 1513 1501 1547
rect 1535 1544 1547 1547
rect 2406 1544 2412 1556
rect 1535 1516 2412 1544
rect 1535 1513 1547 1516
rect 1489 1507 1547 1513
rect 2406 1504 2412 1516
rect 2464 1504 2470 1556
rect 2866 1504 2872 1556
rect 2924 1544 2930 1556
rect 3881 1547 3939 1553
rect 2924 1516 3832 1544
rect 2924 1504 2930 1516
rect 3804 1476 3832 1516
rect 3881 1513 3893 1547
rect 3927 1544 3939 1547
rect 4614 1544 4620 1556
rect 3927 1516 4620 1544
rect 3927 1513 3939 1516
rect 3881 1507 3939 1513
rect 4614 1504 4620 1516
rect 4672 1504 4678 1556
rect 5371 1547 5429 1553
rect 5371 1513 5383 1547
rect 5417 1544 5429 1547
rect 5626 1544 5632 1556
rect 5417 1516 5632 1544
rect 5417 1513 5429 1516
rect 5371 1507 5429 1513
rect 5626 1504 5632 1516
rect 5684 1504 5690 1556
rect 6917 1547 6975 1553
rect 6917 1513 6929 1547
rect 6963 1544 6975 1547
rect 7834 1544 7840 1556
rect 6963 1516 7840 1544
rect 6963 1513 6975 1516
rect 6917 1507 6975 1513
rect 7834 1504 7840 1516
rect 7892 1504 7898 1556
rect 8294 1504 8300 1556
rect 8352 1544 8358 1556
rect 8352 1516 8616 1544
rect 8352 1504 8358 1516
rect 3970 1476 3976 1488
rect 3804 1448 3976 1476
rect 3970 1436 3976 1448
rect 4028 1436 4034 1488
rect 8588 1476 8616 1516
rect 8662 1504 8668 1556
rect 8720 1544 8726 1556
rect 11069 1547 11127 1553
rect 11069 1544 11081 1547
rect 8720 1516 11081 1544
rect 8720 1504 8726 1516
rect 11069 1513 11081 1516
rect 11115 1513 11127 1547
rect 11069 1507 11127 1513
rect 11238 1504 11244 1556
rect 11296 1544 11302 1556
rect 15010 1544 15016 1556
rect 11296 1516 15016 1544
rect 11296 1504 11302 1516
rect 15010 1504 15016 1516
rect 15068 1504 15074 1556
rect 9858 1476 9864 1488
rect 8588 1448 9864 1476
rect 9858 1436 9864 1448
rect 9916 1436 9922 1488
rect 2961 1411 3019 1417
rect 2961 1377 2973 1411
rect 3007 1408 3019 1411
rect 6362 1408 6368 1420
rect 3007 1380 3464 1408
rect 3007 1377 3019 1380
rect 2961 1371 3019 1377
rect 934 1300 940 1352
rect 992 1340 998 1352
rect 1486 1340 1492 1352
rect 992 1312 1492 1340
rect 992 1300 998 1312
rect 1486 1300 1492 1312
rect 1544 1300 1550 1352
rect 3237 1343 3295 1349
rect 3237 1309 3249 1343
rect 3283 1309 3295 1343
rect 3237 1303 3295 1309
rect 1504 1204 1532 1300
rect 2866 1272 2872 1284
rect 2530 1244 2872 1272
rect 2866 1232 2872 1244
rect 2924 1232 2930 1284
rect 3252 1204 3280 1303
rect 1504 1176 3280 1204
rect 3436 1204 3464 1380
rect 3804 1380 6368 1408
rect 3804 1352 3832 1380
rect 3605 1343 3663 1349
rect 3605 1309 3617 1343
rect 3651 1340 3663 1343
rect 3786 1340 3792 1352
rect 3651 1312 3792 1340
rect 3651 1309 3663 1312
rect 3605 1303 3663 1309
rect 3786 1300 3792 1312
rect 3844 1300 3850 1352
rect 3970 1300 3976 1352
rect 4028 1340 4034 1352
rect 5644 1349 5672 1380
rect 6362 1368 6368 1380
rect 6420 1408 6426 1420
rect 6730 1408 6736 1420
rect 6420 1380 6736 1408
rect 6420 1368 6426 1380
rect 6730 1368 6736 1380
rect 6788 1408 6794 1420
rect 8665 1411 8723 1417
rect 8665 1408 8677 1411
rect 6788 1380 8677 1408
rect 6788 1368 6794 1380
rect 8665 1377 8677 1380
rect 8711 1408 8723 1411
rect 8938 1408 8944 1420
rect 8711 1380 8944 1408
rect 8711 1377 8723 1380
rect 8665 1371 8723 1377
rect 8938 1368 8944 1380
rect 8996 1368 9002 1420
rect 9030 1368 9036 1420
rect 9088 1408 9094 1420
rect 9585 1411 9643 1417
rect 9585 1408 9597 1411
rect 9088 1380 9597 1408
rect 9088 1368 9094 1380
rect 5629 1343 5687 1349
rect 4028 1312 4278 1340
rect 4028 1300 4034 1312
rect 5629 1309 5641 1343
rect 5675 1309 5687 1343
rect 5629 1303 5687 1309
rect 5718 1300 5724 1352
rect 5776 1300 5782 1352
rect 5902 1300 5908 1352
rect 5960 1300 5966 1352
rect 5994 1300 6000 1352
rect 6052 1340 6058 1352
rect 6457 1343 6515 1349
rect 6457 1340 6469 1343
rect 6052 1312 6469 1340
rect 6052 1300 6058 1312
rect 6457 1309 6469 1312
rect 6503 1309 6515 1343
rect 6457 1303 6515 1309
rect 6638 1300 6644 1352
rect 6696 1300 6702 1352
rect 9324 1349 9352 1380
rect 9585 1377 9597 1380
rect 9631 1377 9643 1411
rect 9585 1371 9643 1377
rect 11054 1368 11060 1420
rect 11112 1408 11118 1420
rect 11514 1408 11520 1420
rect 11112 1380 11520 1408
rect 11112 1368 11118 1380
rect 11514 1368 11520 1380
rect 11572 1368 11578 1420
rect 11793 1411 11851 1417
rect 11793 1377 11805 1411
rect 11839 1408 11851 1411
rect 11839 1380 14136 1408
rect 11839 1377 11851 1380
rect 11793 1371 11851 1377
rect 14108 1349 14136 1380
rect 9217 1343 9275 1349
rect 9217 1309 9229 1343
rect 9263 1309 9275 1343
rect 9217 1303 9275 1309
rect 9309 1343 9367 1349
rect 9309 1309 9321 1343
rect 9355 1309 9367 1343
rect 9309 1303 9367 1309
rect 11333 1343 11391 1349
rect 11333 1309 11345 1343
rect 11379 1309 11391 1343
rect 11333 1303 11391 1309
rect 14093 1343 14151 1349
rect 14093 1309 14105 1343
rect 14139 1309 14151 1343
rect 14093 1303 14151 1309
rect 3513 1275 3571 1281
rect 3513 1241 3525 1275
rect 3559 1272 3571 1275
rect 4062 1272 4068 1284
rect 3559 1244 4068 1272
rect 3559 1241 3571 1244
rect 3513 1235 3571 1241
rect 4062 1232 4068 1244
rect 4120 1232 4126 1284
rect 6365 1275 6423 1281
rect 6365 1272 6377 1275
rect 5552 1244 6377 1272
rect 5552 1204 5580 1244
rect 6365 1241 6377 1244
rect 6411 1241 6423 1275
rect 8294 1272 8300 1284
rect 7958 1244 8300 1272
rect 6365 1235 6423 1241
rect 8294 1232 8300 1244
rect 8352 1232 8358 1284
rect 8389 1275 8447 1281
rect 8389 1241 8401 1275
rect 8435 1272 8447 1275
rect 9033 1275 9091 1281
rect 9033 1272 9045 1275
rect 8435 1244 9045 1272
rect 8435 1241 8447 1244
rect 8389 1235 8447 1241
rect 9033 1241 9045 1244
rect 9079 1241 9091 1275
rect 9232 1272 9260 1303
rect 9766 1272 9772 1284
rect 9232 1244 9772 1272
rect 9033 1235 9091 1241
rect 9766 1232 9772 1244
rect 9824 1232 9830 1284
rect 10962 1272 10968 1284
rect 10626 1244 10968 1272
rect 10962 1232 10968 1244
rect 11020 1232 11026 1284
rect 3436 1176 5580 1204
rect 5810 1164 5816 1216
rect 5868 1164 5874 1216
rect 10410 1164 10416 1216
rect 10468 1204 10474 1216
rect 11348 1204 11376 1303
rect 14642 1300 14648 1352
rect 14700 1300 14706 1352
rect 12526 1232 12532 1284
rect 12584 1232 12590 1284
rect 10468 1176 11376 1204
rect 13265 1207 13323 1213
rect 10468 1164 10474 1176
rect 13265 1173 13277 1207
rect 13311 1204 13323 1207
rect 14550 1204 14556 1216
rect 13311 1176 14556 1204
rect 13311 1173 13323 1176
rect 13265 1167 13323 1173
rect 14550 1164 14556 1176
rect 14608 1164 14614 1216
rect 1104 1114 22816 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 22816 1114
rect 1104 1040 22816 1062
rect 1762 960 1768 1012
rect 1820 1000 1826 1012
rect 5718 1000 5724 1012
rect 1820 972 5724 1000
rect 1820 960 1826 972
rect 5718 960 5724 972
rect 5776 960 5782 1012
<< via1 >>
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 20214 13574 20266 13626
rect 20278 13574 20330 13626
rect 20342 13574 20394 13626
rect 20406 13574 20458 13626
rect 20470 13574 20522 13626
rect 1492 13175 1544 13184
rect 1492 13141 1501 13175
rect 1501 13141 1535 13175
rect 1535 13141 1544 13175
rect 1492 13132 1544 13141
rect 2964 13243 3016 13252
rect 2964 13209 2973 13243
rect 2973 13209 3007 13243
rect 3007 13209 3016 13243
rect 2964 13200 3016 13209
rect 3700 13268 3752 13320
rect 3884 13200 3936 13252
rect 4160 13311 4212 13320
rect 4160 13277 4174 13311
rect 4174 13277 4208 13311
rect 4208 13277 4212 13311
rect 5540 13404 5592 13456
rect 10232 13447 10284 13456
rect 10232 13413 10241 13447
rect 10241 13413 10275 13447
rect 10275 13413 10284 13447
rect 10232 13404 10284 13413
rect 6184 13336 6236 13388
rect 4160 13268 4212 13277
rect 5540 13311 5592 13320
rect 5540 13277 5549 13311
rect 5549 13277 5583 13311
rect 5583 13277 5592 13311
rect 5540 13268 5592 13277
rect 3148 13132 3200 13184
rect 3332 13132 3384 13184
rect 3792 13132 3844 13184
rect 6092 13200 6144 13252
rect 6736 13268 6788 13320
rect 10232 13268 10284 13320
rect 11152 13311 11204 13320
rect 11152 13277 11161 13311
rect 11161 13277 11195 13311
rect 11195 13277 11204 13311
rect 11152 13268 11204 13277
rect 11704 13268 11756 13320
rect 7012 13200 7064 13252
rect 4344 13132 4396 13184
rect 5632 13132 5684 13184
rect 7564 13200 7616 13252
rect 10692 13200 10744 13252
rect 13268 13268 13320 13320
rect 14740 13311 14792 13320
rect 14740 13277 14749 13311
rect 14749 13277 14783 13311
rect 14783 13277 14792 13311
rect 14740 13268 14792 13277
rect 15476 13311 15528 13320
rect 15476 13277 15485 13311
rect 15485 13277 15519 13311
rect 15519 13277 15528 13311
rect 15476 13268 15528 13277
rect 16120 13268 16172 13320
rect 16580 13268 16632 13320
rect 17408 13311 17460 13320
rect 17408 13277 17417 13311
rect 17417 13277 17451 13311
rect 17451 13277 17460 13311
rect 17408 13268 17460 13277
rect 11980 13243 12032 13252
rect 11980 13209 11989 13243
rect 11989 13209 12023 13243
rect 12023 13209 12032 13243
rect 11980 13200 12032 13209
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9772 13132 9824 13184
rect 10508 13132 10560 13184
rect 11520 13132 11572 13184
rect 11704 13132 11756 13184
rect 20628 13200 20680 13252
rect 21824 13268 21876 13320
rect 21732 13200 21784 13252
rect 22284 13200 22336 13252
rect 14832 13132 14884 13184
rect 15568 13132 15620 13184
rect 16672 13132 16724 13184
rect 16764 13132 16816 13184
rect 18604 13132 18656 13184
rect 19800 13175 19852 13184
rect 19800 13141 19809 13175
rect 19809 13141 19843 13175
rect 19843 13141 19852 13175
rect 19800 13132 19852 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 16214 13030 16266 13082
rect 16278 13030 16330 13082
rect 16342 13030 16394 13082
rect 16406 13030 16458 13082
rect 16470 13030 16522 13082
rect 6092 12971 6144 12980
rect 6092 12937 6101 12971
rect 6101 12937 6135 12971
rect 6135 12937 6144 12971
rect 6092 12928 6144 12937
rect 1492 12860 1544 12912
rect 1768 12699 1820 12708
rect 1768 12665 1777 12699
rect 1777 12665 1811 12699
rect 1811 12665 1820 12699
rect 1768 12656 1820 12665
rect 2044 12588 2096 12640
rect 2228 12767 2280 12776
rect 2228 12733 2237 12767
rect 2237 12733 2271 12767
rect 2271 12733 2280 12767
rect 2228 12724 2280 12733
rect 3148 12724 3200 12776
rect 5080 12860 5132 12912
rect 5172 12860 5224 12912
rect 4344 12835 4396 12844
rect 4344 12801 4353 12835
rect 4353 12801 4387 12835
rect 4387 12801 4396 12835
rect 4344 12792 4396 12801
rect 6368 12792 6420 12844
rect 6736 12860 6788 12912
rect 6920 12792 6972 12844
rect 7196 12928 7248 12980
rect 9404 12928 9456 12980
rect 9680 12928 9732 12980
rect 9496 12860 9548 12912
rect 9772 12903 9824 12912
rect 9772 12869 9781 12903
rect 9781 12869 9815 12903
rect 9815 12869 9824 12903
rect 9772 12860 9824 12869
rect 13268 12971 13320 12980
rect 13268 12937 13277 12971
rect 13277 12937 13311 12971
rect 13311 12937 13320 12971
rect 13268 12928 13320 12937
rect 14740 12971 14792 12980
rect 14740 12937 14749 12971
rect 14749 12937 14783 12971
rect 14783 12937 14792 12971
rect 14740 12928 14792 12937
rect 15476 12971 15528 12980
rect 15476 12937 15485 12971
rect 15485 12937 15519 12971
rect 15519 12937 15528 12971
rect 15476 12928 15528 12937
rect 16120 12928 16172 12980
rect 13820 12860 13872 12912
rect 16672 12903 16724 12912
rect 16672 12869 16681 12903
rect 16681 12869 16715 12903
rect 16715 12869 16724 12903
rect 16672 12860 16724 12869
rect 17868 12903 17920 12912
rect 17868 12869 17877 12903
rect 17877 12869 17911 12903
rect 17911 12869 17920 12903
rect 17868 12860 17920 12869
rect 18604 12903 18656 12912
rect 18604 12869 18613 12903
rect 18613 12869 18647 12903
rect 18647 12869 18656 12903
rect 18604 12860 18656 12869
rect 18880 12903 18932 12912
rect 18880 12869 18889 12903
rect 18889 12869 18923 12903
rect 18923 12869 18932 12903
rect 18880 12860 18932 12869
rect 4620 12767 4672 12776
rect 4620 12733 4629 12767
rect 4629 12733 4663 12767
rect 4663 12733 4672 12767
rect 4620 12724 4672 12733
rect 6184 12724 6236 12776
rect 11520 12835 11572 12844
rect 11520 12801 11529 12835
rect 11529 12801 11563 12835
rect 11563 12801 11572 12835
rect 11520 12792 11572 12801
rect 13452 12835 13504 12844
rect 13452 12801 13461 12835
rect 13461 12801 13495 12835
rect 13495 12801 13504 12835
rect 13452 12792 13504 12801
rect 7472 12724 7524 12776
rect 11152 12724 11204 12776
rect 14832 12792 14884 12844
rect 15568 12792 15620 12844
rect 16028 12792 16080 12844
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 19984 12860 20036 12912
rect 22100 12860 22152 12912
rect 22652 12860 22704 12912
rect 20812 12724 20864 12776
rect 4160 12588 4212 12640
rect 7656 12588 7708 12640
rect 21824 12631 21876 12640
rect 21824 12597 21833 12631
rect 21833 12597 21867 12631
rect 21867 12597 21876 12631
rect 21824 12588 21876 12597
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 20214 12486 20266 12538
rect 20278 12486 20330 12538
rect 20342 12486 20394 12538
rect 20406 12486 20458 12538
rect 20470 12486 20522 12538
rect 2228 12384 2280 12436
rect 2412 12384 2464 12436
rect 2780 12248 2832 12300
rect 1676 12223 1728 12232
rect 1676 12189 1685 12223
rect 1685 12189 1719 12223
rect 1719 12189 1728 12223
rect 1676 12180 1728 12189
rect 3148 12180 3200 12232
rect 3884 12384 3936 12436
rect 4620 12384 4672 12436
rect 6736 12384 6788 12436
rect 10692 12384 10744 12436
rect 13452 12384 13504 12436
rect 16580 12427 16632 12436
rect 16580 12393 16589 12427
rect 16589 12393 16623 12427
rect 16623 12393 16632 12427
rect 16580 12384 16632 12393
rect 17408 12384 17460 12436
rect 5908 12248 5960 12300
rect 6184 12291 6236 12300
rect 6184 12257 6193 12291
rect 6193 12257 6227 12291
rect 6227 12257 6236 12291
rect 6184 12248 6236 12257
rect 2044 12155 2096 12164
rect 2044 12121 2053 12155
rect 2053 12121 2087 12155
rect 2087 12121 2096 12155
rect 2044 12112 2096 12121
rect 3792 12155 3844 12164
rect 3792 12121 3801 12155
rect 3801 12121 3835 12155
rect 3835 12121 3844 12155
rect 3792 12112 3844 12121
rect 3608 12044 3660 12096
rect 3976 12087 4028 12096
rect 3976 12053 3985 12087
rect 3985 12053 4019 12087
rect 4019 12053 4028 12087
rect 3976 12044 4028 12053
rect 6276 12223 6328 12232
rect 6276 12189 6285 12223
rect 6285 12189 6319 12223
rect 6319 12189 6328 12223
rect 6276 12180 6328 12189
rect 9772 12248 9824 12300
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 11888 12248 11940 12300
rect 15752 12248 15804 12300
rect 10876 12223 10928 12232
rect 10876 12189 10885 12223
rect 10885 12189 10919 12223
rect 10919 12189 10928 12223
rect 10876 12180 10928 12189
rect 13728 12223 13780 12232
rect 13728 12189 13737 12223
rect 13737 12189 13771 12223
rect 13771 12189 13780 12223
rect 13728 12180 13780 12189
rect 16764 12223 16816 12232
rect 16764 12189 16773 12223
rect 16773 12189 16807 12223
rect 16807 12189 16816 12223
rect 16764 12180 16816 12189
rect 18328 12223 18380 12232
rect 18328 12189 18337 12223
rect 18337 12189 18371 12223
rect 18371 12189 18380 12223
rect 18328 12180 18380 12189
rect 20076 12291 20128 12300
rect 20076 12257 20085 12291
rect 20085 12257 20119 12291
rect 20119 12257 20128 12291
rect 20076 12248 20128 12257
rect 20628 12248 20680 12300
rect 22284 12291 22336 12300
rect 22284 12257 22293 12291
rect 22293 12257 22327 12291
rect 22327 12257 22336 12291
rect 22284 12248 22336 12257
rect 19800 12180 19852 12232
rect 19984 12180 20036 12232
rect 5448 12112 5500 12164
rect 5632 12112 5684 12164
rect 6552 12155 6604 12164
rect 6552 12121 6561 12155
rect 6561 12121 6595 12155
rect 6595 12121 6604 12155
rect 6552 12112 6604 12121
rect 8116 12112 8168 12164
rect 6736 12044 6788 12096
rect 6828 12044 6880 12096
rect 9496 12112 9548 12164
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 12624 12112 12676 12164
rect 14372 12155 14424 12164
rect 14372 12121 14381 12155
rect 14381 12121 14415 12155
rect 14415 12121 14424 12155
rect 14372 12112 14424 12121
rect 14740 12044 14792 12096
rect 18880 12044 18932 12096
rect 22100 12112 22152 12164
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 16214 11942 16266 11994
rect 16278 11942 16330 11994
rect 16342 11942 16394 11994
rect 16406 11942 16458 11994
rect 16470 11942 16522 11994
rect 2964 11840 3016 11892
rect 1676 11747 1728 11756
rect 1676 11713 1685 11747
rect 1685 11713 1719 11747
rect 1719 11713 1728 11747
rect 1676 11704 1728 11713
rect 2780 11772 2832 11824
rect 3700 11840 3752 11892
rect 6276 11840 6328 11892
rect 3608 11815 3660 11824
rect 3608 11781 3617 11815
rect 3617 11781 3651 11815
rect 3651 11781 3660 11815
rect 3608 11772 3660 11781
rect 5172 11772 5224 11824
rect 5448 11772 5500 11824
rect 6828 11772 6880 11824
rect 8024 11772 8076 11824
rect 8208 11772 8260 11824
rect 10876 11840 10928 11892
rect 11244 11883 11296 11892
rect 11244 11849 11253 11883
rect 11253 11849 11287 11883
rect 11287 11849 11296 11883
rect 11244 11840 11296 11849
rect 14372 11840 14424 11892
rect 18328 11840 18380 11892
rect 19616 11840 19668 11892
rect 20812 11840 20864 11892
rect 10324 11772 10376 11824
rect 1860 11636 1912 11688
rect 2412 11636 2464 11688
rect 3332 11747 3384 11756
rect 3332 11713 3341 11747
rect 3341 11713 3375 11747
rect 3375 11713 3384 11747
rect 3332 11704 3384 11713
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 3976 11636 4028 11688
rect 5816 11704 5868 11756
rect 6276 11704 6328 11756
rect 6736 11747 6788 11756
rect 6736 11713 6745 11747
rect 6745 11713 6779 11747
rect 6779 11713 6788 11747
rect 6736 11704 6788 11713
rect 7012 11704 7064 11756
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 6368 11568 6420 11620
rect 6460 11611 6512 11620
rect 6460 11577 6469 11611
rect 6469 11577 6503 11611
rect 6503 11577 6512 11611
rect 6460 11568 6512 11577
rect 6920 11568 6972 11620
rect 7656 11747 7708 11756
rect 7656 11713 7665 11747
rect 7665 11713 7699 11747
rect 7699 11713 7708 11747
rect 7656 11704 7708 11713
rect 9588 11704 9640 11756
rect 8576 11636 8628 11688
rect 9404 11679 9456 11688
rect 9404 11645 9413 11679
rect 9413 11645 9447 11679
rect 9447 11645 9456 11679
rect 9404 11636 9456 11645
rect 7472 11611 7524 11620
rect 7472 11577 7481 11611
rect 7481 11577 7515 11611
rect 7515 11577 7524 11611
rect 7472 11568 7524 11577
rect 8024 11500 8076 11552
rect 9680 11500 9732 11552
rect 10508 11704 10560 11756
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 11060 11747 11112 11756
rect 11060 11713 11069 11747
rect 11069 11713 11103 11747
rect 11103 11713 11112 11747
rect 11060 11704 11112 11713
rect 12072 11772 12124 11824
rect 11612 11747 11664 11756
rect 11612 11713 11621 11747
rect 11621 11713 11655 11747
rect 11655 11713 11664 11747
rect 11612 11704 11664 11713
rect 13544 11704 13596 11756
rect 10784 11568 10836 11620
rect 10876 11568 10928 11620
rect 12716 11679 12768 11688
rect 12716 11645 12725 11679
rect 12725 11645 12759 11679
rect 12759 11645 12768 11679
rect 12716 11636 12768 11645
rect 13452 11636 13504 11688
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 16672 11747 16724 11756
rect 16672 11713 16681 11747
rect 16681 11713 16715 11747
rect 16715 11713 16724 11747
rect 16672 11704 16724 11713
rect 18880 11747 18932 11756
rect 18880 11713 18889 11747
rect 18889 11713 18923 11747
rect 18923 11713 18932 11747
rect 18880 11704 18932 11713
rect 21824 11704 21876 11756
rect 16028 11568 16080 11620
rect 11152 11500 11204 11552
rect 13360 11500 13412 11552
rect 15384 11543 15436 11552
rect 15384 11509 15393 11543
rect 15393 11509 15427 11543
rect 15427 11509 15436 11543
rect 15384 11500 15436 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 20214 11398 20266 11450
rect 20278 11398 20330 11450
rect 20342 11398 20394 11450
rect 20406 11398 20458 11450
rect 20470 11398 20522 11450
rect 2780 11296 2832 11348
rect 3884 11296 3936 11348
rect 5448 11296 5500 11348
rect 6552 11296 6604 11348
rect 8668 11296 8720 11348
rect 12716 11296 12768 11348
rect 2688 11160 2740 11212
rect 3884 11203 3936 11212
rect 3884 11169 3893 11203
rect 3893 11169 3927 11203
rect 3927 11169 3936 11203
rect 3884 11160 3936 11169
rect 3976 11160 4028 11212
rect 3608 11135 3660 11144
rect 3608 11101 3617 11135
rect 3617 11101 3651 11135
rect 3651 11101 3660 11135
rect 3608 11092 3660 11101
rect 3792 11092 3844 11144
rect 6460 11160 6512 11212
rect 2872 11024 2924 11076
rect 4528 11067 4580 11076
rect 4528 11033 4537 11067
rect 4537 11033 4571 11067
rect 4571 11033 4580 11067
rect 4528 11024 4580 11033
rect 6920 11203 6972 11212
rect 6920 11169 6929 11203
rect 6929 11169 6963 11203
rect 6963 11169 6972 11203
rect 6920 11160 6972 11169
rect 10876 11203 10928 11212
rect 10876 11169 10885 11203
rect 10885 11169 10919 11203
rect 10919 11169 10928 11203
rect 10876 11160 10928 11169
rect 11152 11203 11204 11212
rect 11152 11169 11161 11203
rect 11161 11169 11195 11203
rect 11195 11169 11204 11203
rect 11152 11160 11204 11169
rect 11244 11203 11296 11212
rect 11244 11169 11253 11203
rect 11253 11169 11287 11203
rect 11287 11169 11296 11203
rect 11244 11160 11296 11169
rect 12072 11160 12124 11212
rect 9404 11092 9456 11144
rect 12624 11092 12676 11144
rect 4896 10956 4948 11008
rect 5908 10956 5960 11008
rect 7564 10956 7616 11008
rect 8852 11024 8904 11076
rect 10968 11024 11020 11076
rect 8668 10999 8720 11008
rect 8668 10965 8677 10999
rect 8677 10965 8711 10999
rect 8711 10965 8720 10999
rect 8668 10956 8720 10965
rect 9036 10999 9088 11008
rect 9036 10965 9045 10999
rect 9045 10965 9079 10999
rect 9079 10965 9088 10999
rect 9036 10956 9088 10965
rect 9588 10956 9640 11008
rect 10600 10956 10652 11008
rect 11060 10956 11112 11008
rect 11336 10956 11388 11008
rect 13728 11339 13780 11348
rect 13728 11305 13737 11339
rect 13737 11305 13771 11339
rect 13771 11305 13780 11339
rect 13728 11296 13780 11305
rect 16672 11339 16724 11348
rect 16672 11305 16681 11339
rect 16681 11305 16715 11339
rect 16715 11305 16724 11339
rect 16672 11296 16724 11305
rect 13452 11135 13504 11144
rect 13452 11101 13461 11135
rect 13461 11101 13495 11135
rect 13495 11101 13504 11135
rect 13452 11092 13504 11101
rect 13544 11135 13596 11144
rect 13544 11101 13558 11135
rect 13558 11101 13592 11135
rect 13592 11101 13596 11135
rect 15384 11160 15436 11212
rect 13544 11092 13596 11101
rect 16028 11135 16080 11144
rect 16028 11101 16037 11135
rect 16037 11101 16071 11135
rect 16071 11101 16080 11135
rect 16028 11092 16080 11101
rect 13820 11024 13872 11076
rect 15752 11067 15804 11076
rect 15752 11033 15761 11067
rect 15761 11033 15795 11067
rect 15795 11033 15804 11067
rect 15752 11024 15804 11033
rect 15016 10956 15068 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 16214 10854 16266 10906
rect 16278 10854 16330 10906
rect 16342 10854 16394 10906
rect 16406 10854 16458 10906
rect 16470 10854 16522 10906
rect 1676 10752 1728 10804
rect 3792 10752 3844 10804
rect 5816 10752 5868 10804
rect 2872 10684 2924 10736
rect 4528 10684 4580 10736
rect 4896 10684 4948 10736
rect 1676 10659 1728 10668
rect 1676 10625 1685 10659
rect 1685 10625 1719 10659
rect 1719 10625 1728 10659
rect 1676 10616 1728 10625
rect 5908 10616 5960 10668
rect 9036 10752 9088 10804
rect 9680 10752 9732 10804
rect 8852 10684 8904 10736
rect 9956 10727 10008 10736
rect 9956 10693 9965 10727
rect 9965 10693 9999 10727
rect 9999 10693 10008 10727
rect 9956 10684 10008 10693
rect 9680 10616 9732 10668
rect 10508 10752 10560 10804
rect 11060 10752 11112 10804
rect 10324 10684 10376 10736
rect 1952 10591 2004 10600
rect 1952 10557 1961 10591
rect 1961 10557 1995 10591
rect 1995 10557 2004 10591
rect 1952 10548 2004 10557
rect 4160 10591 4212 10600
rect 4160 10557 4169 10591
rect 4169 10557 4203 10591
rect 4203 10557 4212 10591
rect 4160 10548 4212 10557
rect 5816 10548 5868 10600
rect 6460 10548 6512 10600
rect 8668 10548 8720 10600
rect 10600 10616 10652 10668
rect 10784 10659 10836 10668
rect 10784 10625 10793 10659
rect 10793 10625 10827 10659
rect 10827 10625 10836 10659
rect 10784 10616 10836 10625
rect 11060 10616 11112 10668
rect 11336 10616 11388 10668
rect 11704 10659 11756 10668
rect 11704 10625 11713 10659
rect 11713 10625 11747 10659
rect 11747 10625 11756 10659
rect 11704 10616 11756 10625
rect 11796 10659 11848 10668
rect 11796 10625 11805 10659
rect 11805 10625 11839 10659
rect 11839 10625 11848 10659
rect 11796 10616 11848 10625
rect 15752 10752 15804 10804
rect 13360 10727 13412 10736
rect 13360 10693 13369 10727
rect 13369 10693 13403 10727
rect 13403 10693 13412 10727
rect 13360 10684 13412 10693
rect 13820 10684 13872 10736
rect 15936 10684 15988 10736
rect 11980 10659 12032 10668
rect 11980 10625 11983 10659
rect 11983 10625 12032 10659
rect 11980 10616 12032 10625
rect 15292 10659 15344 10668
rect 15292 10625 15296 10659
rect 15296 10625 15330 10659
rect 15330 10625 15344 10659
rect 15292 10616 15344 10625
rect 13452 10548 13504 10600
rect 15660 10659 15712 10668
rect 15660 10625 15669 10659
rect 15669 10625 15703 10659
rect 15703 10625 15712 10659
rect 15660 10616 15712 10625
rect 15752 10591 15804 10600
rect 15752 10557 15761 10591
rect 15761 10557 15795 10591
rect 15795 10557 15804 10591
rect 15752 10548 15804 10557
rect 4896 10412 4948 10464
rect 6276 10412 6328 10464
rect 8116 10412 8168 10464
rect 11520 10412 11572 10464
rect 11888 10412 11940 10464
rect 12992 10412 13044 10464
rect 13912 10412 13964 10464
rect 16580 10480 16632 10532
rect 17960 10548 18012 10600
rect 15108 10455 15160 10464
rect 15108 10421 15117 10455
rect 15117 10421 15151 10455
rect 15151 10421 15160 10455
rect 15108 10412 15160 10421
rect 16488 10412 16540 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 20214 10310 20266 10362
rect 20278 10310 20330 10362
rect 20342 10310 20394 10362
rect 20406 10310 20458 10362
rect 20470 10310 20522 10362
rect 1952 10208 2004 10260
rect 2872 10208 2924 10260
rect 3608 10208 3660 10260
rect 4068 10208 4120 10260
rect 2504 10140 2556 10192
rect 3792 10140 3844 10192
rect 4804 10140 4856 10192
rect 2136 10047 2188 10056
rect 2136 10013 2145 10047
rect 2145 10013 2179 10047
rect 2179 10013 2188 10047
rect 2136 10004 2188 10013
rect 2504 10047 2556 10056
rect 2504 10013 2513 10047
rect 2513 10013 2547 10047
rect 2547 10013 2556 10047
rect 2504 10004 2556 10013
rect 3884 10072 3936 10124
rect 6000 10208 6052 10260
rect 6920 10208 6972 10260
rect 11336 10208 11388 10260
rect 11612 10208 11664 10260
rect 13452 10208 13504 10260
rect 8024 10140 8076 10192
rect 2872 10004 2924 10056
rect 3700 10004 3752 10056
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 4804 10047 4856 10056
rect 4804 10013 4813 10047
rect 4813 10013 4847 10047
rect 4847 10013 4856 10047
rect 4804 10004 4856 10013
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 5908 10072 5960 10124
rect 2044 9868 2096 9920
rect 4252 9936 4304 9988
rect 4620 9936 4672 9988
rect 7196 10004 7248 10056
rect 7656 10047 7708 10056
rect 7656 10013 7665 10047
rect 7665 10013 7699 10047
rect 7699 10013 7708 10047
rect 7656 10004 7708 10013
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 8116 10047 8168 10056
rect 8116 10013 8125 10047
rect 8125 10013 8159 10047
rect 8159 10013 8168 10047
rect 8116 10004 8168 10013
rect 8576 10140 8628 10192
rect 9772 10115 9824 10124
rect 9772 10081 9781 10115
rect 9781 10081 9815 10115
rect 9815 10081 9824 10115
rect 9772 10072 9824 10081
rect 5908 9936 5960 9988
rect 6276 9936 6328 9988
rect 6644 9868 6696 9920
rect 7104 9868 7156 9920
rect 8760 9936 8812 9988
rect 9496 9936 9548 9988
rect 10508 10047 10560 10056
rect 10508 10013 10517 10047
rect 10517 10013 10551 10047
rect 10551 10013 10560 10047
rect 10508 10004 10560 10013
rect 11520 10115 11572 10124
rect 11520 10081 11529 10115
rect 11529 10081 11563 10115
rect 11563 10081 11572 10115
rect 11520 10072 11572 10081
rect 10876 10047 10928 10056
rect 10876 10013 10890 10047
rect 10890 10013 10924 10047
rect 10924 10013 10928 10047
rect 10876 10004 10928 10013
rect 10232 9936 10284 9988
rect 10784 9979 10836 9988
rect 10784 9945 10793 9979
rect 10793 9945 10827 9979
rect 10827 9945 10836 9979
rect 10784 9936 10836 9945
rect 13084 9936 13136 9988
rect 13268 9936 13320 9988
rect 13544 9979 13596 9988
rect 13544 9945 13553 9979
rect 13553 9945 13587 9979
rect 13587 9945 13596 9979
rect 13544 9936 13596 9945
rect 15660 10208 15712 10260
rect 15752 10208 15804 10260
rect 17960 10251 18012 10260
rect 17960 10217 17969 10251
rect 17969 10217 18003 10251
rect 18003 10217 18012 10251
rect 17960 10208 18012 10217
rect 15108 10072 15160 10124
rect 16488 10115 16540 10124
rect 16488 10081 16497 10115
rect 16497 10081 16531 10115
rect 16531 10081 16540 10115
rect 16488 10072 16540 10081
rect 13912 10047 13964 10056
rect 13912 10013 13921 10047
rect 13921 10013 13955 10047
rect 13955 10013 13964 10047
rect 13912 10004 13964 10013
rect 13176 9868 13228 9920
rect 15936 10004 15988 10056
rect 14832 9936 14884 9988
rect 15016 9936 15068 9988
rect 16580 9936 16632 9988
rect 15476 9868 15528 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 16214 9766 16266 9818
rect 16278 9766 16330 9818
rect 16342 9766 16394 9818
rect 16406 9766 16458 9818
rect 16470 9766 16522 9818
rect 2504 9664 2556 9716
rect 6276 9664 6328 9716
rect 2044 9571 2096 9580
rect 2044 9537 2053 9571
rect 2053 9537 2087 9571
rect 2087 9537 2096 9571
rect 2044 9528 2096 9537
rect 3424 9528 3476 9580
rect 4252 9528 4304 9580
rect 6644 9596 6696 9648
rect 9404 9664 9456 9716
rect 8760 9639 8812 9648
rect 8760 9605 8769 9639
rect 8769 9605 8803 9639
rect 8803 9605 8812 9639
rect 8760 9596 8812 9605
rect 13084 9664 13136 9716
rect 13176 9664 13228 9716
rect 15292 9664 15344 9716
rect 10232 9596 10284 9648
rect 12072 9596 12124 9648
rect 4804 9528 4856 9580
rect 5448 9528 5500 9580
rect 5816 9571 5868 9580
rect 5816 9537 5825 9571
rect 5825 9537 5859 9571
rect 5859 9537 5868 9571
rect 5816 9528 5868 9537
rect 6000 9571 6052 9580
rect 6000 9537 6003 9571
rect 6003 9537 6052 9571
rect 6000 9528 6052 9537
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 10048 9528 10100 9580
rect 10600 9528 10652 9580
rect 10784 9528 10836 9580
rect 2320 9503 2372 9512
rect 2320 9469 2329 9503
rect 2329 9469 2363 9503
rect 2363 9469 2372 9503
rect 2320 9460 2372 9469
rect 1308 9392 1360 9444
rect 3700 9392 3752 9444
rect 7196 9460 7248 9512
rect 7656 9460 7708 9512
rect 9772 9460 9824 9512
rect 10232 9503 10284 9512
rect 10232 9469 10241 9503
rect 10241 9469 10275 9503
rect 10275 9469 10284 9503
rect 10232 9460 10284 9469
rect 10968 9460 11020 9512
rect 11612 9528 11664 9580
rect 11704 9571 11756 9580
rect 11704 9537 11713 9571
rect 11713 9537 11747 9571
rect 11747 9537 11756 9571
rect 11704 9528 11756 9537
rect 11796 9571 11848 9580
rect 11796 9537 11805 9571
rect 11805 9537 11839 9571
rect 11839 9537 11848 9571
rect 11796 9528 11848 9537
rect 11980 9571 12032 9580
rect 11980 9537 11983 9571
rect 11983 9537 12032 9571
rect 11980 9528 12032 9537
rect 13544 9596 13596 9648
rect 13912 9596 13964 9648
rect 15476 9639 15528 9648
rect 15476 9605 15485 9639
rect 15485 9605 15519 9639
rect 15519 9605 15528 9639
rect 15476 9596 15528 9605
rect 16580 9596 16632 9648
rect 17408 9596 17460 9648
rect 12624 9460 12676 9512
rect 13084 9460 13136 9512
rect 13820 9460 13872 9512
rect 15292 9528 15344 9580
rect 14832 9460 14884 9512
rect 11060 9392 11112 9444
rect 15016 9392 15068 9444
rect 15568 9392 15620 9444
rect 1492 9367 1544 9376
rect 1492 9333 1501 9367
rect 1501 9333 1535 9367
rect 1535 9333 1544 9367
rect 1492 9324 1544 9333
rect 3884 9324 3936 9376
rect 3976 9324 4028 9376
rect 6828 9324 6880 9376
rect 10508 9324 10560 9376
rect 11152 9324 11204 9376
rect 11336 9324 11388 9376
rect 15844 9367 15896 9376
rect 15844 9333 15853 9367
rect 15853 9333 15887 9367
rect 15887 9333 15896 9367
rect 15844 9324 15896 9333
rect 16028 9324 16080 9376
rect 16488 9460 16540 9512
rect 18420 9460 18472 9512
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 16948 9435 17000 9444
rect 16948 9401 16957 9435
rect 16957 9401 16991 9435
rect 16991 9401 17000 9435
rect 16948 9392 17000 9401
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 20214 9222 20266 9274
rect 20278 9222 20330 9274
rect 20342 9222 20394 9274
rect 20406 9222 20458 9274
rect 20470 9222 20522 9274
rect 1492 9120 1544 9172
rect 6000 9120 6052 9172
rect 6460 9120 6512 9172
rect 11612 9120 11664 9172
rect 11704 9120 11756 9172
rect 13820 9120 13872 9172
rect 15016 9120 15068 9172
rect 16396 9120 16448 9172
rect 19432 9120 19484 9172
rect 2136 8984 2188 9036
rect 3424 9052 3476 9104
rect 3976 9027 4028 9036
rect 3976 8993 3985 9027
rect 3985 8993 4019 9027
rect 4019 8993 4028 9027
rect 3976 8984 4028 8993
rect 6460 8916 6512 8968
rect 5540 8848 5592 8900
rect 7656 8984 7708 9036
rect 6828 8959 6880 8968
rect 6828 8925 6837 8959
rect 6837 8925 6871 8959
rect 6871 8925 6880 8959
rect 6828 8916 6880 8925
rect 8944 8959 8996 8968
rect 8944 8925 8953 8959
rect 8953 8925 8987 8959
rect 8987 8925 8996 8959
rect 8944 8916 8996 8925
rect 8852 8780 8904 8832
rect 10968 8916 11020 8968
rect 11060 8959 11112 8968
rect 11060 8925 11069 8959
rect 11069 8925 11103 8959
rect 11103 8925 11112 8959
rect 11060 8916 11112 8925
rect 11336 9027 11388 9036
rect 11336 8993 11345 9027
rect 11345 8993 11379 9027
rect 11379 8993 11388 9027
rect 11336 8984 11388 8993
rect 13084 9095 13136 9104
rect 13084 9061 13093 9095
rect 13093 9061 13127 9095
rect 13127 9061 13136 9095
rect 13084 9052 13136 9061
rect 12808 8984 12860 9036
rect 13268 8916 13320 8968
rect 13544 8916 13596 8968
rect 14924 8959 14976 8968
rect 14924 8925 14933 8959
rect 14933 8925 14967 8959
rect 14967 8925 14976 8959
rect 14924 8916 14976 8925
rect 15476 8959 15528 8968
rect 15476 8925 15485 8959
rect 15485 8925 15519 8959
rect 15519 8925 15528 8959
rect 15476 8916 15528 8925
rect 17224 8916 17276 8968
rect 10692 8823 10744 8832
rect 10692 8789 10701 8823
rect 10701 8789 10735 8823
rect 10735 8789 10744 8823
rect 10692 8780 10744 8789
rect 11704 8780 11756 8832
rect 15568 8848 15620 8900
rect 15844 8848 15896 8900
rect 16396 8848 16448 8900
rect 13268 8780 13320 8832
rect 15200 8780 15252 8832
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 16214 8678 16266 8730
rect 16278 8678 16330 8730
rect 16342 8678 16394 8730
rect 16406 8678 16458 8730
rect 16470 8678 16522 8730
rect 2320 8576 2372 8628
rect 5448 8619 5500 8628
rect 5448 8585 5457 8619
rect 5457 8585 5491 8619
rect 5491 8585 5500 8619
rect 5448 8576 5500 8585
rect 1492 8508 1544 8560
rect 3884 8508 3936 8560
rect 5540 8508 5592 8560
rect 9864 8576 9916 8628
rect 10692 8576 10744 8628
rect 1952 8483 2004 8492
rect 1952 8449 2001 8483
rect 2001 8449 2004 8483
rect 1952 8440 2004 8449
rect 2136 8483 2188 8492
rect 2136 8449 2145 8483
rect 2145 8449 2179 8483
rect 2179 8449 2188 8483
rect 2136 8440 2188 8449
rect 2320 8440 2372 8492
rect 1124 8372 1176 8424
rect 1308 8304 1360 8356
rect 1768 8304 1820 8356
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 3056 8440 3108 8492
rect 3240 8483 3292 8492
rect 3240 8449 3249 8483
rect 3249 8449 3283 8483
rect 3283 8449 3292 8483
rect 3240 8440 3292 8449
rect 3608 8440 3660 8492
rect 3700 8483 3752 8492
rect 3700 8449 3709 8483
rect 3709 8449 3743 8483
rect 3743 8449 3752 8483
rect 3700 8440 3752 8449
rect 8944 8440 8996 8492
rect 9772 8508 9824 8560
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 12624 8576 12676 8628
rect 13084 8576 13136 8628
rect 15476 8576 15528 8628
rect 13268 8551 13320 8560
rect 13268 8517 13277 8551
rect 13277 8517 13311 8551
rect 13311 8517 13320 8551
rect 13268 8508 13320 8517
rect 13544 8508 13596 8560
rect 16028 8508 16080 8560
rect 18420 8619 18472 8628
rect 18420 8585 18429 8619
rect 18429 8585 18463 8619
rect 18463 8585 18472 8619
rect 18420 8576 18472 8585
rect 6368 8415 6420 8424
rect 6368 8381 6377 8415
rect 6377 8381 6411 8415
rect 6411 8381 6420 8415
rect 6368 8372 6420 8381
rect 6736 8372 6788 8424
rect 8300 8415 8352 8424
rect 8300 8381 8309 8415
rect 8309 8381 8343 8415
rect 8343 8381 8352 8415
rect 8300 8372 8352 8381
rect 12072 8440 12124 8492
rect 11612 8372 11664 8424
rect 3700 8304 3752 8356
rect 7012 8236 7064 8288
rect 11704 8304 11756 8356
rect 8116 8279 8168 8288
rect 8116 8245 8125 8279
rect 8125 8245 8159 8279
rect 8159 8245 8168 8279
rect 8116 8236 8168 8245
rect 8760 8279 8812 8288
rect 8760 8245 8769 8279
rect 8769 8245 8803 8279
rect 8803 8245 8812 8279
rect 8760 8236 8812 8245
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 12808 8372 12860 8424
rect 16580 8440 16632 8492
rect 17224 8508 17276 8560
rect 17408 8508 17460 8560
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 15936 8347 15988 8356
rect 15936 8313 15945 8347
rect 15945 8313 15979 8347
rect 15979 8313 15988 8347
rect 15936 8304 15988 8313
rect 13360 8236 13412 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 20214 8134 20266 8186
rect 20278 8134 20330 8186
rect 20342 8134 20394 8186
rect 20406 8134 20458 8186
rect 20470 8134 20522 8186
rect 3056 8032 3108 8084
rect 3608 8032 3660 8084
rect 8300 8032 8352 8084
rect 11152 8032 11204 8084
rect 12900 8032 12952 8084
rect 1492 7871 1544 7880
rect 1492 7837 1501 7871
rect 1501 7837 1535 7871
rect 1535 7837 1544 7871
rect 1492 7828 1544 7837
rect 3424 7828 3476 7880
rect 2044 7803 2096 7812
rect 2044 7769 2053 7803
rect 2053 7769 2087 7803
rect 2087 7769 2096 7803
rect 2044 7760 2096 7769
rect 8116 7896 8168 7948
rect 4160 7828 4212 7880
rect 5816 7828 5868 7880
rect 1584 7692 1636 7744
rect 4712 7803 4764 7812
rect 4712 7769 4721 7803
rect 4721 7769 4755 7803
rect 4755 7769 4764 7803
rect 4712 7760 4764 7769
rect 6460 7871 6512 7880
rect 6460 7837 6469 7871
rect 6469 7837 6503 7871
rect 6503 7837 6512 7871
rect 6460 7828 6512 7837
rect 10784 7896 10836 7948
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 11704 7896 11756 7948
rect 13360 7939 13412 7948
rect 13360 7905 13369 7939
rect 13369 7905 13403 7939
rect 13403 7905 13412 7939
rect 13360 7896 13412 7905
rect 16488 8032 16540 8084
rect 14924 7896 14976 7948
rect 14280 7871 14332 7880
rect 14280 7837 14289 7871
rect 14289 7837 14323 7871
rect 14323 7837 14332 7871
rect 14280 7828 14332 7837
rect 3884 7692 3936 7744
rect 8024 7692 8076 7744
rect 10140 7692 10192 7744
rect 13728 7735 13780 7744
rect 13728 7701 13737 7735
rect 13737 7701 13771 7735
rect 13771 7701 13780 7735
rect 13728 7692 13780 7701
rect 14096 7692 14148 7744
rect 15108 7760 15160 7812
rect 15292 7760 15344 7812
rect 15660 7692 15712 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 16214 7590 16266 7642
rect 16278 7590 16330 7642
rect 16342 7590 16394 7642
rect 16406 7590 16458 7642
rect 16470 7590 16522 7642
rect 2044 7488 2096 7540
rect 4160 7488 4212 7540
rect 4712 7488 4764 7540
rect 6460 7488 6512 7540
rect 6736 7488 6788 7540
rect 10140 7488 10192 7540
rect 11428 7488 11480 7540
rect 13452 7488 13504 7540
rect 3884 7463 3936 7472
rect 3884 7429 3893 7463
rect 3893 7429 3927 7463
rect 3927 7429 3936 7463
rect 3884 7420 3936 7429
rect 6368 7420 6420 7472
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 1676 7327 1728 7336
rect 1676 7293 1685 7327
rect 1685 7293 1719 7327
rect 1719 7293 1728 7327
rect 1676 7284 1728 7293
rect 3240 7352 3292 7404
rect 3148 7284 3200 7336
rect 5724 7352 5776 7404
rect 7012 7395 7064 7404
rect 7012 7361 7021 7395
rect 7021 7361 7055 7395
rect 7055 7361 7064 7395
rect 7012 7352 7064 7361
rect 8116 7420 8168 7472
rect 8760 7420 8812 7472
rect 9220 7420 9272 7472
rect 10048 7420 10100 7472
rect 7656 7395 7708 7404
rect 7656 7361 7660 7395
rect 7660 7361 7694 7395
rect 7694 7361 7708 7395
rect 7656 7352 7708 7361
rect 8024 7395 8076 7404
rect 8024 7361 8033 7395
rect 8033 7361 8067 7395
rect 8067 7361 8076 7395
rect 8024 7352 8076 7361
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 13728 7463 13780 7472
rect 13728 7429 13737 7463
rect 13737 7429 13771 7463
rect 13771 7429 13780 7463
rect 13728 7420 13780 7429
rect 8024 7216 8076 7268
rect 7472 7191 7524 7200
rect 7472 7157 7481 7191
rect 7481 7157 7515 7191
rect 7515 7157 7524 7191
rect 7472 7148 7524 7157
rect 9496 7284 9548 7336
rect 11060 7395 11112 7404
rect 11060 7361 11069 7395
rect 11069 7361 11103 7395
rect 11103 7361 11112 7395
rect 11060 7352 11112 7361
rect 14832 7352 14884 7404
rect 15292 7352 15344 7404
rect 15384 7395 15436 7404
rect 15384 7361 15393 7395
rect 15393 7361 15427 7395
rect 15427 7361 15436 7395
rect 15384 7352 15436 7361
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 12900 7284 12952 7336
rect 10692 7216 10744 7268
rect 9496 7148 9548 7200
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 13452 7327 13504 7336
rect 13452 7293 13461 7327
rect 13461 7293 13495 7327
rect 13495 7293 13504 7327
rect 13452 7284 13504 7293
rect 13820 7284 13872 7336
rect 14280 7284 14332 7336
rect 22100 7284 22152 7336
rect 15384 7216 15436 7268
rect 19984 7216 20036 7268
rect 15844 7148 15896 7200
rect 16028 7148 16080 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 20214 7046 20266 7098
rect 20278 7046 20330 7098
rect 20342 7046 20394 7098
rect 20406 7046 20458 7098
rect 20470 7046 20522 7098
rect 7472 6944 7524 6996
rect 3240 6876 3292 6928
rect 1768 6851 1820 6860
rect 1768 6817 1777 6851
rect 1777 6817 1811 6851
rect 1811 6817 1820 6851
rect 1768 6808 1820 6817
rect 3884 6808 3936 6860
rect 3148 6740 3200 6792
rect 3332 6740 3384 6792
rect 3976 6672 4028 6724
rect 4344 6715 4396 6724
rect 4344 6681 4353 6715
rect 4353 6681 4387 6715
rect 4387 6681 4396 6715
rect 4344 6672 4396 6681
rect 7196 6876 7248 6928
rect 9404 6944 9456 6996
rect 9496 6987 9548 6996
rect 9496 6953 9505 6987
rect 9505 6953 9539 6987
rect 9539 6953 9548 6987
rect 9496 6944 9548 6953
rect 11428 6944 11480 6996
rect 12900 6944 12952 6996
rect 15844 6944 15896 6996
rect 6920 6740 6972 6792
rect 15384 6876 15436 6928
rect 13820 6808 13872 6860
rect 14096 6851 14148 6860
rect 14096 6817 14105 6851
rect 14105 6817 14139 6851
rect 14139 6817 14148 6851
rect 14096 6808 14148 6817
rect 15660 6808 15712 6860
rect 16028 6851 16080 6860
rect 16028 6817 16037 6851
rect 16037 6817 16071 6851
rect 16071 6817 16080 6851
rect 16028 6808 16080 6817
rect 9312 6783 9364 6792
rect 9312 6749 9321 6783
rect 9321 6749 9355 6783
rect 9355 6749 9364 6783
rect 9312 6740 9364 6749
rect 5540 6672 5592 6724
rect 5632 6715 5684 6724
rect 5632 6681 5641 6715
rect 5641 6681 5675 6715
rect 5675 6681 5684 6715
rect 5632 6672 5684 6681
rect 5724 6672 5776 6724
rect 4068 6604 4120 6656
rect 7748 6604 7800 6656
rect 9496 6740 9548 6792
rect 9772 6715 9824 6724
rect 9772 6681 9781 6715
rect 9781 6681 9815 6715
rect 9815 6681 9824 6715
rect 9772 6672 9824 6681
rect 10048 6783 10100 6792
rect 10048 6749 10057 6783
rect 10057 6749 10091 6783
rect 10091 6749 10100 6783
rect 10048 6740 10100 6749
rect 11796 6672 11848 6724
rect 13360 6672 13412 6724
rect 11060 6604 11112 6656
rect 11244 6604 11296 6656
rect 14924 6672 14976 6724
rect 15108 6604 15160 6656
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 16214 6502 16266 6554
rect 16278 6502 16330 6554
rect 16342 6502 16394 6554
rect 16406 6502 16458 6554
rect 16470 6502 16522 6554
rect 1676 6443 1728 6452
rect 1676 6409 1685 6443
rect 1685 6409 1719 6443
rect 1719 6409 1728 6443
rect 1676 6400 1728 6409
rect 3148 6400 3200 6452
rect 3976 6400 4028 6452
rect 5540 6443 5592 6452
rect 5540 6409 5549 6443
rect 5549 6409 5583 6443
rect 5583 6409 5592 6443
rect 5540 6400 5592 6409
rect 6736 6400 6788 6452
rect 1584 6307 1636 6316
rect 1584 6273 1593 6307
rect 1593 6273 1627 6307
rect 1627 6273 1636 6307
rect 1584 6264 1636 6273
rect 3608 6332 3660 6384
rect 3792 6332 3844 6384
rect 4068 6375 4120 6384
rect 4068 6341 4077 6375
rect 4077 6341 4111 6375
rect 4111 6341 4120 6375
rect 4068 6332 4120 6341
rect 5632 6332 5684 6384
rect 9312 6400 9364 6452
rect 10048 6400 10100 6452
rect 1952 6264 2004 6316
rect 2136 6307 2188 6316
rect 2136 6273 2140 6307
rect 2140 6273 2174 6307
rect 2174 6273 2188 6307
rect 2136 6264 2188 6273
rect 2228 6307 2280 6316
rect 2228 6273 2237 6307
rect 2237 6273 2271 6307
rect 2271 6273 2280 6307
rect 2228 6264 2280 6273
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 1032 6196 1084 6248
rect 2780 6307 2832 6316
rect 2780 6273 2789 6307
rect 2789 6273 2823 6307
rect 2823 6273 2832 6307
rect 2780 6264 2832 6273
rect 3056 6307 3108 6316
rect 3056 6273 3065 6307
rect 3065 6273 3099 6307
rect 3099 6273 3108 6307
rect 3056 6264 3108 6273
rect 3148 6307 3200 6316
rect 3148 6273 3157 6307
rect 3157 6273 3191 6307
rect 3191 6273 3200 6307
rect 3148 6264 3200 6273
rect 5724 6264 5776 6316
rect 7748 6375 7800 6384
rect 7748 6341 7757 6375
rect 7757 6341 7791 6375
rect 7791 6341 7800 6375
rect 7748 6332 7800 6341
rect 1492 6128 1544 6180
rect 2228 6128 2280 6180
rect 2780 6128 2832 6180
rect 3148 6128 3200 6180
rect 3332 6128 3384 6180
rect 6552 6196 6604 6248
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 7196 6307 7248 6316
rect 7196 6273 7205 6307
rect 7205 6273 7239 6307
rect 7239 6273 7248 6307
rect 7196 6264 7248 6273
rect 8760 6264 8812 6316
rect 11428 6400 11480 6452
rect 11244 6332 11296 6384
rect 13360 6332 13412 6384
rect 14924 6332 14976 6384
rect 10784 6264 10836 6316
rect 11152 6264 11204 6316
rect 6920 6196 6972 6248
rect 5448 6128 5500 6180
rect 9772 6196 9824 6248
rect 11980 6196 12032 6248
rect 2688 6103 2740 6112
rect 2688 6069 2697 6103
rect 2697 6069 2731 6103
rect 2731 6069 2740 6103
rect 2688 6060 2740 6069
rect 3056 6060 3108 6112
rect 4252 6060 4304 6112
rect 7104 6060 7156 6112
rect 9680 6060 9732 6112
rect 10048 6060 10100 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 20214 5958 20266 6010
rect 20278 5958 20330 6010
rect 20342 5958 20394 6010
rect 20406 5958 20458 6010
rect 20470 5958 20522 6010
rect 2136 5856 2188 5908
rect 2688 5720 2740 5772
rect 5448 5856 5500 5908
rect 6552 5856 6604 5908
rect 3608 5788 3660 5840
rect 5724 5788 5776 5840
rect 6920 5788 6972 5840
rect 3884 5720 3936 5772
rect 3332 5652 3384 5704
rect 4068 5652 4120 5704
rect 5540 5763 5592 5772
rect 5540 5729 5549 5763
rect 5549 5729 5583 5763
rect 5583 5729 5592 5763
rect 5540 5720 5592 5729
rect 7656 5899 7708 5908
rect 7656 5865 7665 5899
rect 7665 5865 7699 5899
rect 7699 5865 7708 5899
rect 7656 5856 7708 5865
rect 9772 5856 9824 5908
rect 11980 5856 12032 5908
rect 13544 5856 13596 5908
rect 7380 5788 7432 5840
rect 10140 5788 10192 5840
rect 2044 5627 2096 5636
rect 2044 5593 2053 5627
rect 2053 5593 2087 5627
rect 2087 5593 2096 5627
rect 2044 5584 2096 5593
rect 3424 5584 3476 5636
rect 3608 5584 3660 5636
rect 3792 5584 3844 5636
rect 4712 5627 4764 5636
rect 4712 5593 4721 5627
rect 4721 5593 4755 5627
rect 4755 5593 4764 5627
rect 4712 5584 4764 5593
rect 6184 5695 6236 5704
rect 6184 5661 6193 5695
rect 6193 5661 6227 5695
rect 6227 5661 6236 5695
rect 6184 5652 6236 5661
rect 7104 5695 7156 5704
rect 7104 5661 7113 5695
rect 7113 5661 7147 5695
rect 7147 5661 7156 5695
rect 7104 5652 7156 5661
rect 10048 5763 10100 5772
rect 10048 5729 10057 5763
rect 10057 5729 10091 5763
rect 10091 5729 10100 5763
rect 10048 5720 10100 5729
rect 11060 5720 11112 5772
rect 11336 5720 11388 5772
rect 11704 5720 11756 5772
rect 7564 5695 7616 5704
rect 7564 5661 7567 5695
rect 7567 5661 7616 5695
rect 7564 5652 7616 5661
rect 6552 5584 6604 5636
rect 6736 5584 6788 5636
rect 8576 5652 8628 5704
rect 11796 5652 11848 5704
rect 12532 5652 12584 5704
rect 12716 5652 12768 5704
rect 14924 5652 14976 5704
rect 8852 5584 8904 5636
rect 10692 5627 10744 5636
rect 10692 5593 10701 5627
rect 10701 5593 10735 5627
rect 10735 5593 10744 5627
rect 10692 5584 10744 5593
rect 2320 5516 2372 5568
rect 3056 5516 3108 5568
rect 6276 5516 6328 5568
rect 6920 5516 6972 5568
rect 7104 5516 7156 5568
rect 8668 5559 8720 5568
rect 8668 5525 8677 5559
rect 8677 5525 8711 5559
rect 8711 5525 8720 5559
rect 8668 5516 8720 5525
rect 9036 5559 9088 5568
rect 9036 5525 9045 5559
rect 9045 5525 9079 5559
rect 9079 5525 9088 5559
rect 9036 5516 9088 5525
rect 9312 5516 9364 5568
rect 12716 5516 12768 5568
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 16214 5414 16266 5466
rect 16278 5414 16330 5466
rect 16342 5414 16394 5466
rect 16406 5414 16458 5466
rect 16470 5414 16522 5466
rect 2044 5312 2096 5364
rect 3424 5312 3476 5364
rect 6552 5312 6604 5364
rect 7564 5312 7616 5364
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 9680 5312 9732 5364
rect 4068 5244 4120 5296
rect 4712 5244 4764 5296
rect 8760 5244 8812 5296
rect 9956 5244 10008 5296
rect 10784 5244 10836 5296
rect 3332 5219 3384 5228
rect 3332 5185 3341 5219
rect 3341 5185 3375 5219
rect 3375 5185 3384 5219
rect 3332 5176 3384 5185
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 3976 5219 4028 5228
rect 3976 5185 3990 5219
rect 3990 5185 4024 5219
rect 4024 5185 4028 5219
rect 3976 5176 4028 5185
rect 5724 5176 5776 5228
rect 3884 5040 3936 5092
rect 3792 4972 3844 5024
rect 4068 4972 4120 5024
rect 6368 4972 6420 5024
rect 6736 4972 6788 5024
rect 7104 5219 7156 5228
rect 7104 5185 7113 5219
rect 7113 5185 7147 5219
rect 7147 5185 7156 5219
rect 7104 5176 7156 5185
rect 9036 5176 9088 5228
rect 12532 5244 12584 5296
rect 13544 5244 13596 5296
rect 14924 5244 14976 5296
rect 7748 5108 7800 5160
rect 10048 5108 10100 5160
rect 10140 5108 10192 5160
rect 12624 5219 12676 5228
rect 12624 5185 12633 5219
rect 12633 5185 12667 5219
rect 12667 5185 12676 5219
rect 12624 5176 12676 5185
rect 13084 5176 13136 5228
rect 13636 5151 13688 5160
rect 13636 5117 13645 5151
rect 13645 5117 13679 5151
rect 13679 5117 13688 5151
rect 13636 5108 13688 5117
rect 11704 5083 11756 5092
rect 11704 5049 11713 5083
rect 11713 5049 11747 5083
rect 11747 5049 11756 5083
rect 11704 5040 11756 5049
rect 9312 4972 9364 5024
rect 11612 5015 11664 5024
rect 11612 4981 11621 5015
rect 11621 4981 11655 5015
rect 11655 4981 11664 5015
rect 11612 4972 11664 4981
rect 11796 4972 11848 5024
rect 13452 4972 13504 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 20214 4870 20266 4922
rect 20278 4870 20330 4922
rect 20342 4870 20394 4922
rect 20406 4870 20458 4922
rect 20470 4870 20522 4922
rect 3884 4768 3936 4820
rect 6000 4768 6052 4820
rect 6644 4768 6696 4820
rect 12716 4768 12768 4820
rect 13636 4768 13688 4820
rect 3332 4632 3384 4684
rect 3792 4675 3844 4684
rect 3792 4641 3801 4675
rect 3801 4641 3835 4675
rect 3835 4641 3844 4675
rect 3792 4632 3844 4641
rect 7748 4743 7800 4752
rect 7748 4709 7757 4743
rect 7757 4709 7791 4743
rect 7791 4709 7800 4743
rect 7748 4700 7800 4709
rect 5540 4632 5592 4684
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 3148 4564 3200 4616
rect 2044 4539 2096 4548
rect 2044 4505 2053 4539
rect 2053 4505 2087 4539
rect 2087 4505 2096 4539
rect 2044 4496 2096 4505
rect 5908 4607 5960 4616
rect 5908 4573 5917 4607
rect 5917 4573 5951 4607
rect 5951 4573 5960 4607
rect 5908 4564 5960 4573
rect 4436 4428 4488 4480
rect 4712 4428 4764 4480
rect 5816 4471 5868 4480
rect 5816 4437 5825 4471
rect 5825 4437 5859 4471
rect 5859 4437 5868 4471
rect 5816 4428 5868 4437
rect 6828 4496 6880 4548
rect 8116 4564 8168 4616
rect 11612 4632 11664 4684
rect 12716 4632 12768 4684
rect 13360 4632 13412 4684
rect 9220 4564 9272 4616
rect 9588 4564 9640 4616
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 14280 4607 14332 4616
rect 14280 4573 14289 4607
rect 14289 4573 14323 4607
rect 14323 4573 14332 4607
rect 14280 4564 14332 4573
rect 8760 4496 8812 4548
rect 10876 4496 10928 4548
rect 13084 4496 13136 4548
rect 8852 4428 8904 4480
rect 9680 4471 9732 4480
rect 9680 4437 9689 4471
rect 9689 4437 9723 4471
rect 9723 4437 9732 4471
rect 9680 4428 9732 4437
rect 12072 4428 12124 4480
rect 14096 4428 14148 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 16214 4326 16266 4378
rect 16278 4326 16330 4378
rect 16342 4326 16394 4378
rect 16406 4326 16458 4378
rect 16470 4326 16522 4378
rect 2044 4224 2096 4276
rect 2964 4224 3016 4276
rect 2136 4088 2188 4140
rect 4436 4156 4488 4208
rect 5540 4156 5592 4208
rect 6736 4156 6788 4208
rect 10048 4224 10100 4276
rect 13544 4267 13596 4276
rect 13544 4233 13553 4267
rect 13553 4233 13587 4267
rect 13587 4233 13596 4267
rect 13544 4224 13596 4233
rect 9956 4156 10008 4208
rect 10784 4156 10836 4208
rect 12072 4199 12124 4208
rect 12072 4165 12081 4199
rect 12081 4165 12115 4199
rect 12115 4165 12124 4199
rect 12072 4156 12124 4165
rect 3056 4131 3108 4140
rect 3056 4097 3060 4131
rect 3060 4097 3094 4131
rect 3094 4097 3108 4131
rect 3056 4088 3108 4097
rect 3516 4131 3568 4140
rect 2780 4020 2832 4072
rect 2964 4020 3016 4072
rect 3516 4097 3525 4131
rect 3525 4097 3559 4131
rect 3559 4097 3568 4131
rect 3516 4088 3568 4097
rect 3700 4088 3752 4140
rect 3884 4131 3936 4140
rect 3884 4097 3893 4131
rect 3893 4097 3927 4131
rect 3927 4097 3936 4131
rect 3884 4088 3936 4097
rect 3608 4020 3660 4072
rect 6000 4131 6052 4140
rect 6000 4097 6009 4131
rect 6009 4097 6043 4131
rect 6043 4097 6052 4131
rect 6000 4088 6052 4097
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 1308 3884 1360 3936
rect 2412 3995 2464 4004
rect 2412 3961 2421 3995
rect 2421 3961 2455 3995
rect 2455 3961 2464 3995
rect 2412 3952 2464 3961
rect 3240 3952 3292 4004
rect 3608 3927 3660 3936
rect 3608 3893 3617 3927
rect 3617 3893 3651 3927
rect 3651 3893 3660 3927
rect 3608 3884 3660 3893
rect 5264 3884 5316 3936
rect 6736 4063 6788 4072
rect 6736 4029 6745 4063
rect 6745 4029 6779 4063
rect 6779 4029 6788 4063
rect 6736 4020 6788 4029
rect 8668 4063 8720 4072
rect 8668 4029 8677 4063
rect 8677 4029 8711 4063
rect 8711 4029 8720 4063
rect 8668 4020 8720 4029
rect 8760 4020 8812 4072
rect 11796 4131 11848 4140
rect 11796 4097 11805 4131
rect 11805 4097 11839 4131
rect 11839 4097 11848 4131
rect 11796 4088 11848 4097
rect 13084 4088 13136 4140
rect 10416 4020 10468 4072
rect 13912 4131 13964 4140
rect 13912 4097 13921 4131
rect 13921 4097 13955 4131
rect 13955 4097 13964 4131
rect 13912 4088 13964 4097
rect 13268 4020 13320 4072
rect 14924 4063 14976 4072
rect 14924 4029 14933 4063
rect 14933 4029 14967 4063
rect 14967 4029 14976 4063
rect 14924 4020 14976 4029
rect 15660 4020 15712 4072
rect 6920 3884 6972 3936
rect 8116 3884 8168 3936
rect 10048 3952 10100 4004
rect 10968 3952 11020 4004
rect 8760 3884 8812 3936
rect 10416 3927 10468 3936
rect 10416 3893 10425 3927
rect 10425 3893 10459 3927
rect 10459 3893 10468 3927
rect 10416 3884 10468 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 20214 3782 20266 3834
rect 20278 3782 20330 3834
rect 20342 3782 20394 3834
rect 20406 3782 20458 3834
rect 20470 3782 20522 3834
rect 2780 3680 2832 3732
rect 3332 3680 3384 3732
rect 4528 3612 4580 3664
rect 6736 3680 6788 3732
rect 9036 3680 9088 3732
rect 9496 3680 9548 3732
rect 3056 3544 3108 3596
rect 3148 3476 3200 3528
rect 3424 3476 3476 3528
rect 3884 3544 3936 3596
rect 4712 3544 4764 3596
rect 5816 3544 5868 3596
rect 6552 3544 6604 3596
rect 10968 3612 11020 3664
rect 8576 3544 8628 3596
rect 11888 3544 11940 3596
rect 2044 3451 2096 3460
rect 2044 3417 2053 3451
rect 2053 3417 2087 3451
rect 2087 3417 2096 3451
rect 2044 3408 2096 3417
rect 2964 3340 3016 3392
rect 4804 3519 4856 3528
rect 4804 3485 4813 3519
rect 4813 3485 4847 3519
rect 4847 3485 4856 3519
rect 4804 3476 4856 3485
rect 8944 3519 8996 3528
rect 8944 3485 8953 3519
rect 8953 3485 8987 3519
rect 8987 3485 8996 3519
rect 8944 3476 8996 3485
rect 9036 3476 9088 3528
rect 3700 3340 3752 3392
rect 4620 3408 4672 3460
rect 5264 3451 5316 3460
rect 5264 3417 5273 3451
rect 5273 3417 5307 3451
rect 5307 3417 5316 3451
rect 5264 3408 5316 3417
rect 5448 3340 5500 3392
rect 5632 3340 5684 3392
rect 6828 3408 6880 3460
rect 8668 3408 8720 3460
rect 8852 3340 8904 3392
rect 8944 3340 8996 3392
rect 9680 3408 9732 3460
rect 10784 3408 10836 3460
rect 11980 3451 12032 3460
rect 11980 3417 11989 3451
rect 11989 3417 12023 3451
rect 12023 3417 12032 3451
rect 11980 3408 12032 3417
rect 9956 3340 10008 3392
rect 13084 3408 13136 3460
rect 14096 3587 14148 3596
rect 14096 3553 14105 3587
rect 14105 3553 14139 3587
rect 14139 3553 14148 3587
rect 14096 3544 14148 3553
rect 14280 3408 14332 3460
rect 15660 3408 15712 3460
rect 15844 3383 15896 3392
rect 15844 3349 15853 3383
rect 15853 3349 15887 3383
rect 15887 3349 15896 3383
rect 15844 3340 15896 3349
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 16214 3238 16266 3290
rect 16278 3238 16330 3290
rect 16342 3238 16394 3290
rect 16406 3238 16458 3290
rect 16470 3238 16522 3290
rect 1492 3136 1544 3188
rect 2780 3068 2832 3120
rect 3148 3068 3200 3120
rect 3700 3043 3752 3052
rect 3700 3009 3704 3043
rect 3704 3009 3738 3043
rect 3738 3009 3752 3043
rect 3700 3000 3752 3009
rect 3792 3043 3844 3052
rect 3792 3009 3801 3043
rect 3801 3009 3835 3043
rect 3835 3009 3844 3043
rect 3792 3000 3844 3009
rect 4712 3068 4764 3120
rect 6828 3136 6880 3188
rect 8576 3136 8628 3188
rect 9588 3136 9640 3188
rect 8300 3068 8352 3120
rect 8668 3068 8720 3120
rect 9956 3068 10008 3120
rect 4068 3043 4120 3052
rect 4068 3009 4077 3043
rect 4077 3009 4111 3043
rect 4111 3009 4120 3043
rect 4068 3000 4120 3009
rect 10416 3068 10468 3120
rect 10968 3000 11020 3052
rect 14280 3068 14332 3120
rect 11520 3000 11572 3052
rect 13268 3000 13320 3052
rect 2044 2932 2096 2984
rect 3056 2975 3108 2984
rect 3056 2941 3065 2975
rect 3065 2941 3099 2975
rect 3099 2941 3108 2975
rect 3056 2932 3108 2941
rect 3516 2839 3568 2848
rect 3516 2805 3525 2839
rect 3525 2805 3559 2839
rect 3559 2805 3568 2839
rect 3516 2796 3568 2805
rect 3884 2796 3936 2848
rect 4160 2932 4212 2984
rect 6460 2975 6512 2984
rect 6460 2941 6469 2975
rect 6469 2941 6503 2975
rect 6503 2941 6512 2975
rect 6460 2932 6512 2941
rect 8116 2932 8168 2984
rect 10508 2932 10560 2984
rect 12624 2932 12676 2984
rect 14924 3043 14976 3052
rect 14924 3009 14933 3043
rect 14933 3009 14967 3043
rect 14967 3009 14976 3043
rect 14924 3000 14976 3009
rect 15844 3136 15896 3188
rect 4620 2796 4672 2848
rect 8944 2864 8996 2916
rect 11060 2907 11112 2916
rect 11060 2873 11069 2907
rect 11069 2873 11103 2907
rect 11103 2873 11112 2907
rect 11060 2864 11112 2873
rect 9220 2796 9272 2848
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 11980 2796 12032 2848
rect 13544 2932 13596 2984
rect 13360 2864 13412 2916
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 15660 2796 15712 2848
rect 22192 2796 22244 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 20214 2694 20266 2746
rect 20278 2694 20330 2746
rect 20342 2694 20394 2746
rect 20406 2694 20458 2746
rect 20470 2694 20522 2746
rect 4528 2592 4580 2644
rect 4712 2592 4764 2644
rect 5724 2592 5776 2644
rect 3332 2524 3384 2576
rect 10140 2592 10192 2644
rect 3516 2456 3568 2508
rect 3608 2456 3660 2508
rect 1492 2431 1544 2440
rect 1492 2397 1501 2431
rect 1501 2397 1535 2431
rect 1535 2397 1544 2431
rect 1492 2388 1544 2397
rect 5724 2388 5776 2440
rect 2044 2363 2096 2372
rect 2044 2329 2053 2363
rect 2053 2329 2087 2363
rect 2087 2329 2096 2363
rect 2044 2320 2096 2329
rect 2780 2320 2832 2372
rect 2136 2252 2188 2304
rect 4620 2320 4672 2372
rect 5540 2252 5592 2304
rect 6092 2252 6144 2304
rect 8576 2456 8628 2508
rect 9772 2524 9824 2576
rect 10048 2567 10100 2576
rect 10048 2533 10057 2567
rect 10057 2533 10091 2567
rect 10091 2533 10100 2567
rect 10048 2524 10100 2533
rect 8300 2388 8352 2440
rect 9036 2431 9088 2440
rect 9036 2397 9045 2431
rect 9045 2397 9079 2431
rect 9079 2397 9088 2431
rect 9036 2388 9088 2397
rect 9404 2431 9456 2440
rect 9404 2397 9418 2431
rect 9418 2397 9452 2431
rect 9452 2397 9456 2431
rect 9404 2388 9456 2397
rect 6828 2320 6880 2372
rect 8668 2295 8720 2304
rect 8668 2261 8677 2295
rect 8677 2261 8711 2295
rect 8711 2261 8720 2295
rect 8668 2252 8720 2261
rect 8944 2320 8996 2372
rect 10324 2388 10376 2440
rect 12348 2592 12400 2644
rect 12624 2592 12676 2644
rect 12716 2592 12768 2644
rect 13912 2592 13964 2644
rect 14004 2592 14056 2644
rect 11980 2524 12032 2576
rect 14188 2524 14240 2576
rect 11060 2456 11112 2508
rect 11612 2456 11664 2508
rect 13728 2456 13780 2508
rect 13912 2456 13964 2508
rect 13820 2431 13872 2440
rect 13820 2397 13829 2431
rect 13829 2397 13863 2431
rect 13863 2397 13872 2431
rect 13820 2388 13872 2397
rect 14096 2431 14148 2440
rect 14096 2397 14105 2431
rect 14105 2397 14139 2431
rect 14139 2397 14148 2431
rect 14096 2388 14148 2397
rect 9496 2252 9548 2304
rect 10600 2252 10652 2304
rect 10968 2320 11020 2372
rect 12256 2320 12308 2372
rect 11060 2252 11112 2304
rect 11888 2252 11940 2304
rect 22100 2320 22152 2372
rect 23020 2320 23072 2372
rect 13728 2252 13780 2304
rect 15016 2252 15068 2304
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 16214 2150 16266 2202
rect 16278 2150 16330 2202
rect 16342 2150 16394 2202
rect 16406 2150 16458 2202
rect 16470 2150 16522 2202
rect 2044 2048 2096 2100
rect 3424 2048 3476 2100
rect 3976 2048 4028 2100
rect 6460 2048 6512 2100
rect 6644 2048 6696 2100
rect 2872 1980 2924 2032
rect 4620 1980 4672 2032
rect 6552 2023 6604 2032
rect 6552 1989 6561 2023
rect 6561 1989 6595 2023
rect 6595 1989 6604 2023
rect 6552 1980 6604 1989
rect 8300 1980 8352 2032
rect 9404 2048 9456 2100
rect 11520 2048 11572 2100
rect 11612 1980 11664 2032
rect 11888 1980 11940 2032
rect 11980 2023 12032 2032
rect 11980 1989 11989 2023
rect 11989 1989 12023 2023
rect 12023 1989 12032 2023
rect 11980 1980 12032 1989
rect 2136 1955 2188 1964
rect 2136 1921 2145 1955
rect 2145 1921 2179 1955
rect 2179 1921 2188 1955
rect 2136 1912 2188 1921
rect 3976 1912 4028 1964
rect 4068 1955 4120 1964
rect 4068 1921 4077 1955
rect 4077 1921 4111 1955
rect 4111 1921 4120 1955
rect 4068 1912 4120 1921
rect 5908 1912 5960 1964
rect 2412 1887 2464 1896
rect 2412 1853 2421 1887
rect 2421 1853 2455 1887
rect 2455 1853 2464 1887
rect 2412 1844 2464 1853
rect 2780 1844 2832 1896
rect 1768 1819 1820 1828
rect 1768 1785 1777 1819
rect 1777 1785 1811 1819
rect 1811 1785 1820 1819
rect 1768 1776 1820 1785
rect 4160 1844 4212 1896
rect 4620 1887 4672 1896
rect 4620 1853 4629 1887
rect 4629 1853 4663 1887
rect 4663 1853 4672 1887
rect 4620 1844 4672 1853
rect 6000 1844 6052 1896
rect 6736 1955 6788 1964
rect 6736 1921 6750 1955
rect 6750 1921 6784 1955
rect 6784 1921 6788 1955
rect 6736 1912 6788 1921
rect 12624 1912 12676 1964
rect 14924 2048 14976 2100
rect 15016 2048 15068 2100
rect 14188 1912 14240 1964
rect 15016 1912 15068 1964
rect 20260 1955 20312 1964
rect 20260 1921 20269 1955
rect 20269 1921 20303 1955
rect 20303 1921 20312 1955
rect 20260 1912 20312 1921
rect 22192 1912 22244 1964
rect 7840 1887 7892 1896
rect 7840 1853 7849 1887
rect 7849 1853 7883 1887
rect 7883 1853 7892 1887
rect 7840 1844 7892 1853
rect 9496 1887 9548 1896
rect 9496 1853 9505 1887
rect 9505 1853 9539 1887
rect 9539 1853 9548 1887
rect 9496 1844 9548 1853
rect 10508 1844 10560 1896
rect 10784 1844 10836 1896
rect 12072 1844 12124 1896
rect 13544 1844 13596 1896
rect 14556 1887 14608 1896
rect 14556 1853 14565 1887
rect 14565 1853 14599 1887
rect 14599 1853 14608 1887
rect 14556 1844 14608 1853
rect 15660 1887 15712 1896
rect 15660 1853 15669 1887
rect 15669 1853 15703 1887
rect 15703 1853 15712 1887
rect 15660 1844 15712 1853
rect 17500 1887 17552 1896
rect 17500 1853 17509 1887
rect 17509 1853 17543 1887
rect 17543 1853 17552 1887
rect 17500 1844 17552 1853
rect 19340 1887 19392 1896
rect 19340 1853 19349 1887
rect 19349 1853 19383 1887
rect 19383 1853 19392 1887
rect 19340 1844 19392 1853
rect 21180 1887 21232 1896
rect 21180 1853 21189 1887
rect 21189 1853 21223 1887
rect 21223 1853 21232 1887
rect 21180 1844 21232 1853
rect 6736 1776 6788 1828
rect 6920 1819 6972 1828
rect 6920 1785 6929 1819
rect 6929 1785 6963 1819
rect 6963 1785 6972 1819
rect 6920 1776 6972 1785
rect 10140 1708 10192 1760
rect 14648 1708 14700 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 20214 1606 20266 1658
rect 20278 1606 20330 1658
rect 20342 1606 20394 1658
rect 20406 1606 20458 1658
rect 20470 1606 20522 1658
rect 2412 1504 2464 1556
rect 2872 1504 2924 1556
rect 4620 1504 4672 1556
rect 5632 1504 5684 1556
rect 7840 1504 7892 1556
rect 8300 1504 8352 1556
rect 3976 1436 4028 1488
rect 8668 1504 8720 1556
rect 11244 1504 11296 1556
rect 15016 1504 15068 1556
rect 9864 1436 9916 1488
rect 940 1300 992 1352
rect 1492 1300 1544 1352
rect 2872 1232 2924 1284
rect 3792 1300 3844 1352
rect 3976 1300 4028 1352
rect 6368 1368 6420 1420
rect 6736 1368 6788 1420
rect 8944 1368 8996 1420
rect 9036 1368 9088 1420
rect 5724 1343 5776 1352
rect 5724 1309 5733 1343
rect 5733 1309 5767 1343
rect 5767 1309 5776 1343
rect 5724 1300 5776 1309
rect 5908 1343 5960 1352
rect 5908 1309 5917 1343
rect 5917 1309 5951 1343
rect 5951 1309 5960 1343
rect 5908 1300 5960 1309
rect 6000 1300 6052 1352
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 11060 1368 11112 1420
rect 11520 1411 11572 1420
rect 11520 1377 11529 1411
rect 11529 1377 11563 1411
rect 11563 1377 11572 1411
rect 11520 1368 11572 1377
rect 4068 1232 4120 1284
rect 8300 1232 8352 1284
rect 9772 1232 9824 1284
rect 10968 1232 11020 1284
rect 5816 1207 5868 1216
rect 5816 1173 5825 1207
rect 5825 1173 5859 1207
rect 5859 1173 5868 1207
rect 5816 1164 5868 1173
rect 10416 1164 10468 1216
rect 14648 1343 14700 1352
rect 14648 1309 14657 1343
rect 14657 1309 14691 1343
rect 14691 1309 14700 1343
rect 14648 1300 14700 1309
rect 12532 1232 12584 1284
rect 14556 1164 14608 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 16214 1062 16266 1114
rect 16278 1062 16330 1114
rect 16342 1062 16394 1114
rect 16406 1062 16458 1114
rect 16470 1062 16522 1114
rect 1768 960 1820 1012
rect 5724 960 5776 1012
<< metal2 >>
rect 1030 14362 1086 15000
rect 2318 14362 2374 15000
rect 3606 14362 3662 15000
rect 1030 14334 1164 14362
rect 1030 14200 1086 14334
rect 1136 8430 1164 14334
rect 2318 14334 2636 14362
rect 2318 14200 2374 14334
rect 1492 13184 1544 13190
rect 1492 13126 1544 13132
rect 1504 12918 1532 13126
rect 1492 12912 1544 12918
rect 1492 12854 1544 12860
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 1768 12708 1820 12714
rect 1768 12650 1820 12656
rect 1676 12232 1728 12238
rect 1676 12174 1728 12180
rect 1688 11762 1716 12174
rect 1676 11756 1728 11762
rect 1676 11698 1728 11704
rect 1688 10810 1716 11698
rect 1780 11676 1808 12650
rect 2044 12640 2096 12646
rect 2044 12582 2096 12588
rect 2056 12170 2084 12582
rect 2240 12442 2268 12718
rect 2228 12436 2280 12442
rect 2228 12378 2280 12384
rect 2412 12436 2464 12442
rect 2412 12378 2464 12384
rect 2044 12164 2096 12170
rect 2044 12106 2096 12112
rect 2424 11694 2452 12378
rect 1860 11688 1912 11694
rect 1780 11648 1860 11676
rect 1780 11529 1808 11648
rect 1860 11630 1912 11636
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 1766 11520 1822 11529
rect 1766 11455 1822 11464
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 1688 10674 1716 10746
rect 1676 10668 1728 10674
rect 1676 10610 1728 10616
rect 1952 10600 2004 10606
rect 1952 10542 2004 10548
rect 1964 10266 1992 10542
rect 1952 10260 2004 10266
rect 1952 10202 2004 10208
rect 2504 10192 2556 10198
rect 2504 10134 2556 10140
rect 2516 10062 2544 10134
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2504 10056 2556 10062
rect 2504 9998 2556 10004
rect 2044 9920 2096 9926
rect 2044 9862 2096 9868
rect 2056 9586 2084 9862
rect 2044 9580 2096 9586
rect 2044 9522 2096 9528
rect 1308 9444 1360 9450
rect 1308 9386 1360 9392
rect 1124 8424 1176 8430
rect 1124 8366 1176 8372
rect 1136 6914 1164 8366
rect 1320 8362 1348 9386
rect 1492 9376 1544 9382
rect 1492 9318 1544 9324
rect 1504 9178 1532 9318
rect 1492 9172 1544 9178
rect 1492 9114 1544 9120
rect 2148 9042 2176 9998
rect 2516 9722 2544 9998
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2332 8634 2360 9454
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 1492 8560 1544 8566
rect 1492 8502 1544 8508
rect 1308 8356 1360 8362
rect 1308 8298 1360 8304
rect 1044 6886 1164 6914
rect 1044 6254 1072 6886
rect 1032 6248 1084 6254
rect 1032 6190 1084 6196
rect 1320 5817 1348 8298
rect 1504 7886 1532 8502
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 2320 8492 2372 8498
rect 2320 8434 2372 8440
rect 1768 8356 1820 8362
rect 1768 8298 1820 8304
rect 1582 8256 1638 8265
rect 1582 8191 1638 8200
rect 1492 7880 1544 7886
rect 1492 7822 1544 7828
rect 1400 7404 1452 7410
rect 1504 7392 1532 7822
rect 1596 7750 1624 8191
rect 1584 7744 1636 7750
rect 1584 7686 1636 7692
rect 1452 7364 1532 7392
rect 1400 7346 1452 7352
rect 1504 6186 1532 7364
rect 1596 6322 1624 7686
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1688 6458 1716 7278
rect 1780 6866 1808 8298
rect 1768 6860 1820 6866
rect 1768 6802 1820 6808
rect 1676 6452 1728 6458
rect 1676 6394 1728 6400
rect 1964 6322 1992 8434
rect 2044 7812 2096 7818
rect 2044 7754 2096 7760
rect 2056 7546 2084 7754
rect 2044 7540 2096 7546
rect 2044 7482 2096 7488
rect 2148 6914 2176 8434
rect 2148 6886 2268 6914
rect 2240 6322 2268 6886
rect 2332 6322 2360 8434
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1952 6316 2004 6322
rect 1952 6258 2004 6264
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2228 6316 2280 6322
rect 2228 6258 2280 6264
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 1492 6180 1544 6186
rect 1492 6122 1544 6128
rect 2148 5914 2176 6258
rect 2240 6186 2268 6258
rect 2228 6180 2280 6186
rect 2228 6122 2280 6128
rect 2136 5908 2188 5914
rect 2136 5850 2188 5856
rect 1306 5808 1362 5817
rect 1306 5743 1362 5752
rect 2044 5636 2096 5642
rect 2044 5578 2096 5584
rect 2056 5370 2084 5578
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2044 4548 2096 4554
rect 2044 4490 2096 4496
rect 2056 4282 2084 4490
rect 2044 4276 2096 4282
rect 2044 4218 2096 4224
rect 2148 4146 2176 5850
rect 2332 5574 2360 6258
rect 2320 5568 2372 5574
rect 2320 5510 2372 5516
rect 2410 4176 2466 4185
rect 2136 4140 2188 4146
rect 2410 4111 2466 4120
rect 2136 4082 2188 4088
rect 2424 4010 2452 4111
rect 2412 4004 2464 4010
rect 2412 3946 2464 3952
rect 1308 3936 1360 3942
rect 1308 3878 1360 3884
rect 1320 3369 1348 3878
rect 2424 3641 2452 3946
rect 2410 3632 2466 3641
rect 2410 3567 2466 3576
rect 2044 3460 2096 3466
rect 2044 3402 2096 3408
rect 1306 3360 1362 3369
rect 1306 3295 1362 3304
rect 1492 3188 1544 3194
rect 1492 3130 1544 3136
rect 1504 2446 1532 3130
rect 2056 2990 2084 3402
rect 2044 2984 2096 2990
rect 2044 2926 2096 2932
rect 1766 2544 1822 2553
rect 1766 2479 1822 2488
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1504 1358 1532 2382
rect 1780 1834 1808 2479
rect 2608 2417 2636 14334
rect 3528 14334 3662 14362
rect 2964 13252 3016 13258
rect 2964 13194 3016 13200
rect 2780 12300 2832 12306
rect 2780 12242 2832 12248
rect 2792 11830 2820 12242
rect 2976 11898 3004 13194
rect 3148 13184 3200 13190
rect 3148 13126 3200 13132
rect 3332 13184 3384 13190
rect 3332 13126 3384 13132
rect 3160 12782 3188 13126
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 3160 12238 3188 12718
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2964 11892 3016 11898
rect 2964 11834 3016 11840
rect 2780 11824 2832 11830
rect 2780 11766 2832 11772
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2700 11218 2728 11630
rect 2792 11354 2820 11766
rect 3344 11762 3372 13126
rect 3332 11756 3384 11762
rect 3332 11698 3384 11704
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2688 11212 2740 11218
rect 2688 11154 2740 11160
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2884 10742 2912 11018
rect 2872 10736 2924 10742
rect 2872 10678 2924 10684
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2884 10062 2912 10202
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2884 9674 2912 9998
rect 2700 9646 2912 9674
rect 2700 8498 2728 9646
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3436 9110 3464 9522
rect 3424 9104 3476 9110
rect 3424 9046 3476 9052
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 3056 8492 3108 8498
rect 3056 8434 3108 8440
rect 3240 8492 3292 8498
rect 3240 8434 3292 8440
rect 3068 8090 3096 8434
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3252 7410 3280 8434
rect 3424 7880 3476 7886
rect 3424 7822 3476 7828
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 7336 3200 7342
rect 3148 7278 3200 7284
rect 3160 6798 3188 7278
rect 3252 6934 3280 7346
rect 3240 6928 3292 6934
rect 3240 6870 3292 6876
rect 3148 6792 3200 6798
rect 3148 6734 3200 6740
rect 3332 6792 3384 6798
rect 3332 6734 3384 6740
rect 3160 6610 3188 6734
rect 3160 6582 3280 6610
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3160 6322 3188 6394
rect 2780 6316 2832 6322
rect 2780 6258 2832 6264
rect 3056 6316 3108 6322
rect 3056 6258 3108 6264
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 2792 6186 2820 6258
rect 2780 6180 2832 6186
rect 2780 6122 2832 6128
rect 3068 6118 3096 6258
rect 3160 6186 3188 6258
rect 3148 6180 3200 6186
rect 3148 6122 3200 6128
rect 2688 6112 2740 6118
rect 2688 6054 2740 6060
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 2700 5778 2728 6054
rect 2688 5772 2740 5778
rect 2688 5714 2740 5720
rect 3068 5574 3096 6054
rect 3056 5568 3108 5574
rect 3056 5510 3108 5516
rect 3252 5284 3280 6582
rect 3344 6186 3372 6734
rect 3332 6180 3384 6186
rect 3332 6122 3384 6128
rect 3344 5710 3372 6122
rect 3332 5704 3384 5710
rect 3332 5646 3384 5652
rect 3160 5256 3280 5284
rect 2964 5160 3016 5166
rect 2964 5102 3016 5108
rect 2976 4282 3004 5102
rect 3160 4622 3188 5256
rect 3344 5234 3372 5646
rect 3436 5642 3464 7822
rect 3424 5636 3476 5642
rect 3424 5578 3476 5584
rect 3436 5370 3464 5578
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3332 5228 3384 5234
rect 3252 5188 3332 5216
rect 3148 4616 3200 4622
rect 3148 4558 3200 4564
rect 2964 4276 3016 4282
rect 2964 4218 3016 4224
rect 3056 4140 3108 4146
rect 3056 4082 3108 4088
rect 2780 4072 2832 4078
rect 2780 4014 2832 4020
rect 2964 4072 3016 4078
rect 2964 4014 3016 4020
rect 2792 3738 2820 4014
rect 2780 3732 2832 3738
rect 2780 3674 2832 3680
rect 2976 3398 3004 4014
rect 3068 3602 3096 4082
rect 3056 3596 3108 3602
rect 3056 3538 3108 3544
rect 3160 3534 3188 4558
rect 3252 4010 3280 5188
rect 3332 5170 3384 5176
rect 3332 4684 3384 4690
rect 3332 4626 3384 4632
rect 3240 4004 3292 4010
rect 3240 3946 3292 3952
rect 3344 3738 3372 4626
rect 3528 4298 3556 14334
rect 3606 14200 3662 14334
rect 4894 14362 4950 15000
rect 6182 14362 6238 15000
rect 7470 14362 7526 15000
rect 8758 14362 8814 15000
rect 10046 14362 10102 15000
rect 11334 14362 11390 15000
rect 12622 14362 12678 15000
rect 4894 14334 5028 14362
rect 4894 14200 4950 14334
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3700 13320 3752 13326
rect 3700 13262 3752 13268
rect 4160 13320 4212 13326
rect 4160 13262 4212 13268
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3620 11830 3648 12038
rect 3712 11898 3740 13262
rect 3884 13252 3936 13258
rect 3884 13194 3936 13200
rect 3792 13184 3844 13190
rect 3792 13126 3844 13132
rect 3804 12170 3832 13126
rect 3896 12442 3924 13194
rect 4172 12646 4200 13262
rect 4344 13184 4396 13190
rect 4344 13126 4396 13132
rect 4356 12850 4384 13126
rect 4344 12844 4396 12850
rect 4344 12786 4396 12792
rect 4620 12776 4672 12782
rect 4620 12718 4672 12724
rect 4160 12640 4212 12646
rect 4160 12582 4212 12588
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 12718
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 4620 12436 4672 12442
rect 4620 12378 4672 12384
rect 3792 12164 3844 12170
rect 3792 12106 3844 12112
rect 3700 11892 3752 11898
rect 3700 11834 3752 11840
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3804 11150 3832 12106
rect 3896 11354 3924 12378
rect 3976 12096 4028 12102
rect 3976 12038 4028 12044
rect 3988 11694 4016 12038
rect 3976 11688 4028 11694
rect 3976 11630 4028 11636
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 3896 11218 3924 11290
rect 3988 11218 4016 11630
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3976 11212 4028 11218
rect 3976 11154 4028 11160
rect 3608 11144 3660 11150
rect 3608 11086 3660 11092
rect 3792 11144 3844 11150
rect 3792 11086 3844 11092
rect 3620 10266 3648 11086
rect 3804 10810 3832 11086
rect 4528 11076 4580 11082
rect 4528 11018 4580 11024
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 4540 10742 4568 11018
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4908 10742 4936 10950
rect 4528 10736 4580 10742
rect 4528 10678 4580 10684
rect 4896 10736 4948 10742
rect 4896 10678 4948 10684
rect 4160 10600 4212 10606
rect 4080 10548 4160 10554
rect 4080 10542 4212 10548
rect 4080 10526 4200 10542
rect 4080 10266 4108 10526
rect 4908 10470 4936 10678
rect 4896 10464 4948 10470
rect 4896 10406 4948 10412
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 4068 10260 4120 10266
rect 4068 10202 4120 10208
rect 3792 10192 3844 10198
rect 3792 10134 3844 10140
rect 4804 10192 4856 10198
rect 4804 10134 4856 10140
rect 3804 10062 3832 10134
rect 3884 10124 3936 10130
rect 3884 10066 3936 10072
rect 3700 10056 3752 10062
rect 3700 9998 3752 10004
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3712 9908 3740 9998
rect 3896 9908 3924 10066
rect 4816 10062 4844 10134
rect 4804 10056 4856 10062
rect 4804 9998 4856 10004
rect 4252 9988 4304 9994
rect 4252 9930 4304 9936
rect 4620 9988 4672 9994
rect 4620 9930 4672 9936
rect 3712 9880 3924 9908
rect 4264 9586 4292 9930
rect 4252 9580 4304 9586
rect 4252 9522 4304 9528
rect 3700 9444 3752 9450
rect 3700 9386 3752 9392
rect 3712 8498 3740 9386
rect 3884 9376 3936 9382
rect 3884 9318 3936 9324
rect 3976 9376 4028 9382
rect 3976 9318 4028 9324
rect 3896 8566 3924 9318
rect 3988 9042 4016 9318
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 3884 8560 3936 8566
rect 3884 8502 3936 8508
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3620 8090 3648 8434
rect 3700 8356 3752 8362
rect 3700 8298 3752 8304
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3620 6390 3648 8026
rect 3608 6384 3660 6390
rect 3608 6326 3660 6332
rect 3608 5840 3660 5846
rect 3608 5782 3660 5788
rect 3620 5642 3648 5782
rect 3608 5636 3660 5642
rect 3608 5578 3660 5584
rect 3436 4270 3556 4298
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3436 3618 3464 4270
rect 3712 4146 3740 8298
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7478 3924 7686
rect 4172 7546 4200 7822
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3884 6860 3936 6866
rect 3884 6802 3936 6808
rect 3792 6384 3844 6390
rect 3896 6338 3924 6802
rect 3976 6724 4028 6730
rect 3976 6666 4028 6672
rect 4344 6724 4396 6730
rect 4344 6666 4396 6672
rect 3988 6458 4016 6666
rect 4068 6656 4120 6662
rect 4356 6610 4384 6666
rect 4068 6598 4120 6604
rect 3976 6452 4028 6458
rect 3976 6394 4028 6400
rect 3844 6332 3924 6338
rect 3792 6326 3924 6332
rect 3804 6310 3924 6326
rect 3896 5778 3924 6310
rect 3884 5772 3936 5778
rect 3884 5714 3936 5720
rect 3792 5636 3844 5642
rect 3792 5578 3844 5584
rect 3804 5114 3832 5578
rect 3896 5216 3924 5714
rect 3988 5692 4016 6394
rect 4080 6390 4108 6598
rect 4264 6582 4384 6610
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 4264 6118 4292 6582
rect 4252 6112 4304 6118
rect 4252 6054 4304 6060
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4068 5704 4120 5710
rect 3988 5664 4068 5692
rect 4068 5646 4120 5652
rect 4080 5302 4108 5646
rect 4068 5296 4120 5302
rect 4068 5238 4120 5244
rect 3976 5228 4028 5234
rect 3896 5188 3976 5216
rect 3976 5170 4028 5176
rect 3804 5098 3924 5114
rect 3804 5092 3936 5098
rect 3804 5086 3884 5092
rect 3884 5034 3936 5040
rect 3792 5024 3844 5030
rect 3792 4966 3844 4972
rect 3804 4690 3832 4966
rect 3896 4826 3924 5034
rect 4068 5024 4120 5030
rect 4068 4966 4120 4972
rect 3884 4820 3936 4826
rect 3884 4762 3936 4768
rect 3792 4684 3844 4690
rect 3792 4626 3844 4632
rect 3516 4140 3568 4146
rect 3516 4082 3568 4088
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3344 3590 3464 3618
rect 3148 3528 3200 3534
rect 3148 3470 3200 3476
rect 2964 3392 3016 3398
rect 2964 3334 3016 3340
rect 3160 3126 3188 3470
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 3148 3120 3200 3126
rect 3148 3062 3200 3068
rect 2792 2774 2820 3062
rect 3056 2984 3108 2990
rect 3054 2952 3056 2961
rect 3108 2952 3110 2961
rect 3054 2887 3110 2896
rect 2792 2746 2912 2774
rect 2594 2408 2650 2417
rect 2044 2372 2096 2378
rect 2594 2343 2650 2352
rect 2780 2372 2832 2378
rect 2044 2314 2096 2320
rect 2780 2314 2832 2320
rect 2056 2106 2084 2314
rect 2136 2304 2188 2310
rect 2136 2246 2188 2252
rect 2044 2100 2096 2106
rect 2044 2042 2096 2048
rect 2148 1970 2176 2246
rect 2792 2122 2820 2314
rect 2884 2122 2912 2746
rect 3344 2582 3372 3590
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3332 2576 3384 2582
rect 3332 2518 3384 2524
rect 2792 2094 2912 2122
rect 3436 2106 3464 3470
rect 3528 2854 3556 4082
rect 3608 4072 3660 4078
rect 3896 4049 3924 4082
rect 3882 4040 3938 4049
rect 3660 4020 3740 4026
rect 3608 4014 3740 4020
rect 3620 3998 3740 4014
rect 3608 3936 3660 3942
rect 3608 3878 3660 3884
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3528 2514 3556 2790
rect 3620 2514 3648 3878
rect 3712 3398 3740 3998
rect 3882 3975 3938 3984
rect 3884 3596 3936 3602
rect 3884 3538 3936 3544
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3792 3052 3844 3058
rect 3792 2994 3844 3000
rect 3516 2508 3568 2514
rect 3516 2450 3568 2456
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 2884 2038 2912 2094
rect 3424 2100 3476 2106
rect 3424 2042 3476 2048
rect 2872 2032 2924 2038
rect 3712 2009 3740 2994
rect 2872 1974 2924 1980
rect 3698 2000 3754 2009
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 2780 1896 2832 1902
rect 2780 1838 2832 1844
rect 1768 1828 1820 1834
rect 1768 1770 1820 1776
rect 940 1352 992 1358
rect 940 1294 992 1300
rect 1492 1352 1544 1358
rect 1492 1294 1544 1300
rect 952 800 980 1294
rect 1780 1018 1808 1770
rect 2424 1562 2452 1838
rect 2412 1556 2464 1562
rect 2412 1498 2464 1504
rect 1768 1012 1820 1018
rect 1768 954 1820 960
rect 2792 800 2820 1838
rect 2884 1562 2912 1974
rect 3698 1935 3754 1944
rect 2872 1556 2924 1562
rect 2872 1498 2924 1504
rect 2884 1290 2912 1498
rect 3804 1358 3832 2994
rect 3896 2854 3924 3538
rect 4080 3074 4108 4966
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4436 4480 4488 4486
rect 4436 4422 4488 4428
rect 4448 4214 4476 4422
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4528 3664 4580 3670
rect 4528 3606 4580 3612
rect 4540 3505 4568 3606
rect 4526 3496 4582 3505
rect 4632 3466 4660 9930
rect 4816 9586 4844 9998
rect 4804 9580 4856 9586
rect 4804 9522 4856 9528
rect 4712 7812 4764 7818
rect 4712 7754 4764 7760
rect 4724 7546 4752 7754
rect 5000 7562 5028 14334
rect 6182 14334 6592 14362
rect 6182 14200 6238 14334
rect 5540 13456 5592 13462
rect 5540 13398 5592 13404
rect 5552 13326 5580 13398
rect 6184 13388 6236 13394
rect 6184 13330 6236 13336
rect 5540 13320 5592 13326
rect 5540 13262 5592 13268
rect 5080 12912 5132 12918
rect 5172 12912 5224 12918
rect 5132 12872 5172 12900
rect 5080 12854 5132 12860
rect 5172 12854 5224 12860
rect 5184 11830 5212 12854
rect 5552 12345 5580 13262
rect 6092 13252 6144 13258
rect 6092 13194 6144 13200
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5538 12336 5594 12345
rect 5538 12271 5594 12280
rect 5644 12170 5672 13126
rect 6104 12986 6132 13194
rect 6092 12980 6144 12986
rect 6092 12922 6144 12928
rect 6196 12782 6224 13330
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6184 12776 6236 12782
rect 6184 12718 6236 12724
rect 6196 12306 6224 12718
rect 5908 12300 5960 12306
rect 5908 12242 5960 12248
rect 6184 12300 6236 12306
rect 6184 12242 6236 12248
rect 5448 12164 5500 12170
rect 5448 12106 5500 12112
rect 5632 12164 5684 12170
rect 5632 12106 5684 12112
rect 5460 11830 5488 12106
rect 5172 11824 5224 11830
rect 5172 11766 5224 11772
rect 5448 11824 5500 11830
rect 5448 11766 5500 11772
rect 5460 11354 5488 11766
rect 5816 11756 5868 11762
rect 5816 11698 5868 11704
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5828 10810 5856 11698
rect 5920 11014 5948 12242
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6288 11898 6316 12174
rect 6276 11892 6328 11898
rect 6276 11834 6328 11840
rect 6276 11756 6328 11762
rect 6276 11698 6328 11704
rect 5908 11008 5960 11014
rect 5908 10950 5960 10956
rect 5816 10804 5868 10810
rect 5816 10746 5868 10752
rect 5920 10674 5948 10950
rect 5908 10668 5960 10674
rect 5908 10610 5960 10616
rect 5816 10600 5868 10606
rect 6288 10588 6316 11698
rect 6380 11626 6408 12786
rect 6564 12434 6592 14334
rect 7470 14334 7880 14362
rect 7470 14200 7526 14334
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12918 6776 13262
rect 7012 13252 7064 13258
rect 7012 13194 7064 13200
rect 7564 13252 7616 13258
rect 7564 13194 7616 13200
rect 6736 12912 6788 12918
rect 7024 12866 7052 13194
rect 7196 12980 7248 12986
rect 7196 12922 7248 12928
rect 7208 12866 7236 12922
rect 6736 12854 6788 12860
rect 6932 12850 7236 12866
rect 6920 12844 7236 12850
rect 6972 12838 7236 12844
rect 6920 12786 6972 12792
rect 7472 12776 7524 12782
rect 7472 12718 7524 12724
rect 6736 12436 6788 12442
rect 6564 12406 6684 12434
rect 6552 12164 6604 12170
rect 6552 12106 6604 12112
rect 6368 11620 6420 11626
rect 6368 11562 6420 11568
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6472 11218 6500 11562
rect 6564 11354 6592 12106
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6656 11234 6684 12406
rect 6736 12378 6788 12384
rect 6748 12102 6776 12378
rect 6736 12096 6788 12102
rect 6736 12038 6788 12044
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6748 11762 6776 12038
rect 6840 11830 6868 12038
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 6920 11620 6972 11626
rect 6920 11562 6972 11568
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6564 11206 6684 11234
rect 6932 11218 6960 11562
rect 6920 11212 6972 11218
rect 6460 10600 6512 10606
rect 6288 10560 6460 10588
rect 5816 10542 5868 10548
rect 6460 10542 6512 10548
rect 5828 10130 5856 10542
rect 6276 10464 6328 10470
rect 6276 10406 6328 10412
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5920 9994 5948 10066
rect 5908 9988 5960 9994
rect 5908 9930 5960 9936
rect 5446 9888 5502 9897
rect 5446 9823 5502 9832
rect 5460 9586 5488 9823
rect 5920 9602 5948 9930
rect 5828 9586 5948 9602
rect 6012 9586 6040 10202
rect 6288 9994 6316 10406
rect 6276 9988 6328 9994
rect 6276 9930 6328 9936
rect 6288 9722 6316 9930
rect 6564 9738 6592 11206
rect 6920 11154 6972 11160
rect 6932 10266 6960 11154
rect 6920 10260 6972 10266
rect 6920 10202 6972 10208
rect 6644 9920 6696 9926
rect 7024 9897 7052 11698
rect 7116 9926 7144 11698
rect 7484 11626 7512 12718
rect 7472 11620 7524 11626
rect 7472 11562 7524 11568
rect 7576 11014 7604 13194
rect 7656 12640 7708 12646
rect 7656 12582 7708 12588
rect 7668 11762 7696 12582
rect 7852 12434 7880 14334
rect 8758 14334 9168 14362
rect 8758 14200 8814 14334
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8214 13084 8522 13093
rect 8214 13082 8220 13084
rect 8276 13082 8300 13084
rect 8356 13082 8380 13084
rect 8436 13082 8460 13084
rect 8516 13082 8522 13084
rect 8276 13030 8278 13082
rect 8458 13030 8460 13082
rect 8214 13028 8220 13030
rect 8276 13028 8300 13030
rect 8356 13028 8380 13030
rect 8436 13028 8460 13030
rect 8516 13028 8522 13030
rect 8214 13019 8522 13028
rect 7852 12406 7972 12434
rect 7656 11756 7708 11762
rect 7656 11698 7708 11704
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7838 10568 7894 10577
rect 7838 10503 7894 10512
rect 7852 10062 7880 10503
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7104 9920 7156 9926
rect 6644 9862 6696 9868
rect 7010 9888 7066 9897
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6472 9710 6592 9738
rect 5448 9580 5500 9586
rect 5448 9522 5500 9528
rect 5816 9580 5948 9586
rect 5868 9574 5948 9580
rect 6000 9580 6052 9586
rect 5816 9522 5868 9528
rect 6000 9522 6052 9528
rect 5460 8634 5488 9522
rect 6012 9178 6040 9522
rect 6472 9466 6500 9710
rect 6656 9654 6684 9862
rect 7104 9862 7156 9868
rect 7010 9823 7066 9832
rect 6644 9648 6696 9654
rect 6644 9590 6696 9596
rect 6472 9438 6592 9466
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6472 9081 6500 9114
rect 6458 9072 6514 9081
rect 6458 9007 6514 9016
rect 6472 8974 6500 9007
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 5540 8900 5592 8906
rect 5540 8842 5592 8848
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5552 8566 5580 8842
rect 5540 8560 5592 8566
rect 5540 8502 5592 8508
rect 6368 8424 6420 8430
rect 6368 8366 6420 8372
rect 5816 7880 5868 7886
rect 5816 7822 5868 7828
rect 4712 7540 4764 7546
rect 5000 7534 5120 7562
rect 4712 7482 4764 7488
rect 4712 5636 4764 5642
rect 4712 5578 4764 5584
rect 4724 5302 4752 5578
rect 4712 5296 4764 5302
rect 4712 5238 4764 5244
rect 4710 4720 4766 4729
rect 4710 4655 4766 4664
rect 4724 4486 4752 4655
rect 4712 4480 4764 4486
rect 4712 4422 4764 4428
rect 4724 3602 4752 4422
rect 4802 3904 4858 3913
rect 4802 3839 4858 3848
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4816 3534 4844 3839
rect 4804 3528 4856 3534
rect 4804 3470 4856 3476
rect 4526 3431 4582 3440
rect 4620 3460 4672 3466
rect 4620 3402 4672 3408
rect 3988 3058 4108 3074
rect 3988 3052 4120 3058
rect 3988 3046 4068 3052
rect 3884 2848 3936 2854
rect 3884 2790 3936 2796
rect 3988 2106 4016 3046
rect 4068 2994 4120 3000
rect 4160 2984 4212 2990
rect 4080 2932 4160 2938
rect 4080 2926 4212 2932
rect 4080 2910 4200 2926
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 4080 1970 4108 2910
rect 4632 2854 4660 3402
rect 4712 3120 4764 3126
rect 4712 3062 4764 3068
rect 4620 2848 4672 2854
rect 4620 2790 4672 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 4528 2644 4580 2650
rect 4528 2586 4580 2592
rect 4540 2394 4568 2586
rect 4632 2530 4660 2790
rect 4724 2650 4752 3062
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 4632 2502 4752 2530
rect 4540 2378 4660 2394
rect 4540 2372 4672 2378
rect 4540 2366 4620 2372
rect 4620 2314 4672 2320
rect 4632 2038 4660 2314
rect 4620 2032 4672 2038
rect 4620 1974 4672 1980
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 4068 1964 4120 1970
rect 4068 1906 4120 1912
rect 3988 1494 4016 1906
rect 4160 1896 4212 1902
rect 4080 1844 4160 1850
rect 4080 1838 4212 1844
rect 4620 1896 4672 1902
rect 4620 1838 4672 1844
rect 4080 1822 4200 1838
rect 3976 1488 4028 1494
rect 3976 1430 4028 1436
rect 3988 1358 4016 1430
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 3976 1352 4028 1358
rect 3976 1294 4028 1300
rect 4080 1290 4108 1822
rect 4214 1660 4522 1669
rect 4214 1658 4220 1660
rect 4276 1658 4300 1660
rect 4356 1658 4380 1660
rect 4436 1658 4460 1660
rect 4516 1658 4522 1660
rect 4276 1606 4278 1658
rect 4458 1606 4460 1658
rect 4214 1604 4220 1606
rect 4276 1604 4300 1606
rect 4356 1604 4380 1606
rect 4436 1604 4460 1606
rect 4516 1604 4522 1606
rect 4214 1595 4522 1604
rect 4632 1562 4660 1838
rect 4620 1556 4672 1562
rect 4620 1498 4672 1504
rect 4724 1442 4752 2502
rect 5092 1601 5120 7534
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5736 6730 5764 7346
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5632 6724 5684 6730
rect 5632 6666 5684 6672
rect 5724 6724 5776 6730
rect 5724 6666 5776 6672
rect 5552 6458 5580 6666
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5460 5914 5488 6122
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5552 5778 5580 6394
rect 5644 6390 5672 6666
rect 5632 6384 5684 6390
rect 5632 6326 5684 6332
rect 5724 6316 5776 6322
rect 5828 6304 5856 7822
rect 6380 7478 6408 8366
rect 6460 7880 6512 7886
rect 6460 7822 6512 7828
rect 6472 7546 6500 7822
rect 6460 7540 6512 7546
rect 6460 7482 6512 7488
rect 6368 7472 6420 7478
rect 6564 7426 6592 9438
rect 6368 7414 6420 7420
rect 6472 7398 6592 7426
rect 6182 6624 6238 6633
rect 6182 6559 6238 6568
rect 5776 6276 5856 6304
rect 5724 6258 5776 6264
rect 5736 5846 5764 6258
rect 5724 5840 5776 5846
rect 6196 5817 6224 6559
rect 5724 5782 5776 5788
rect 6182 5808 6238 5817
rect 5540 5772 5592 5778
rect 5540 5714 5592 5720
rect 5552 4690 5580 5714
rect 5736 5234 5764 5782
rect 6182 5743 6238 5752
rect 6196 5710 6224 5743
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 5724 5228 5776 5234
rect 5724 5170 5776 5176
rect 6000 4820 6052 4826
rect 6000 4762 6052 4768
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5908 4616 5960 4622
rect 5908 4558 5960 4564
rect 5816 4480 5868 4486
rect 5816 4422 5868 4428
rect 5540 4208 5592 4214
rect 5540 4150 5592 4156
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 3466 5304 3878
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 5448 3392 5500 3398
rect 5448 3334 5500 3340
rect 5460 3074 5488 3334
rect 5552 3210 5580 4150
rect 5828 3602 5856 4422
rect 5920 4049 5948 4558
rect 6012 4146 6040 4762
rect 6288 4690 6316 5510
rect 6368 5024 6420 5030
rect 6368 4966 6420 4972
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6000 4140 6052 4146
rect 6000 4082 6052 4088
rect 5906 4040 5962 4049
rect 5906 3975 5962 3984
rect 5816 3596 5868 3602
rect 5816 3538 5868 3544
rect 5632 3392 5684 3398
rect 5684 3340 5764 3346
rect 5632 3334 5764 3340
rect 5644 3318 5764 3334
rect 5552 3182 5672 3210
rect 5460 3046 5580 3074
rect 5552 2310 5580 3046
rect 5540 2304 5592 2310
rect 5540 2246 5592 2252
rect 5078 1592 5134 1601
rect 5644 1562 5672 3182
rect 5736 2650 5764 3318
rect 5814 2952 5870 2961
rect 5814 2887 5870 2896
rect 5724 2644 5776 2650
rect 5724 2586 5776 2592
rect 5736 2446 5764 2586
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5078 1527 5134 1536
rect 5632 1556 5684 1562
rect 5632 1498 5684 1504
rect 4632 1414 4752 1442
rect 2872 1284 2924 1290
rect 2872 1226 2924 1232
rect 4068 1284 4120 1290
rect 4068 1226 4120 1232
rect 4632 800 4660 1414
rect 5724 1352 5776 1358
rect 5724 1294 5776 1300
rect 5736 1018 5764 1294
rect 5828 1222 5856 2887
rect 5920 1970 5948 3975
rect 6092 2304 6144 2310
rect 6092 2246 6144 2252
rect 5998 2000 6054 2009
rect 5908 1964 5960 1970
rect 5998 1935 6054 1944
rect 5908 1906 5960 1912
rect 6012 1902 6040 1935
rect 6000 1896 6052 1902
rect 6000 1838 6052 1844
rect 6012 1358 6040 1838
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 5816 1216 5868 1222
rect 5816 1158 5868 1164
rect 5920 1170 5948 1294
rect 6104 1170 6132 2246
rect 6380 1873 6408 4966
rect 6472 4706 6500 7398
rect 6552 6248 6604 6254
rect 6552 6190 6604 6196
rect 6564 5914 6592 6190
rect 6552 5908 6604 5914
rect 6552 5850 6604 5856
rect 6564 5642 6592 5850
rect 6552 5636 6604 5642
rect 6552 5578 6604 5584
rect 6564 5370 6592 5578
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6656 4826 6684 9590
rect 7208 9518 7236 9998
rect 7668 9518 7696 9998
rect 7852 9897 7880 9998
rect 7838 9888 7894 9897
rect 7838 9823 7894 9832
rect 7196 9512 7248 9518
rect 7196 9454 7248 9460
rect 7656 9512 7708 9518
rect 7656 9454 7708 9460
rect 6828 9376 6880 9382
rect 6828 9318 6880 9324
rect 6840 8974 6868 9318
rect 7668 9042 7696 9454
rect 7656 9036 7708 9042
rect 7656 8978 7708 8984
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6736 8424 6788 8430
rect 6736 8366 6788 8372
rect 6748 7546 6776 8366
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6736 7540 6788 7546
rect 6736 7482 6788 7488
rect 7024 7449 7052 8230
rect 7010 7440 7066 7449
rect 7010 7375 7012 7384
rect 7064 7375 7066 7384
rect 7656 7404 7708 7410
rect 7012 7346 7064 7352
rect 7656 7346 7708 7352
rect 7472 7200 7524 7206
rect 7472 7142 7524 7148
rect 7484 7002 7512 7142
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 6920 6792 6972 6798
rect 6920 6734 6972 6740
rect 6736 6452 6788 6458
rect 6736 6394 6788 6400
rect 6748 6304 6776 6394
rect 6828 6316 6880 6322
rect 6748 6276 6828 6304
rect 6748 5642 6776 6276
rect 6828 6258 6880 6264
rect 6932 6254 6960 6734
rect 7208 6322 7236 6870
rect 7196 6316 7248 6322
rect 7024 6276 7196 6304
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6932 5846 6960 6190
rect 6920 5840 6972 5846
rect 6920 5782 6972 5788
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6920 5568 6972 5574
rect 7024 5556 7052 6276
rect 7196 6258 7248 6264
rect 7104 6112 7156 6118
rect 7104 6054 7156 6060
rect 7116 5710 7144 6054
rect 7668 5914 7696 7346
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7760 6390 7788 6598
rect 7748 6384 7800 6390
rect 7748 6326 7800 6332
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7380 5840 7432 5846
rect 7378 5808 7380 5817
rect 7432 5808 7434 5817
rect 7378 5743 7434 5752
rect 7104 5704 7156 5710
rect 7104 5646 7156 5652
rect 7564 5704 7616 5710
rect 7564 5646 7616 5652
rect 6972 5528 7052 5556
rect 7104 5568 7156 5574
rect 6920 5510 6972 5516
rect 7104 5510 7156 5516
rect 7116 5234 7144 5510
rect 7576 5370 7604 5646
rect 7564 5364 7616 5370
rect 7564 5306 7616 5312
rect 7104 5228 7156 5234
rect 7104 5170 7156 5176
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 6736 5024 6788 5030
rect 6736 4966 6788 4972
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 6472 4678 6684 4706
rect 6552 3596 6604 3602
rect 6552 3538 6604 3544
rect 6460 2984 6512 2990
rect 6460 2926 6512 2932
rect 6472 2106 6500 2926
rect 6460 2100 6512 2106
rect 6460 2042 6512 2048
rect 6564 2038 6592 3538
rect 6656 2106 6684 4678
rect 6748 4214 6776 4966
rect 7760 4758 7788 5102
rect 7748 4752 7800 4758
rect 7748 4694 7800 4700
rect 6828 4548 6880 4554
rect 6828 4490 6880 4496
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6736 4072 6788 4078
rect 6736 4014 6788 4020
rect 6748 3738 6776 4014
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6734 3496 6790 3505
rect 6840 3466 6868 4490
rect 6920 3936 6972 3942
rect 6920 3878 6972 3884
rect 6734 3431 6790 3440
rect 6828 3460 6880 3466
rect 6748 3210 6776 3431
rect 6828 3402 6880 3408
rect 6748 3194 6868 3210
rect 6748 3188 6880 3194
rect 6748 3182 6828 3188
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6552 2032 6604 2038
rect 6552 1974 6604 1980
rect 6748 1970 6776 3182
rect 6828 3130 6880 3136
rect 6828 2372 6880 2378
rect 6828 2314 6880 2320
rect 6736 1964 6788 1970
rect 6736 1906 6788 1912
rect 6840 1873 6868 2314
rect 6366 1864 6422 1873
rect 6366 1799 6422 1808
rect 6642 1864 6698 1873
rect 6826 1864 6882 1873
rect 6642 1799 6698 1808
rect 6736 1828 6788 1834
rect 6368 1420 6420 1426
rect 6368 1362 6420 1368
rect 6380 1272 6408 1362
rect 6656 1358 6684 1799
rect 6932 1834 6960 3878
rect 7944 2774 7972 12406
rect 8116 12164 8168 12170
rect 8116 12106 8168 12112
rect 8024 11824 8076 11830
rect 8024 11766 8076 11772
rect 8128 11778 8156 12106
rect 8214 11996 8522 12005
rect 8214 11994 8220 11996
rect 8276 11994 8300 11996
rect 8356 11994 8380 11996
rect 8436 11994 8460 11996
rect 8516 11994 8522 11996
rect 8276 11942 8278 11994
rect 8458 11942 8460 11994
rect 8214 11940 8220 11942
rect 8276 11940 8300 11942
rect 8356 11940 8380 11942
rect 8436 11940 8460 11942
rect 8516 11940 8522 11942
rect 8214 11931 8522 11940
rect 8208 11824 8260 11830
rect 8128 11772 8208 11778
rect 8128 11766 8260 11772
rect 8036 11676 8064 11766
rect 8128 11750 8248 11766
rect 8588 11694 8616 13126
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 8576 11688 8628 11694
rect 8036 11648 8156 11676
rect 8024 11552 8076 11558
rect 8024 11494 8076 11500
rect 8036 10198 8064 11494
rect 8128 10470 8156 11648
rect 8576 11630 8628 11636
rect 8680 11354 8708 12038
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 8852 11076 8904 11082
rect 8852 11018 8904 11024
rect 8668 11008 8720 11014
rect 8668 10950 8720 10956
rect 8214 10908 8522 10917
rect 8214 10906 8220 10908
rect 8276 10906 8300 10908
rect 8356 10906 8380 10908
rect 8436 10906 8460 10908
rect 8516 10906 8522 10908
rect 8276 10854 8278 10906
rect 8458 10854 8460 10906
rect 8214 10852 8220 10854
rect 8276 10852 8300 10854
rect 8356 10852 8380 10854
rect 8436 10852 8460 10854
rect 8516 10852 8522 10854
rect 8214 10843 8522 10852
rect 8680 10606 8708 10950
rect 8864 10742 8892 11018
rect 9036 11008 9088 11014
rect 9036 10950 9088 10956
rect 9048 10810 9076 10950
rect 9036 10804 9088 10810
rect 9036 10746 9088 10752
rect 8852 10736 8904 10742
rect 8852 10678 8904 10684
rect 8668 10600 8720 10606
rect 8668 10542 8720 10548
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8024 10192 8076 10198
rect 8024 10134 8076 10140
rect 8128 10062 8156 10406
rect 8576 10192 8628 10198
rect 8576 10134 8628 10140
rect 8116 10056 8168 10062
rect 8116 9998 8168 10004
rect 8214 9820 8522 9829
rect 8214 9818 8220 9820
rect 8276 9818 8300 9820
rect 8356 9818 8380 9820
rect 8436 9818 8460 9820
rect 8516 9818 8522 9820
rect 8276 9766 8278 9818
rect 8458 9766 8460 9818
rect 8214 9764 8220 9766
rect 8276 9764 8300 9766
rect 8356 9764 8380 9766
rect 8436 9764 8460 9766
rect 8516 9764 8522 9766
rect 8214 9755 8522 9764
rect 8588 9704 8616 10134
rect 8760 9988 8812 9994
rect 8760 9930 8812 9936
rect 8496 9676 8616 9704
rect 8496 9586 8524 9676
rect 8772 9654 8800 9930
rect 8760 9648 8812 9654
rect 8760 9590 8812 9596
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 8864 8838 8892 10678
rect 8944 8968 8996 8974
rect 8944 8910 8996 8916
rect 8852 8832 8904 8838
rect 8852 8774 8904 8780
rect 8214 8732 8522 8741
rect 8214 8730 8220 8732
rect 8276 8730 8300 8732
rect 8356 8730 8380 8732
rect 8436 8730 8460 8732
rect 8516 8730 8522 8732
rect 8276 8678 8278 8730
rect 8458 8678 8460 8730
rect 8214 8676 8220 8678
rect 8276 8676 8300 8678
rect 8356 8676 8380 8678
rect 8436 8676 8460 8678
rect 8516 8676 8522 8678
rect 8214 8667 8522 8676
rect 8956 8498 8984 8910
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8116 8288 8168 8294
rect 8116 8230 8168 8236
rect 8128 7954 8156 8230
rect 8312 8090 8340 8366
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 8300 8084 8352 8090
rect 8300 8026 8352 8032
rect 8116 7948 8168 7954
rect 8116 7890 8168 7896
rect 8312 7834 8340 8026
rect 8128 7806 8340 7834
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8036 7410 8064 7686
rect 8128 7478 8156 7806
rect 8214 7644 8522 7653
rect 8214 7642 8220 7644
rect 8276 7642 8300 7644
rect 8356 7642 8380 7644
rect 8436 7642 8460 7644
rect 8516 7642 8522 7644
rect 8276 7590 8278 7642
rect 8458 7590 8460 7642
rect 8214 7588 8220 7590
rect 8276 7588 8300 7590
rect 8356 7588 8380 7590
rect 8436 7588 8460 7590
rect 8516 7588 8522 7590
rect 8214 7579 8522 7588
rect 8772 7478 8800 8230
rect 8116 7472 8168 7478
rect 8116 7414 8168 7420
rect 8760 7472 8812 7478
rect 8760 7414 8812 7420
rect 8024 7404 8076 7410
rect 8024 7346 8076 7352
rect 8036 7274 8064 7346
rect 8024 7268 8076 7274
rect 8024 7210 8076 7216
rect 8214 6556 8522 6565
rect 8214 6554 8220 6556
rect 8276 6554 8300 6556
rect 8356 6554 8380 6556
rect 8436 6554 8460 6556
rect 8516 6554 8522 6556
rect 8276 6502 8278 6554
rect 8458 6502 8460 6554
rect 8214 6500 8220 6502
rect 8276 6500 8300 6502
rect 8356 6500 8380 6502
rect 8436 6500 8460 6502
rect 8516 6500 8522 6502
rect 8214 6491 8522 6500
rect 8760 6316 8812 6322
rect 8760 6258 8812 6264
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8214 5468 8522 5477
rect 8214 5466 8220 5468
rect 8276 5466 8300 5468
rect 8356 5466 8380 5468
rect 8436 5466 8460 5468
rect 8516 5466 8522 5468
rect 8276 5414 8278 5466
rect 8458 5414 8460 5466
rect 8214 5412 8220 5414
rect 8276 5412 8300 5414
rect 8356 5412 8380 5414
rect 8436 5412 8460 5414
rect 8516 5412 8522 5414
rect 8214 5403 8522 5412
rect 8116 4616 8168 4622
rect 8116 4558 8168 4564
rect 8128 4162 8156 4558
rect 8214 4380 8522 4389
rect 8214 4378 8220 4380
rect 8276 4378 8300 4380
rect 8356 4378 8380 4380
rect 8436 4378 8460 4380
rect 8516 4378 8522 4380
rect 8276 4326 8278 4378
rect 8458 4326 8460 4378
rect 8214 4324 8220 4326
rect 8276 4324 8300 4326
rect 8356 4324 8380 4326
rect 8436 4324 8460 4326
rect 8516 4324 8522 4326
rect 8214 4315 8522 4324
rect 8588 4162 8616 5646
rect 8668 5568 8720 5574
rect 8668 5510 8720 5516
rect 8128 4134 8340 4162
rect 8404 4146 8616 4162
rect 8116 3936 8168 3942
rect 8312 3913 8340 4134
rect 8392 4140 8616 4146
rect 8444 4134 8616 4140
rect 8392 4082 8444 4088
rect 8680 4078 8708 5510
rect 8772 5302 8800 6258
rect 8852 5636 8904 5642
rect 8852 5578 8904 5584
rect 8864 5370 8892 5578
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8760 5296 8812 5302
rect 8760 5238 8812 5244
rect 9048 5234 9076 5510
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 8760 4548 8812 4554
rect 8760 4490 8812 4496
rect 8772 4078 8800 4490
rect 8852 4480 8904 4486
rect 8852 4422 8904 4428
rect 8668 4072 8720 4078
rect 8668 4014 8720 4020
rect 8760 4072 8812 4078
rect 8760 4014 8812 4020
rect 8772 3942 8800 4014
rect 8760 3936 8812 3942
rect 8116 3878 8168 3884
rect 8298 3904 8354 3913
rect 8128 2990 8156 3878
rect 8760 3878 8812 3884
rect 8298 3839 8354 3848
rect 8576 3596 8628 3602
rect 8576 3538 8628 3544
rect 8214 3292 8522 3301
rect 8214 3290 8220 3292
rect 8276 3290 8300 3292
rect 8356 3290 8380 3292
rect 8436 3290 8460 3292
rect 8516 3290 8522 3292
rect 8276 3238 8278 3290
rect 8458 3238 8460 3290
rect 8214 3236 8220 3238
rect 8276 3236 8300 3238
rect 8356 3236 8380 3238
rect 8436 3236 8460 3238
rect 8516 3236 8522 3238
rect 8214 3227 8522 3236
rect 8588 3194 8616 3538
rect 8668 3460 8720 3466
rect 8668 3402 8720 3408
rect 8576 3188 8628 3194
rect 8576 3130 8628 3136
rect 8300 3120 8352 3126
rect 8300 3062 8352 3068
rect 8116 2984 8168 2990
rect 8116 2926 8168 2932
rect 7944 2746 8064 2774
rect 8036 2009 8064 2746
rect 8312 2446 8340 3062
rect 8588 2514 8616 3130
rect 8680 3126 8708 3402
rect 8864 3398 8892 4422
rect 9036 3732 9088 3738
rect 9036 3674 9088 3680
rect 8942 3632 8998 3641
rect 8942 3567 8998 3576
rect 8956 3534 8984 3567
rect 9048 3534 9076 3674
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 8852 3392 8904 3398
rect 8852 3334 8904 3340
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8668 3120 8720 3126
rect 8668 3062 8720 3068
rect 8956 2922 8984 3334
rect 9140 2961 9168 14334
rect 10046 14334 10456 14362
rect 10046 14200 10102 14334
rect 10232 13456 10284 13462
rect 10232 13398 10284 13404
rect 10244 13326 10272 13398
rect 10232 13320 10284 13326
rect 10230 13288 10232 13297
rect 10284 13288 10286 13297
rect 10230 13223 10286 13232
rect 9772 13184 9824 13190
rect 9772 13126 9824 13132
rect 9404 12980 9456 12986
rect 9404 12922 9456 12928
rect 9680 12980 9732 12986
rect 9680 12922 9732 12928
rect 9416 11694 9444 12922
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9508 12170 9536 12854
rect 9692 12434 9720 12922
rect 9784 12918 9812 13126
rect 9772 12912 9824 12918
rect 9772 12854 9824 12860
rect 9692 12406 9812 12434
rect 9784 12306 9812 12406
rect 9772 12300 9824 12306
rect 9772 12242 9824 12248
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9404 11144 9456 11150
rect 9508 11132 9536 12106
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9456 11104 9536 11132
rect 9404 11086 9456 11092
rect 9416 9722 9444 11086
rect 9600 11014 9628 11698
rect 9680 11552 9732 11558
rect 9680 11494 9732 11500
rect 9588 11008 9640 11014
rect 9588 10950 9640 10956
rect 9600 10690 9628 10950
rect 9692 10810 9720 11494
rect 9680 10804 9732 10810
rect 9680 10746 9732 10752
rect 9600 10674 9720 10690
rect 9600 10668 9732 10674
rect 9600 10662 9680 10668
rect 9600 10577 9628 10662
rect 9680 10610 9732 10616
rect 9586 10568 9642 10577
rect 9586 10503 9642 10512
rect 9784 10248 9812 12242
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 10336 10742 10364 11766
rect 9956 10736 10008 10742
rect 10324 10736 10376 10742
rect 10008 10696 10324 10724
rect 9956 10678 10008 10684
rect 10324 10678 10376 10684
rect 9784 10220 9904 10248
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9496 9988 9548 9994
rect 9496 9930 9548 9936
rect 9404 9716 9456 9722
rect 9404 9658 9456 9664
rect 9508 8498 9536 9930
rect 9784 9518 9812 10066
rect 9876 9602 9904 10220
rect 10232 9988 10284 9994
rect 10232 9930 10284 9936
rect 10244 9654 10272 9930
rect 10232 9648 10284 9654
rect 9876 9586 10088 9602
rect 10232 9590 10284 9596
rect 9876 9580 10100 9586
rect 9876 9574 10048 9580
rect 9772 9512 9824 9518
rect 9772 9454 9824 9460
rect 9784 8566 9812 9454
rect 9876 8634 9904 9574
rect 10048 9522 10100 9528
rect 10244 9518 10272 9590
rect 10232 9512 10284 9518
rect 10232 9454 10284 9460
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9772 8560 9824 8566
rect 9772 8502 9824 8508
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10152 7546 10180 7686
rect 10140 7540 10192 7546
rect 10140 7482 10192 7488
rect 9220 7472 9272 7478
rect 9220 7414 9272 7420
rect 10048 7472 10100 7478
rect 10048 7414 10100 7420
rect 9232 5556 9260 7414
rect 9496 7336 9548 7342
rect 9496 7278 9548 7284
rect 9508 7206 9536 7278
rect 9496 7200 9548 7206
rect 9496 7142 9548 7148
rect 9508 7002 9536 7142
rect 9404 6996 9456 7002
rect 9404 6938 9456 6944
rect 9496 6996 9548 7002
rect 9496 6938 9548 6944
rect 9416 6882 9444 6938
rect 9416 6854 9536 6882
rect 9508 6798 9536 6854
rect 10060 6798 10088 7414
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 9324 6458 9352 6734
rect 9772 6724 9824 6730
rect 9772 6666 9824 6672
rect 9784 6610 9812 6666
rect 9784 6582 9904 6610
rect 9312 6452 9364 6458
rect 9312 6394 9364 6400
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9312 5568 9364 5574
rect 9232 5528 9312 5556
rect 9312 5510 9364 5516
rect 9324 5030 9352 5510
rect 9692 5370 9720 6054
rect 9784 5914 9812 6190
rect 9876 6100 9904 6582
rect 10060 6458 10088 6734
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 10048 6112 10100 6118
rect 9876 6072 10048 6100
rect 10048 6054 10100 6060
rect 9772 5908 9824 5914
rect 9772 5850 9824 5856
rect 10060 5778 10088 6054
rect 10152 5846 10180 7346
rect 10140 5840 10192 5846
rect 10140 5782 10192 5788
rect 10048 5772 10100 5778
rect 10048 5714 10100 5720
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9956 5296 10008 5302
rect 9956 5238 10008 5244
rect 9312 5024 9364 5030
rect 9312 4966 9364 4972
rect 9220 4616 9272 4622
rect 9220 4558 9272 4564
rect 9126 2952 9182 2961
rect 8944 2916 8996 2922
rect 9126 2887 9182 2896
rect 8944 2858 8996 2864
rect 9232 2854 9260 4558
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 8576 2508 8628 2514
rect 8576 2450 8628 2456
rect 8300 2440 8352 2446
rect 8300 2382 8352 2388
rect 8214 2204 8522 2213
rect 8214 2202 8220 2204
rect 8276 2202 8300 2204
rect 8356 2202 8380 2204
rect 8436 2202 8460 2204
rect 8516 2202 8522 2204
rect 8276 2150 8278 2202
rect 8458 2150 8460 2202
rect 8214 2148 8220 2150
rect 8276 2148 8300 2150
rect 8356 2148 8380 2150
rect 8436 2148 8460 2150
rect 8516 2148 8522 2150
rect 8214 2139 8522 2148
rect 8300 2032 8352 2038
rect 8022 2000 8078 2009
rect 8300 1974 8352 1980
rect 8022 1935 8078 1944
rect 7840 1896 7892 1902
rect 7840 1838 7892 1844
rect 6826 1799 6882 1808
rect 6920 1828 6972 1834
rect 6736 1770 6788 1776
rect 6920 1770 6972 1776
rect 6748 1426 6776 1770
rect 7852 1562 7880 1838
rect 8312 1562 8340 1974
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 8300 1556 8352 1562
rect 8300 1498 8352 1504
rect 6736 1420 6788 1426
rect 6736 1362 6788 1368
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 8312 1290 8340 1498
rect 8300 1284 8352 1290
rect 6380 1244 6500 1272
rect 5920 1142 6132 1170
rect 5724 1012 5776 1018
rect 5724 954 5776 960
rect 6472 800 6500 1244
rect 8300 1226 8352 1232
rect 8214 1116 8522 1125
rect 8214 1114 8220 1116
rect 8276 1114 8300 1116
rect 8356 1114 8380 1116
rect 8436 1114 8460 1116
rect 8516 1114 8522 1116
rect 8276 1062 8278 1114
rect 8458 1062 8460 1114
rect 8214 1060 8220 1062
rect 8276 1060 8300 1062
rect 8356 1060 8380 1062
rect 8436 1060 8460 1062
rect 8516 1060 8522 1062
rect 8214 1051 8522 1060
rect 8312 870 8432 898
rect 8312 800 8340 870
rect 938 0 994 800
rect 2778 0 2834 800
rect 4618 0 4674 800
rect 6458 0 6514 800
rect 8298 0 8354 800
rect 8404 762 8432 870
rect 8588 762 8616 2450
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8944 2372 8996 2378
rect 8944 2314 8996 2320
rect 8668 2304 8720 2310
rect 8668 2246 8720 2252
rect 8680 1562 8708 2246
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 8956 1426 8984 2314
rect 9048 1426 9076 2382
rect 9324 1873 9352 4966
rect 9588 4616 9640 4622
rect 9588 4558 9640 4564
rect 9494 3904 9550 3913
rect 9494 3839 9550 3848
rect 9508 3738 9536 3839
rect 9496 3732 9548 3738
rect 9496 3674 9548 3680
rect 9600 3194 9628 4558
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9692 3466 9720 4422
rect 9968 4214 9996 5238
rect 10048 5160 10100 5166
rect 10048 5102 10100 5108
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10060 4282 10088 5102
rect 10152 4622 10180 5102
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 10048 4276 10100 4282
rect 10048 4218 10100 4224
rect 9956 4208 10008 4214
rect 9956 4150 10008 4156
rect 9680 3460 9732 3466
rect 9680 3402 9732 3408
rect 9968 3398 9996 4150
rect 10048 4004 10100 4010
rect 10048 3946 10100 3952
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 9588 3188 9640 3194
rect 9588 3130 9640 3136
rect 9968 3126 9996 3334
rect 9956 3120 10008 3126
rect 9956 3062 10008 3068
rect 9968 2774 9996 3062
rect 9876 2746 9996 2774
rect 9772 2576 9824 2582
rect 9772 2518 9824 2524
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9416 2106 9444 2382
rect 9496 2304 9548 2310
rect 9496 2246 9548 2252
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9508 1902 9536 2246
rect 9496 1896 9548 1902
rect 9310 1864 9366 1873
rect 9496 1838 9548 1844
rect 9310 1799 9366 1808
rect 8944 1420 8996 1426
rect 8944 1362 8996 1368
rect 9036 1420 9088 1426
rect 9036 1362 9088 1368
rect 9784 1290 9812 2518
rect 9876 1494 9904 2746
rect 10060 2582 10088 3946
rect 10152 2650 10180 4558
rect 10428 4078 10456 14334
rect 11334 14334 11468 14362
rect 11334 14200 11390 14334
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10508 13184 10560 13190
rect 10508 13126 10560 13132
rect 10520 12306 10548 13126
rect 10704 12442 10732 13194
rect 11164 12782 11192 13262
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10692 12436 10744 12442
rect 10692 12378 10744 12384
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10876 12232 10928 12238
rect 10876 12174 10928 12180
rect 10888 11898 10916 12174
rect 10876 11892 10928 11898
rect 10876 11834 10928 11840
rect 11244 11892 11296 11898
rect 11244 11834 11296 11840
rect 10508 11756 10560 11762
rect 10508 11698 10560 11704
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 11060 11756 11112 11762
rect 11060 11698 11112 11704
rect 10520 10810 10548 11698
rect 10796 11626 10824 11698
rect 10784 11620 10836 11626
rect 10784 11562 10836 11568
rect 10876 11620 10928 11626
rect 10876 11562 10928 11568
rect 10600 11008 10652 11014
rect 10600 10950 10652 10956
rect 10508 10804 10560 10810
rect 10508 10746 10560 10752
rect 10612 10674 10640 10950
rect 10796 10674 10824 11562
rect 10888 11218 10916 11562
rect 10876 11212 10928 11218
rect 10876 11154 10928 11160
rect 10968 11076 11020 11082
rect 10968 11018 11020 11024
rect 10600 10668 10652 10674
rect 10600 10610 10652 10616
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10508 10056 10560 10062
rect 10508 9998 10560 10004
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10520 9382 10548 9998
rect 10784 9988 10836 9994
rect 10784 9930 10836 9936
rect 10796 9586 10824 9930
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10784 9580 10836 9586
rect 10784 9522 10836 9528
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10612 9217 10640 9522
rect 10888 9466 10916 9998
rect 10980 9518 11008 11018
rect 11072 11014 11100 11698
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 11218 11192 11494
rect 11256 11218 11284 11834
rect 11152 11212 11204 11218
rect 11152 11154 11204 11160
rect 11244 11212 11296 11218
rect 11244 11154 11296 11160
rect 11060 11008 11112 11014
rect 11060 10950 11112 10956
rect 11336 11008 11388 11014
rect 11336 10950 11388 10956
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 11072 10674 11100 10746
rect 11348 10674 11376 10950
rect 11060 10668 11112 10674
rect 11060 10610 11112 10616
rect 11336 10668 11388 10674
rect 11336 10610 11388 10616
rect 11348 10266 11376 10610
rect 11336 10260 11388 10266
rect 11336 10202 11388 10208
rect 10704 9438 10916 9466
rect 10968 9512 11020 9518
rect 10968 9454 11020 9460
rect 10598 9208 10654 9217
rect 10598 9143 10654 9152
rect 10704 8838 10732 9438
rect 10980 8974 11008 9454
rect 11060 9444 11112 9450
rect 11060 9386 11112 9392
rect 11072 8974 11100 9386
rect 11152 9376 11204 9382
rect 11152 9318 11204 9324
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 10968 8968 11020 8974
rect 10968 8910 11020 8916
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10692 8832 10744 8838
rect 10692 8774 10744 8780
rect 10704 8634 10732 8774
rect 10692 8628 10744 8634
rect 10692 8570 10744 8576
rect 11164 8090 11192 9318
rect 11348 9042 11376 9318
rect 11336 9036 11388 9042
rect 11336 8978 11388 8984
rect 11152 8084 11204 8090
rect 11152 8026 11204 8032
rect 11440 7970 11468 14334
rect 12622 14334 12848 14362
rect 12622 14200 12678 14334
rect 12214 13628 12522 13637
rect 12214 13626 12220 13628
rect 12276 13626 12300 13628
rect 12356 13626 12380 13628
rect 12436 13626 12460 13628
rect 12516 13626 12522 13628
rect 12276 13574 12278 13626
rect 12458 13574 12460 13626
rect 12214 13572 12220 13574
rect 12276 13572 12300 13574
rect 12356 13572 12380 13574
rect 12436 13572 12460 13574
rect 12516 13572 12522 13574
rect 12214 13563 12522 13572
rect 11704 13320 11756 13326
rect 11704 13262 11756 13268
rect 11716 13190 11744 13262
rect 11980 13252 12032 13258
rect 11980 13194 12032 13200
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11704 13184 11756 13190
rect 11704 13126 11756 13132
rect 11532 12850 11560 13126
rect 11520 12844 11572 12850
rect 11520 12786 11572 12792
rect 11992 12434 12020 13194
rect 12214 12540 12522 12549
rect 12214 12538 12220 12540
rect 12276 12538 12300 12540
rect 12356 12538 12380 12540
rect 12436 12538 12460 12540
rect 12516 12538 12522 12540
rect 12276 12486 12278 12538
rect 12458 12486 12460 12538
rect 12214 12484 12220 12486
rect 12276 12484 12300 12486
rect 12356 12484 12380 12486
rect 12436 12484 12460 12486
rect 12516 12484 12522 12486
rect 12214 12475 12522 12484
rect 11992 12406 12112 12434
rect 11888 12300 11940 12306
rect 11888 12242 11940 12248
rect 11612 11756 11664 11762
rect 11612 11698 11664 11704
rect 11624 10713 11652 11698
rect 11610 10704 11666 10713
rect 11610 10639 11666 10648
rect 11704 10668 11756 10674
rect 11704 10610 11756 10616
rect 11796 10668 11848 10674
rect 11796 10610 11848 10616
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 10130 11560 10406
rect 11612 10260 11664 10266
rect 11612 10202 11664 10208
rect 11520 10124 11572 10130
rect 11520 10066 11572 10072
rect 11624 9586 11652 10202
rect 11716 9586 11744 10610
rect 11808 9586 11836 10610
rect 11900 10470 11928 12242
rect 12084 11830 12112 12406
rect 12624 12164 12676 12170
rect 12624 12106 12676 12112
rect 12072 11824 12124 11830
rect 12072 11766 12124 11772
rect 12084 11218 12112 11766
rect 12214 11452 12522 11461
rect 12214 11450 12220 11452
rect 12276 11450 12300 11452
rect 12356 11450 12380 11452
rect 12436 11450 12460 11452
rect 12516 11450 12522 11452
rect 12276 11398 12278 11450
rect 12458 11398 12460 11450
rect 12214 11396 12220 11398
rect 12276 11396 12300 11398
rect 12356 11396 12380 11398
rect 12436 11396 12460 11398
rect 12516 11396 12522 11398
rect 12214 11387 12522 11396
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12636 11150 12664 12106
rect 12716 11688 12768 11694
rect 12716 11630 12768 11636
rect 12728 11354 12756 11630
rect 12716 11348 12768 11354
rect 12716 11290 12768 11296
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 11888 10464 11940 10470
rect 11888 10406 11940 10412
rect 11992 9586 12020 10610
rect 12214 10364 12522 10373
rect 12214 10362 12220 10364
rect 12276 10362 12300 10364
rect 12356 10362 12380 10364
rect 12436 10362 12460 10364
rect 12516 10362 12522 10364
rect 12276 10310 12278 10362
rect 12458 10310 12460 10362
rect 12214 10308 12220 10310
rect 12276 10308 12300 10310
rect 12356 10308 12380 10310
rect 12436 10308 12460 10310
rect 12516 10308 12522 10310
rect 12214 10299 12522 10308
rect 12072 9648 12124 9654
rect 12072 9590 12124 9596
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11796 9580 11848 9586
rect 11796 9522 11848 9528
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11702 9208 11758 9217
rect 11612 9172 11664 9178
rect 11702 9143 11704 9152
rect 11612 9114 11664 9120
rect 11756 9143 11758 9152
rect 11704 9114 11756 9120
rect 11624 8786 11652 9114
rect 11704 8832 11756 8838
rect 11624 8780 11704 8786
rect 11624 8774 11756 8780
rect 11624 8758 11744 8774
rect 11624 8430 11652 8758
rect 11612 8424 11664 8430
rect 11612 8366 11664 8372
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 10784 7948 10836 7954
rect 10784 7890 10836 7896
rect 11348 7942 11468 7970
rect 11716 7954 11744 8298
rect 11808 8106 11836 9522
rect 12084 8498 12112 9590
rect 12624 9512 12676 9518
rect 12624 9454 12676 9460
rect 12214 9276 12522 9285
rect 12214 9274 12220 9276
rect 12276 9274 12300 9276
rect 12356 9274 12380 9276
rect 12436 9274 12460 9276
rect 12516 9274 12522 9276
rect 12276 9222 12278 9274
rect 12458 9222 12460 9274
rect 12214 9220 12220 9222
rect 12276 9220 12300 9222
rect 12356 9220 12380 9222
rect 12436 9220 12460 9222
rect 12516 9220 12522 9222
rect 12214 9211 12522 9220
rect 12636 8634 12664 9454
rect 12820 9160 12848 14334
rect 13910 14200 13966 15000
rect 15198 14200 15254 15000
rect 16486 14362 16542 15000
rect 16040 14334 16542 14362
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 14740 13320 14792 13326
rect 14740 13262 14792 13268
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 13280 12986 13308 13262
rect 14752 12986 14780 13262
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 13268 12980 13320 12986
rect 13268 12922 13320 12928
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 13820 12912 13872 12918
rect 13820 12854 13872 12860
rect 13452 12844 13504 12850
rect 13452 12786 13504 12792
rect 13464 12442 13492 12786
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13728 12232 13780 12238
rect 13728 12174 13780 12180
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13372 10742 13400 11494
rect 13464 11150 13492 11630
rect 13556 11150 13584 11698
rect 13740 11354 13768 12174
rect 13728 11348 13780 11354
rect 13728 11290 13780 11296
rect 13452 11144 13504 11150
rect 13452 11086 13504 11092
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 13464 10606 13492 11086
rect 13832 11082 13860 12854
rect 14844 12850 14872 13126
rect 15488 12986 15516 13262
rect 15568 13184 15620 13190
rect 15568 13126 15620 13132
rect 15476 12980 15528 12986
rect 15476 12922 15528 12928
rect 15580 12850 15608 13126
rect 16040 12850 16068 14334
rect 16486 14200 16542 14334
rect 17774 14362 17830 15000
rect 19062 14362 19118 15000
rect 20350 14362 20406 15000
rect 17774 14334 17908 14362
rect 17774 14200 17830 14334
rect 16120 13320 16172 13326
rect 16120 13262 16172 13268
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 16132 12986 16160 13262
rect 16214 13084 16522 13093
rect 16214 13082 16220 13084
rect 16276 13082 16300 13084
rect 16356 13082 16380 13084
rect 16436 13082 16460 13084
rect 16516 13082 16522 13084
rect 16276 13030 16278 13082
rect 16458 13030 16460 13082
rect 16214 13028 16220 13030
rect 16276 13028 16300 13030
rect 16356 13028 16380 13030
rect 16436 13028 16460 13030
rect 16516 13028 16522 13030
rect 16214 13019 16522 13028
rect 16120 12980 16172 12986
rect 16120 12922 16172 12928
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 15568 12844 15620 12850
rect 15568 12786 15620 12792
rect 16028 12844 16080 12850
rect 16028 12786 16080 12792
rect 16592 12442 16620 13262
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16764 13184 16816 13190
rect 16764 13126 16816 13132
rect 16684 12918 16712 13126
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16580 12436 16632 12442
rect 16580 12378 16632 12384
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 14372 12164 14424 12170
rect 14372 12106 14424 12112
rect 14384 11898 14412 12106
rect 14740 12096 14792 12102
rect 14740 12038 14792 12044
rect 14372 11892 14424 11898
rect 14372 11834 14424 11840
rect 13820 11076 13872 11082
rect 13820 11018 13872 11024
rect 13832 10742 13860 11018
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13452 10600 13504 10606
rect 13452 10542 13504 10548
rect 12992 10464 13044 10470
rect 12992 10406 13044 10412
rect 12820 9132 12940 9160
rect 12808 9036 12860 9042
rect 12808 8978 12860 8984
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12072 8492 12124 8498
rect 12072 8434 12124 8440
rect 12820 8430 12848 8978
rect 12808 8424 12860 8430
rect 12808 8366 12860 8372
rect 12214 8188 12522 8197
rect 12214 8186 12220 8188
rect 12276 8186 12300 8188
rect 12356 8186 12380 8188
rect 12436 8186 12460 8188
rect 12516 8186 12522 8188
rect 12276 8134 12278 8186
rect 12458 8134 12460 8186
rect 12214 8132 12220 8134
rect 12276 8132 12300 8134
rect 12356 8132 12380 8134
rect 12436 8132 12460 8134
rect 12516 8132 12522 8134
rect 12214 8123 12522 8132
rect 11808 8078 11928 8106
rect 12912 8090 12940 9132
rect 13004 8498 13032 10406
rect 13464 10266 13492 10542
rect 13452 10260 13504 10266
rect 13452 10202 13504 10208
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 13268 9988 13320 9994
rect 13268 9930 13320 9936
rect 13544 9988 13596 9994
rect 13544 9930 13596 9936
rect 13096 9722 13124 9930
rect 13176 9920 13228 9926
rect 13176 9862 13228 9868
rect 13188 9722 13216 9862
rect 13084 9716 13136 9722
rect 13084 9658 13136 9664
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13084 9512 13136 9518
rect 13084 9454 13136 9460
rect 13096 9110 13124 9454
rect 13084 9104 13136 9110
rect 13084 9046 13136 9052
rect 13096 8634 13124 9046
rect 13280 8974 13308 9930
rect 13556 9654 13584 9930
rect 13544 9648 13596 9654
rect 13832 9636 13860 10678
rect 13912 10464 13964 10470
rect 13912 10406 13964 10412
rect 13924 10062 13952 10406
rect 13912 10056 13964 10062
rect 13910 10024 13912 10033
rect 13964 10024 13966 10033
rect 13910 9959 13966 9968
rect 13912 9648 13964 9654
rect 13832 9608 13912 9636
rect 13544 9590 13596 9596
rect 13912 9590 13964 9596
rect 13820 9512 13872 9518
rect 13820 9454 13872 9460
rect 13832 9178 13860 9454
rect 13820 9172 13872 9178
rect 13872 9132 13952 9160
rect 13820 9114 13872 9120
rect 13268 8968 13320 8974
rect 13268 8910 13320 8916
rect 13544 8968 13596 8974
rect 13544 8910 13596 8916
rect 13268 8832 13320 8838
rect 13268 8774 13320 8780
rect 13084 8628 13136 8634
rect 13084 8570 13136 8576
rect 13280 8566 13308 8774
rect 13556 8566 13584 8910
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13544 8560 13596 8566
rect 13544 8502 13596 8508
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13360 8288 13412 8294
rect 13360 8230 13412 8236
rect 11704 7948 11756 7954
rect 10692 7268 10744 7274
rect 10692 7210 10744 7216
rect 10704 5642 10732 7210
rect 10796 6322 10824 7890
rect 11060 7404 11112 7410
rect 11060 7346 11112 7352
rect 11072 6662 11100 7346
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11060 6656 11112 6662
rect 11060 6598 11112 6604
rect 10784 6316 10836 6322
rect 10784 6258 10836 6264
rect 10692 5636 10744 5642
rect 10692 5578 10744 5584
rect 10796 5302 10824 6258
rect 11072 5778 11100 6598
rect 11164 6322 11192 7142
rect 11244 6656 11296 6662
rect 11244 6598 11296 6604
rect 11256 6390 11284 6598
rect 11244 6384 11296 6390
rect 11244 6326 11296 6332
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11348 5778 11376 7942
rect 11704 7890 11756 7896
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11440 7546 11468 7822
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11428 6996 11480 7002
rect 11428 6938 11480 6944
rect 11440 6458 11468 6938
rect 11796 6724 11848 6730
rect 11796 6666 11848 6672
rect 11428 6452 11480 6458
rect 11428 6394 11480 6400
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11336 5772 11388 5778
rect 11336 5714 11388 5720
rect 11704 5772 11756 5778
rect 11704 5714 11756 5720
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10796 4570 10824 5238
rect 11716 5098 11744 5714
rect 11808 5710 11836 6666
rect 11796 5704 11848 5710
rect 11796 5646 11848 5652
rect 11704 5092 11756 5098
rect 11704 5034 11756 5040
rect 11612 5024 11664 5030
rect 11612 4966 11664 4972
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11624 4690 11652 4966
rect 11612 4684 11664 4690
rect 11612 4626 11664 4632
rect 10796 4554 10916 4570
rect 10796 4548 10928 4554
rect 10796 4542 10876 4548
rect 10796 4214 10824 4542
rect 10876 4490 10928 4496
rect 10784 4208 10836 4214
rect 10784 4150 10836 4156
rect 10416 4072 10468 4078
rect 10416 4014 10468 4020
rect 10416 3936 10468 3942
rect 10416 3878 10468 3884
rect 10428 3126 10456 3878
rect 10796 3466 10824 4150
rect 11808 4146 11836 4966
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 10968 4004 11020 4010
rect 10968 3946 11020 3952
rect 10980 3670 11008 3946
rect 10968 3664 11020 3670
rect 10968 3606 11020 3612
rect 10784 3460 10836 3466
rect 10784 3402 10836 3408
rect 10416 3120 10468 3126
rect 10416 3062 10468 3068
rect 10508 2984 10560 2990
rect 10508 2926 10560 2932
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 10048 2576 10100 2582
rect 10048 2518 10100 2524
rect 10322 2544 10378 2553
rect 10322 2479 10378 2488
rect 10336 2446 10364 2479
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 10140 1760 10192 1766
rect 10140 1702 10192 1708
rect 9864 1488 9916 1494
rect 9864 1430 9916 1436
rect 9772 1284 9824 1290
rect 9772 1226 9824 1232
rect 10152 800 10180 1702
rect 10428 1222 10456 2790
rect 10520 1902 10548 2926
rect 10796 2774 10824 3402
rect 10980 3058 11008 3606
rect 11900 3602 11928 8078
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12912 7342 12940 8026
rect 13372 7954 13400 8230
rect 13360 7948 13412 7954
rect 13360 7890 13412 7896
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13464 7342 13492 7482
rect 12900 7336 12952 7342
rect 12900 7278 12952 7284
rect 13452 7336 13504 7342
rect 13452 7278 13504 7284
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12214 7100 12522 7109
rect 12214 7098 12220 7100
rect 12276 7098 12300 7100
rect 12356 7098 12380 7100
rect 12436 7098 12460 7100
rect 12516 7098 12522 7100
rect 12276 7046 12278 7098
rect 12458 7046 12460 7098
rect 12214 7044 12220 7046
rect 12276 7044 12300 7046
rect 12356 7044 12380 7046
rect 12436 7044 12460 7046
rect 12516 7044 12522 7046
rect 12214 7035 12522 7044
rect 12912 7002 12940 7142
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13372 6390 13400 6666
rect 13360 6384 13412 6390
rect 13360 6326 13412 6332
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 11992 5914 12020 6190
rect 12214 6012 12522 6021
rect 12214 6010 12220 6012
rect 12276 6010 12300 6012
rect 12356 6010 12380 6012
rect 12436 6010 12460 6012
rect 12516 6010 12522 6012
rect 12276 5958 12278 6010
rect 12458 5958 12460 6010
rect 12214 5956 12220 5958
rect 12276 5956 12300 5958
rect 12356 5956 12380 5958
rect 12436 5956 12460 5958
rect 12516 5956 12522 5958
rect 12214 5947 12522 5956
rect 11980 5908 12032 5914
rect 11980 5850 12032 5856
rect 12532 5704 12584 5710
rect 12716 5704 12768 5710
rect 12532 5646 12584 5652
rect 12636 5652 12716 5658
rect 12636 5646 12768 5652
rect 12544 5302 12572 5646
rect 12636 5630 12756 5646
rect 12532 5296 12584 5302
rect 12532 5238 12584 5244
rect 12636 5234 12664 5630
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 12624 5228 12676 5234
rect 12624 5170 12676 5176
rect 12214 4924 12522 4933
rect 12214 4922 12220 4924
rect 12276 4922 12300 4924
rect 12356 4922 12380 4924
rect 12436 4922 12460 4924
rect 12516 4922 12522 4924
rect 12276 4870 12278 4922
rect 12458 4870 12460 4922
rect 12214 4868 12220 4870
rect 12276 4868 12300 4870
rect 12356 4868 12380 4870
rect 12436 4868 12460 4870
rect 12516 4868 12522 4870
rect 12214 4859 12522 4868
rect 12636 4706 12664 5170
rect 12728 4826 12756 5510
rect 13096 5234 13124 5510
rect 13084 5228 13136 5234
rect 13084 5170 13136 5176
rect 13464 5030 13492 7278
rect 13556 5914 13584 8502
rect 13728 7744 13780 7750
rect 13728 7686 13780 7692
rect 13740 7478 13768 7686
rect 13728 7472 13780 7478
rect 13728 7414 13780 7420
rect 13820 7336 13872 7342
rect 13820 7278 13872 7284
rect 13832 6866 13860 7278
rect 13820 6860 13872 6866
rect 13820 6802 13872 6808
rect 13544 5908 13596 5914
rect 13544 5850 13596 5856
rect 13544 5296 13596 5302
rect 13544 5238 13596 5244
rect 13452 5024 13504 5030
rect 13452 4966 13504 4972
rect 12716 4820 12768 4826
rect 12716 4762 12768 4768
rect 12636 4690 12756 4706
rect 12636 4684 12768 4690
rect 12636 4678 12716 4684
rect 12716 4626 12768 4632
rect 13360 4684 13412 4690
rect 13360 4626 13412 4632
rect 13084 4548 13136 4554
rect 13084 4490 13136 4496
rect 12072 4480 12124 4486
rect 12072 4422 12124 4428
rect 12084 4214 12112 4422
rect 12072 4208 12124 4214
rect 12072 4150 12124 4156
rect 13096 4146 13124 4490
rect 13084 4140 13136 4146
rect 13084 4082 13136 4088
rect 13268 4072 13320 4078
rect 13268 4014 13320 4020
rect 12214 3836 12522 3845
rect 12214 3834 12220 3836
rect 12276 3834 12300 3836
rect 12356 3834 12380 3836
rect 12436 3834 12460 3836
rect 12516 3834 12522 3836
rect 12276 3782 12278 3834
rect 12458 3782 12460 3834
rect 12214 3780 12220 3782
rect 12276 3780 12300 3782
rect 12356 3780 12380 3782
rect 12436 3780 12460 3782
rect 12516 3780 12522 3782
rect 12214 3771 12522 3780
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 13084 3460 13136 3466
rect 13280 3448 13308 4014
rect 13136 3420 13308 3448
rect 13084 3402 13136 3408
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 10796 2746 11008 2774
rect 10980 2378 11008 2746
rect 11072 2514 11100 2858
rect 11060 2508 11112 2514
rect 11060 2450 11112 2456
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 10600 2304 10652 2310
rect 10652 2252 10824 2258
rect 10600 2246 10824 2252
rect 10612 2230 10824 2246
rect 10796 1902 10824 2230
rect 10508 1896 10560 1902
rect 10784 1896 10836 1902
rect 10508 1838 10560 1844
rect 10782 1864 10784 1873
rect 10836 1864 10838 1873
rect 10782 1799 10838 1808
rect 10980 1290 11008 2314
rect 11060 2304 11112 2310
rect 11060 2246 11112 2252
rect 11072 1426 11100 2246
rect 11532 2106 11560 2994
rect 11992 2854 12020 3402
rect 13280 3058 13308 3420
rect 13268 3052 13320 3058
rect 13268 2994 13320 3000
rect 12624 2984 12676 2990
rect 12624 2926 12676 2932
rect 11980 2848 12032 2854
rect 11980 2790 12032 2796
rect 12214 2748 12522 2757
rect 12214 2746 12220 2748
rect 12276 2746 12300 2748
rect 12356 2746 12380 2748
rect 12436 2746 12460 2748
rect 12516 2746 12522 2748
rect 12276 2694 12278 2746
rect 12458 2694 12460 2746
rect 12214 2692 12220 2694
rect 12276 2692 12300 2694
rect 12356 2692 12380 2694
rect 12436 2692 12460 2694
rect 12516 2692 12522 2694
rect 12214 2683 12522 2692
rect 12636 2650 12664 2926
rect 13372 2922 13400 4626
rect 13556 4282 13584 5238
rect 13636 5160 13688 5166
rect 13636 5102 13688 5108
rect 13648 4826 13676 5102
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13924 4146 13952 9132
rect 14280 7880 14332 7886
rect 14280 7822 14332 7828
rect 14096 7744 14148 7750
rect 14096 7686 14148 7692
rect 14108 6866 14136 7686
rect 14292 7342 14320 7822
rect 14752 7392 14780 12038
rect 15764 11762 15792 12242
rect 16776 12238 16804 13126
rect 17420 12442 17448 13262
rect 17880 12918 17908 14334
rect 18892 14334 19118 14362
rect 18604 13184 18656 13190
rect 18604 13126 18656 13132
rect 18616 12918 18644 13126
rect 18892 12918 18920 14334
rect 19062 14200 19118 14334
rect 20088 14334 20406 14362
rect 19800 13184 19852 13190
rect 19800 13126 19852 13132
rect 17868 12912 17920 12918
rect 17868 12854 17920 12860
rect 18604 12912 18656 12918
rect 18604 12854 18656 12860
rect 18880 12912 18932 12918
rect 18880 12854 18932 12860
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 17408 12436 17460 12442
rect 17408 12378 17460 12384
rect 16764 12232 16816 12238
rect 16764 12174 16816 12180
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 16214 11996 16522 12005
rect 16214 11994 16220 11996
rect 16276 11994 16300 11996
rect 16356 11994 16380 11996
rect 16436 11994 16460 11996
rect 16516 11994 16522 11996
rect 16276 11942 16278 11994
rect 16458 11942 16460 11994
rect 16214 11940 16220 11942
rect 16276 11940 16300 11942
rect 16356 11940 16380 11942
rect 16436 11940 16460 11942
rect 16516 11940 16522 11942
rect 16214 11931 16522 11940
rect 18340 11898 18368 12174
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 18892 11762 18920 12038
rect 19628 11898 19656 12786
rect 19812 12238 19840 13126
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 19996 12238 20024 12854
rect 20088 12306 20116 14334
rect 20350 14200 20406 14334
rect 21638 14362 21694 15000
rect 22926 14362 22982 15000
rect 21638 14334 21772 14362
rect 21638 14200 21694 14334
rect 20214 13628 20522 13637
rect 20214 13626 20220 13628
rect 20276 13626 20300 13628
rect 20356 13626 20380 13628
rect 20436 13626 20460 13628
rect 20516 13626 20522 13628
rect 20276 13574 20278 13626
rect 20458 13574 20460 13626
rect 20214 13572 20220 13574
rect 20276 13572 20300 13574
rect 20356 13572 20380 13574
rect 20436 13572 20460 13574
rect 20516 13572 20522 13574
rect 20214 13563 20522 13572
rect 21744 13258 21772 14334
rect 22664 14334 22982 14362
rect 21824 13320 21876 13326
rect 21824 13262 21876 13268
rect 20628 13252 20680 13258
rect 20628 13194 20680 13200
rect 21732 13252 21784 13258
rect 21732 13194 21784 13200
rect 20214 12540 20522 12549
rect 20214 12538 20220 12540
rect 20276 12538 20300 12540
rect 20356 12538 20380 12540
rect 20436 12538 20460 12540
rect 20516 12538 20522 12540
rect 20276 12486 20278 12538
rect 20458 12486 20460 12538
rect 20214 12484 20220 12486
rect 20276 12484 20300 12486
rect 20356 12484 20380 12486
rect 20436 12484 20460 12486
rect 20516 12484 20522 12486
rect 20214 12475 20522 12484
rect 20640 12306 20668 13194
rect 20812 12776 20864 12782
rect 20812 12718 20864 12724
rect 20076 12300 20128 12306
rect 20076 12242 20128 12248
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 19800 12232 19852 12238
rect 19800 12174 19852 12180
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19616 11892 19668 11898
rect 19616 11834 19668 11840
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 18880 11756 18932 11762
rect 18880 11698 18932 11704
rect 16028 11620 16080 11626
rect 16028 11562 16080 11568
rect 15384 11552 15436 11558
rect 15384 11494 15436 11500
rect 15396 11218 15424 11494
rect 15384 11212 15436 11218
rect 15384 11154 15436 11160
rect 16040 11150 16068 11562
rect 16684 11354 16712 11698
rect 16672 11348 16724 11354
rect 16672 11290 16724 11296
rect 16028 11144 16080 11150
rect 16028 11086 16080 11092
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15016 11008 15068 11014
rect 15016 10950 15068 10956
rect 15028 9994 15056 10950
rect 15764 10810 15792 11018
rect 16214 10908 16522 10917
rect 16214 10906 16220 10908
rect 16276 10906 16300 10908
rect 16356 10906 16380 10908
rect 16436 10906 16460 10908
rect 16516 10906 16522 10908
rect 16276 10854 16278 10906
rect 16458 10854 16460 10906
rect 16214 10852 16220 10854
rect 16276 10852 16300 10854
rect 16356 10852 16380 10854
rect 16436 10852 16460 10854
rect 16516 10852 16522 10854
rect 16214 10843 16522 10852
rect 15752 10804 15804 10810
rect 15752 10746 15804 10752
rect 15936 10736 15988 10742
rect 15936 10678 15988 10684
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15660 10668 15712 10674
rect 15660 10610 15712 10616
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 10130 15148 10406
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 14832 9988 14884 9994
rect 14832 9930 14884 9936
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 14844 9518 14872 9930
rect 14832 9512 14884 9518
rect 14832 9454 14884 9460
rect 15028 9450 15056 9930
rect 15304 9722 15332 10610
rect 15672 10266 15700 10610
rect 15752 10600 15804 10606
rect 15752 10542 15804 10548
rect 15764 10266 15792 10542
rect 15660 10260 15712 10266
rect 15660 10202 15712 10208
rect 15752 10260 15804 10266
rect 15752 10202 15804 10208
rect 15948 10062 15976 10678
rect 17960 10600 18012 10606
rect 17960 10542 18012 10548
rect 16580 10532 16632 10538
rect 16580 10474 16632 10480
rect 16488 10464 16540 10470
rect 16488 10406 16540 10412
rect 16500 10130 16528 10406
rect 16488 10124 16540 10130
rect 16488 10066 16540 10072
rect 15936 10056 15988 10062
rect 15936 9998 15988 10004
rect 15476 9920 15528 9926
rect 15476 9862 15528 9868
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 9586 15332 9658
rect 15488 9654 15516 9862
rect 15476 9648 15528 9654
rect 15476 9590 15528 9596
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 15568 9444 15620 9450
rect 15568 9386 15620 9392
rect 15028 9178 15056 9386
rect 15016 9172 15068 9178
rect 15016 9114 15068 9120
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 15476 8968 15528 8974
rect 15476 8910 15528 8916
rect 14936 7954 14964 8910
rect 15200 8832 15252 8838
rect 15200 8774 15252 8780
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 15212 7834 15240 8774
rect 15488 8634 15516 8910
rect 15580 8906 15608 9386
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15856 8906 15884 9318
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15476 8628 15528 8634
rect 15476 8570 15528 8576
rect 15948 8362 15976 9998
rect 16592 9994 16620 10474
rect 17972 10266 18000 10542
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 16580 9988 16632 9994
rect 16580 9930 16632 9936
rect 16214 9820 16522 9829
rect 16214 9818 16220 9820
rect 16276 9818 16300 9820
rect 16356 9818 16380 9820
rect 16436 9818 16460 9820
rect 16516 9818 16522 9820
rect 16276 9766 16278 9818
rect 16458 9766 16460 9818
rect 16214 9764 16220 9766
rect 16276 9764 16300 9766
rect 16356 9764 16380 9766
rect 16436 9764 16460 9766
rect 16516 9764 16522 9766
rect 16214 9755 16522 9764
rect 16592 9654 16620 9930
rect 16580 9648 16632 9654
rect 16408 9608 16580 9636
rect 16028 9376 16080 9382
rect 16028 9318 16080 9324
rect 16040 8566 16068 9318
rect 16408 9178 16436 9608
rect 16580 9590 16632 9596
rect 17408 9648 17460 9654
rect 17408 9590 17460 9596
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16408 8906 16436 9114
rect 16500 8922 16528 9454
rect 16948 9444 17000 9450
rect 16948 9386 17000 9392
rect 16396 8900 16448 8906
rect 16500 8894 16620 8922
rect 16396 8842 16448 8848
rect 16214 8732 16522 8741
rect 16214 8730 16220 8732
rect 16276 8730 16300 8732
rect 16356 8730 16380 8732
rect 16436 8730 16460 8732
rect 16516 8730 16522 8732
rect 16276 8678 16278 8730
rect 16458 8678 16460 8730
rect 16214 8676 16220 8678
rect 16276 8676 16300 8678
rect 16356 8676 16380 8678
rect 16436 8676 16460 8678
rect 16516 8676 16522 8678
rect 16214 8667 16522 8676
rect 16028 8560 16080 8566
rect 16592 8514 16620 8894
rect 16028 8502 16080 8508
rect 16500 8498 16620 8514
rect 16500 8492 16632 8498
rect 16500 8486 16580 8492
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 16500 8090 16528 8486
rect 16580 8434 16632 8440
rect 16960 8430 16988 9386
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17236 8566 17264 8910
rect 17420 8566 17448 9590
rect 18420 9512 18472 9518
rect 18420 9454 18472 9460
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 18432 8634 18460 9454
rect 19444 9178 19472 9454
rect 19432 9172 19484 9178
rect 19432 9114 19484 9120
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17408 8560 17460 8566
rect 17408 8502 17460 8508
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 15120 7818 15240 7834
rect 15108 7812 15240 7818
rect 15160 7806 15240 7812
rect 15292 7812 15344 7818
rect 15108 7754 15160 7760
rect 15292 7754 15344 7760
rect 15304 7410 15332 7754
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 7410 15700 7686
rect 16214 7644 16522 7653
rect 16214 7642 16220 7644
rect 16276 7642 16300 7644
rect 16356 7642 16380 7644
rect 16436 7642 16460 7644
rect 16516 7642 16522 7644
rect 16276 7590 16278 7642
rect 16458 7590 16460 7642
rect 16214 7588 16220 7590
rect 16276 7588 16300 7590
rect 16356 7588 16380 7590
rect 16436 7588 16460 7590
rect 16516 7588 16522 7590
rect 16214 7579 16522 7588
rect 14832 7404 14884 7410
rect 14752 7364 14832 7392
rect 15292 7404 15344 7410
rect 14884 7364 14964 7392
rect 14832 7346 14884 7352
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14936 6730 14964 7364
rect 15292 7346 15344 7352
rect 15384 7404 15436 7410
rect 15384 7346 15436 7352
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15396 7274 15424 7346
rect 15384 7268 15436 7274
rect 15384 7210 15436 7216
rect 15396 6934 15424 7210
rect 15384 6928 15436 6934
rect 15384 6870 15436 6876
rect 15672 6866 15700 7346
rect 19996 7274 20024 12174
rect 20824 11898 20852 12718
rect 21836 12646 21864 13262
rect 22284 13252 22336 13258
rect 22284 13194 22336 13200
rect 22100 12912 22152 12918
rect 22100 12854 22152 12860
rect 21824 12640 21876 12646
rect 21824 12582 21876 12588
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 21836 11762 21864 12582
rect 22112 12170 22140 12854
rect 22296 12306 22324 13194
rect 22664 12918 22692 14334
rect 22926 14200 22982 14334
rect 22652 12912 22704 12918
rect 22652 12854 22704 12860
rect 22284 12300 22336 12306
rect 22284 12242 22336 12248
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 21824 11756 21876 11762
rect 21824 11698 21876 11704
rect 20214 11452 20522 11461
rect 20214 11450 20220 11452
rect 20276 11450 20300 11452
rect 20356 11450 20380 11452
rect 20436 11450 20460 11452
rect 20516 11450 20522 11452
rect 20276 11398 20278 11450
rect 20458 11398 20460 11450
rect 20214 11396 20220 11398
rect 20276 11396 20300 11398
rect 20356 11396 20380 11398
rect 20436 11396 20460 11398
rect 20516 11396 20522 11398
rect 20214 11387 20522 11396
rect 20214 10364 20522 10373
rect 20214 10362 20220 10364
rect 20276 10362 20300 10364
rect 20356 10362 20380 10364
rect 20436 10362 20460 10364
rect 20516 10362 20522 10364
rect 20276 10310 20278 10362
rect 20458 10310 20460 10362
rect 20214 10308 20220 10310
rect 20276 10308 20300 10310
rect 20356 10308 20380 10310
rect 20436 10308 20460 10310
rect 20516 10308 20522 10310
rect 20214 10299 20522 10308
rect 20214 9276 20522 9285
rect 20214 9274 20220 9276
rect 20276 9274 20300 9276
rect 20356 9274 20380 9276
rect 20436 9274 20460 9276
rect 20516 9274 20522 9276
rect 20276 9222 20278 9274
rect 20458 9222 20460 9274
rect 20214 9220 20220 9222
rect 20276 9220 20300 9222
rect 20356 9220 20380 9222
rect 20436 9220 20460 9222
rect 20516 9220 20522 9222
rect 20214 9211 20522 9220
rect 20214 8188 20522 8197
rect 20214 8186 20220 8188
rect 20276 8186 20300 8188
rect 20356 8186 20380 8188
rect 20436 8186 20460 8188
rect 20516 8186 20522 8188
rect 20276 8134 20278 8186
rect 20458 8134 20460 8186
rect 20214 8132 20220 8134
rect 20276 8132 20300 8134
rect 20356 8132 20380 8134
rect 20436 8132 20460 8134
rect 20516 8132 20522 8134
rect 20214 8123 20522 8132
rect 22098 7440 22154 7449
rect 22098 7375 22154 7384
rect 22112 7342 22140 7375
rect 22100 7336 22152 7342
rect 22100 7278 22152 7284
rect 19984 7268 20036 7274
rect 19984 7210 20036 7216
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 16028 7200 16080 7206
rect 16028 7142 16080 7148
rect 15856 7002 15884 7142
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 16040 6866 16068 7142
rect 20214 7100 20522 7109
rect 20214 7098 20220 7100
rect 20276 7098 20300 7100
rect 20356 7098 20380 7100
rect 20436 7098 20460 7100
rect 20516 7098 20522 7100
rect 20276 7046 20278 7098
rect 20458 7046 20460 7098
rect 20214 7044 20220 7046
rect 20276 7044 20300 7046
rect 20356 7044 20380 7046
rect 20436 7044 20460 7046
rect 20516 7044 20522 7046
rect 20214 7035 20522 7044
rect 15660 6860 15712 6866
rect 15660 6802 15712 6808
rect 16028 6860 16080 6866
rect 16028 6802 16080 6808
rect 14924 6724 14976 6730
rect 14924 6666 14976 6672
rect 14936 6610 14964 6666
rect 15108 6656 15160 6662
rect 14936 6604 15108 6610
rect 14936 6598 15160 6604
rect 14936 6582 15148 6598
rect 14936 6390 14964 6582
rect 16214 6556 16522 6565
rect 16214 6554 16220 6556
rect 16276 6554 16300 6556
rect 16356 6554 16380 6556
rect 16436 6554 16460 6556
rect 16516 6554 16522 6556
rect 16276 6502 16278 6554
rect 16458 6502 16460 6554
rect 16214 6500 16220 6502
rect 16276 6500 16300 6502
rect 16356 6500 16380 6502
rect 16436 6500 16460 6502
rect 16516 6500 16522 6502
rect 16214 6491 16522 6500
rect 14924 6384 14976 6390
rect 14924 6326 14976 6332
rect 14936 5710 14964 6326
rect 20214 6012 20522 6021
rect 20214 6010 20220 6012
rect 20276 6010 20300 6012
rect 20356 6010 20380 6012
rect 20436 6010 20460 6012
rect 20516 6010 20522 6012
rect 20276 5958 20278 6010
rect 20458 5958 20460 6010
rect 20214 5956 20220 5958
rect 20276 5956 20300 5958
rect 20356 5956 20380 5958
rect 20436 5956 20460 5958
rect 20516 5956 20522 5958
rect 20214 5947 20522 5956
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14936 5302 14964 5646
rect 16214 5468 16522 5477
rect 16214 5466 16220 5468
rect 16276 5466 16300 5468
rect 16356 5466 16380 5468
rect 16436 5466 16460 5468
rect 16516 5466 16522 5468
rect 16276 5414 16278 5466
rect 16458 5414 16460 5466
rect 16214 5412 16220 5414
rect 16276 5412 16300 5414
rect 16356 5412 16380 5414
rect 16436 5412 16460 5414
rect 16516 5412 16522 5414
rect 16214 5403 16522 5412
rect 14924 5296 14976 5302
rect 14924 5238 14976 5244
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14096 4480 14148 4486
rect 14096 4422 14148 4428
rect 13912 4140 13964 4146
rect 13912 4082 13964 4088
rect 13544 2984 13596 2990
rect 13544 2926 13596 2932
rect 13360 2916 13412 2922
rect 13360 2858 13412 2864
rect 12348 2644 12400 2650
rect 12348 2586 12400 2592
rect 12624 2644 12676 2650
rect 12624 2586 12676 2592
rect 12716 2644 12768 2650
rect 12716 2586 12768 2592
rect 11980 2576 12032 2582
rect 11978 2544 11980 2553
rect 12360 2553 12388 2586
rect 12728 2553 12756 2586
rect 12032 2544 12034 2553
rect 11612 2508 11664 2514
rect 11978 2479 12034 2488
rect 12346 2544 12402 2553
rect 12346 2479 12402 2488
rect 12714 2544 12770 2553
rect 12714 2479 12770 2488
rect 11612 2450 11664 2456
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 11242 1592 11298 1601
rect 11242 1527 11244 1536
rect 11296 1527 11298 1536
rect 11244 1498 11296 1504
rect 11532 1426 11560 2042
rect 11624 2038 11652 2450
rect 12256 2372 12308 2378
rect 12256 2314 12308 2320
rect 11888 2304 11940 2310
rect 11888 2246 11940 2252
rect 11900 2038 11928 2246
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11888 2032 11940 2038
rect 11888 1974 11940 1980
rect 11980 2032 12032 2038
rect 11980 1974 12032 1980
rect 11060 1420 11112 1426
rect 11060 1362 11112 1368
rect 11520 1420 11572 1426
rect 11520 1362 11572 1368
rect 10968 1284 11020 1290
rect 10968 1226 11020 1232
rect 10416 1216 10468 1222
rect 10416 1158 10468 1164
rect 11992 800 12020 1974
rect 12268 1952 12296 2314
rect 12176 1924 12296 1952
rect 12624 1964 12676 1970
rect 12072 1896 12124 1902
rect 12176 1884 12204 1924
rect 12624 1906 12676 1912
rect 12124 1856 12204 1884
rect 12072 1838 12124 1844
rect 12214 1660 12522 1669
rect 12214 1658 12220 1660
rect 12276 1658 12300 1660
rect 12356 1658 12380 1660
rect 12436 1658 12460 1660
rect 12516 1658 12522 1660
rect 12276 1606 12278 1658
rect 12458 1606 12460 1658
rect 12214 1604 12220 1606
rect 12276 1604 12300 1606
rect 12356 1604 12380 1606
rect 12436 1604 12460 1606
rect 12516 1604 12522 1606
rect 12214 1595 12522 1604
rect 12636 1306 12664 1906
rect 13556 1902 13584 2926
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 13728 2508 13780 2514
rect 13728 2450 13780 2456
rect 13740 2310 13768 2450
rect 13832 2446 13860 2790
rect 13924 2650 13952 4082
rect 14108 3602 14136 4422
rect 14096 3596 14148 3602
rect 14096 3538 14148 3544
rect 14292 3466 14320 4558
rect 14936 4078 14964 5238
rect 20214 4924 20522 4933
rect 20214 4922 20220 4924
rect 20276 4922 20300 4924
rect 20356 4922 20380 4924
rect 20436 4922 20460 4924
rect 20516 4922 20522 4924
rect 20276 4870 20278 4922
rect 20458 4870 20460 4922
rect 20214 4868 20220 4870
rect 20276 4868 20300 4870
rect 20356 4868 20380 4870
rect 20436 4868 20460 4870
rect 20516 4868 20522 4870
rect 20214 4859 20522 4868
rect 16214 4380 16522 4389
rect 16214 4378 16220 4380
rect 16276 4378 16300 4380
rect 16356 4378 16380 4380
rect 16436 4378 16460 4380
rect 16516 4378 16522 4380
rect 16276 4326 16278 4378
rect 16458 4326 16460 4378
rect 16214 4324 16220 4326
rect 16276 4324 16300 4326
rect 16356 4324 16380 4326
rect 16436 4324 16460 4326
rect 16516 4324 16522 4326
rect 16214 4315 16522 4324
rect 14924 4072 14976 4078
rect 14924 4014 14976 4020
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15672 3466 15700 4014
rect 20214 3836 20522 3845
rect 20214 3834 20220 3836
rect 20276 3834 20300 3836
rect 20356 3834 20380 3836
rect 20436 3834 20460 3836
rect 20516 3834 20522 3836
rect 20276 3782 20278 3834
rect 20458 3782 20460 3834
rect 20214 3780 20220 3782
rect 20276 3780 20300 3782
rect 20356 3780 20380 3782
rect 20436 3780 20460 3782
rect 20516 3780 20522 3782
rect 20214 3771 20522 3780
rect 14280 3460 14332 3466
rect 14280 3402 14332 3408
rect 15660 3460 15712 3466
rect 15660 3402 15712 3408
rect 14292 3126 14320 3402
rect 14280 3120 14332 3126
rect 14280 3062 14332 3068
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14002 2952 14058 2961
rect 14002 2887 14058 2896
rect 14016 2650 14044 2887
rect 13912 2644 13964 2650
rect 13912 2586 13964 2592
rect 14004 2644 14056 2650
rect 14004 2586 14056 2592
rect 14188 2576 14240 2582
rect 14188 2518 14240 2524
rect 13912 2508 13964 2514
rect 13912 2450 13964 2456
rect 13820 2440 13872 2446
rect 13820 2382 13872 2388
rect 13728 2304 13780 2310
rect 13728 2246 13780 2252
rect 13544 1896 13596 1902
rect 13544 1838 13596 1844
rect 12544 1290 12664 1306
rect 12532 1284 12664 1290
rect 12584 1278 12664 1284
rect 12532 1226 12584 1232
rect 13924 1170 13952 2450
rect 14096 2440 14148 2446
rect 14094 2408 14096 2417
rect 14148 2408 14150 2417
rect 14094 2343 14150 2352
rect 14200 1970 14228 2518
rect 14936 2106 14964 2994
rect 15672 2854 15700 3402
rect 15844 3392 15896 3398
rect 15844 3334 15896 3340
rect 15856 3194 15884 3334
rect 16214 3292 16522 3301
rect 16214 3290 16220 3292
rect 16276 3290 16300 3292
rect 16356 3290 16380 3292
rect 16436 3290 16460 3292
rect 16516 3290 16522 3292
rect 16276 3238 16278 3290
rect 16458 3238 16460 3290
rect 16214 3236 16220 3238
rect 16276 3236 16300 3238
rect 16356 3236 16380 3238
rect 16436 3236 16460 3238
rect 16516 3236 16522 3238
rect 16214 3227 16522 3236
rect 15844 3188 15896 3194
rect 15844 3130 15896 3136
rect 15660 2848 15712 2854
rect 15660 2790 15712 2796
rect 22192 2848 22244 2854
rect 22192 2790 22244 2796
rect 20214 2748 20522 2757
rect 20214 2746 20220 2748
rect 20276 2746 20300 2748
rect 20356 2746 20380 2748
rect 20436 2746 20460 2748
rect 20516 2746 20522 2748
rect 20276 2694 20278 2746
rect 20458 2694 20460 2746
rect 20214 2692 20220 2694
rect 20276 2692 20300 2694
rect 20356 2692 20380 2694
rect 20436 2692 20460 2694
rect 20516 2692 20522 2694
rect 20214 2683 20522 2692
rect 22098 2544 22154 2553
rect 22098 2479 22154 2488
rect 22112 2378 22140 2479
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 15028 2106 15056 2246
rect 16214 2204 16522 2213
rect 16214 2202 16220 2204
rect 16276 2202 16300 2204
rect 16356 2202 16380 2204
rect 16436 2202 16460 2204
rect 16516 2202 16522 2204
rect 16276 2150 16278 2202
rect 16458 2150 16460 2202
rect 16214 2148 16220 2150
rect 16276 2148 16300 2150
rect 16356 2148 16380 2150
rect 16436 2148 16460 2150
rect 16516 2148 16522 2150
rect 16214 2139 16522 2148
rect 14924 2100 14976 2106
rect 14924 2042 14976 2048
rect 15016 2100 15068 2106
rect 15016 2042 15068 2048
rect 20258 2000 20314 2009
rect 14188 1964 14240 1970
rect 14188 1906 14240 1912
rect 15016 1964 15068 1970
rect 22204 1970 22232 2790
rect 23020 2372 23072 2378
rect 23020 2314 23072 2320
rect 20258 1935 20260 1944
rect 15016 1906 15068 1912
rect 20312 1935 20314 1944
rect 22192 1964 22244 1970
rect 20260 1906 20312 1912
rect 22192 1906 22244 1912
rect 14556 1896 14608 1902
rect 14556 1838 14608 1844
rect 14568 1222 14596 1838
rect 14648 1760 14700 1766
rect 14648 1702 14700 1708
rect 14660 1358 14688 1702
rect 15028 1562 15056 1906
rect 15660 1896 15712 1902
rect 15660 1838 15712 1844
rect 17500 1896 17552 1902
rect 17500 1838 17552 1844
rect 19340 1896 19392 1902
rect 19340 1838 19392 1844
rect 21180 1896 21232 1902
rect 21180 1838 21232 1844
rect 15016 1556 15068 1562
rect 15016 1498 15068 1504
rect 14648 1352 14700 1358
rect 14648 1294 14700 1300
rect 13832 1142 13952 1170
rect 14556 1216 14608 1222
rect 14556 1158 14608 1164
rect 13832 800 13860 1142
rect 15672 800 15700 1838
rect 16214 1116 16522 1125
rect 16214 1114 16220 1116
rect 16276 1114 16300 1116
rect 16356 1114 16380 1116
rect 16436 1114 16460 1116
rect 16516 1114 16522 1116
rect 16276 1062 16278 1114
rect 16458 1062 16460 1114
rect 16214 1060 16220 1062
rect 16276 1060 16300 1062
rect 16356 1060 16380 1062
rect 16436 1060 16460 1062
rect 16516 1060 16522 1062
rect 16214 1051 16522 1060
rect 17512 800 17540 1838
rect 19352 800 19380 1838
rect 20214 1660 20522 1669
rect 20214 1658 20220 1660
rect 20276 1658 20300 1660
rect 20356 1658 20380 1660
rect 20436 1658 20460 1660
rect 20516 1658 20522 1660
rect 20276 1606 20278 1658
rect 20458 1606 20460 1658
rect 20214 1604 20220 1606
rect 20276 1604 20300 1606
rect 20356 1604 20380 1606
rect 20436 1604 20460 1606
rect 20516 1604 20522 1606
rect 20214 1595 20522 1604
rect 21192 800 21220 1838
rect 23032 800 23060 2314
rect 8404 734 8616 762
rect 10138 0 10194 800
rect 11978 0 12034 800
rect 13818 0 13874 800
rect 15658 0 15714 800
rect 17498 0 17554 800
rect 19338 0 19394 800
rect 21178 0 21234 800
rect 23018 0 23074 800
<< via2 >>
rect 1766 11464 1822 11520
rect 1582 8200 1638 8256
rect 1306 5752 1362 5808
rect 2410 4120 2466 4176
rect 2410 3576 2466 3632
rect 1306 3304 1362 3360
rect 1766 2488 1822 2544
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 3054 2932 3056 2952
rect 3056 2932 3108 2952
rect 3108 2932 3110 2952
rect 3054 2896 3110 2932
rect 2594 2352 2650 2408
rect 3882 3984 3938 4040
rect 3698 1944 3754 2000
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4526 3440 4582 3496
rect 5538 12280 5594 12336
rect 5446 9832 5502 9888
rect 8220 13082 8276 13084
rect 8300 13082 8356 13084
rect 8380 13082 8436 13084
rect 8460 13082 8516 13084
rect 8220 13030 8266 13082
rect 8266 13030 8276 13082
rect 8300 13030 8330 13082
rect 8330 13030 8342 13082
rect 8342 13030 8356 13082
rect 8380 13030 8394 13082
rect 8394 13030 8406 13082
rect 8406 13030 8436 13082
rect 8460 13030 8470 13082
rect 8470 13030 8516 13082
rect 8220 13028 8276 13030
rect 8300 13028 8356 13030
rect 8380 13028 8436 13030
rect 8460 13028 8516 13030
rect 7838 10512 7894 10568
rect 7010 9832 7066 9888
rect 6458 9016 6514 9072
rect 4710 4664 4766 4720
rect 4802 3848 4858 3904
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4220 1658 4276 1660
rect 4300 1658 4356 1660
rect 4380 1658 4436 1660
rect 4460 1658 4516 1660
rect 4220 1606 4266 1658
rect 4266 1606 4276 1658
rect 4300 1606 4330 1658
rect 4330 1606 4342 1658
rect 4342 1606 4356 1658
rect 4380 1606 4394 1658
rect 4394 1606 4406 1658
rect 4406 1606 4436 1658
rect 4460 1606 4470 1658
rect 4470 1606 4516 1658
rect 4220 1604 4276 1606
rect 4300 1604 4356 1606
rect 4380 1604 4436 1606
rect 4460 1604 4516 1606
rect 6182 6568 6238 6624
rect 6182 5752 6238 5808
rect 5906 3984 5962 4040
rect 5078 1536 5134 1592
rect 5814 2896 5870 2952
rect 5998 1944 6054 2000
rect 7838 9832 7894 9888
rect 7010 7404 7066 7440
rect 7010 7384 7012 7404
rect 7012 7384 7064 7404
rect 7064 7384 7066 7404
rect 7378 5788 7380 5808
rect 7380 5788 7432 5808
rect 7432 5788 7434 5808
rect 7378 5752 7434 5788
rect 6734 3440 6790 3496
rect 6366 1808 6422 1864
rect 6642 1808 6698 1864
rect 6826 1808 6882 1864
rect 8220 11994 8276 11996
rect 8300 11994 8356 11996
rect 8380 11994 8436 11996
rect 8460 11994 8516 11996
rect 8220 11942 8266 11994
rect 8266 11942 8276 11994
rect 8300 11942 8330 11994
rect 8330 11942 8342 11994
rect 8342 11942 8356 11994
rect 8380 11942 8394 11994
rect 8394 11942 8406 11994
rect 8406 11942 8436 11994
rect 8460 11942 8470 11994
rect 8470 11942 8516 11994
rect 8220 11940 8276 11942
rect 8300 11940 8356 11942
rect 8380 11940 8436 11942
rect 8460 11940 8516 11942
rect 8220 10906 8276 10908
rect 8300 10906 8356 10908
rect 8380 10906 8436 10908
rect 8460 10906 8516 10908
rect 8220 10854 8266 10906
rect 8266 10854 8276 10906
rect 8300 10854 8330 10906
rect 8330 10854 8342 10906
rect 8342 10854 8356 10906
rect 8380 10854 8394 10906
rect 8394 10854 8406 10906
rect 8406 10854 8436 10906
rect 8460 10854 8470 10906
rect 8470 10854 8516 10906
rect 8220 10852 8276 10854
rect 8300 10852 8356 10854
rect 8380 10852 8436 10854
rect 8460 10852 8516 10854
rect 8220 9818 8276 9820
rect 8300 9818 8356 9820
rect 8380 9818 8436 9820
rect 8460 9818 8516 9820
rect 8220 9766 8266 9818
rect 8266 9766 8276 9818
rect 8300 9766 8330 9818
rect 8330 9766 8342 9818
rect 8342 9766 8356 9818
rect 8380 9766 8394 9818
rect 8394 9766 8406 9818
rect 8406 9766 8436 9818
rect 8460 9766 8470 9818
rect 8470 9766 8516 9818
rect 8220 9764 8276 9766
rect 8300 9764 8356 9766
rect 8380 9764 8436 9766
rect 8460 9764 8516 9766
rect 8220 8730 8276 8732
rect 8300 8730 8356 8732
rect 8380 8730 8436 8732
rect 8460 8730 8516 8732
rect 8220 8678 8266 8730
rect 8266 8678 8276 8730
rect 8300 8678 8330 8730
rect 8330 8678 8342 8730
rect 8342 8678 8356 8730
rect 8380 8678 8394 8730
rect 8394 8678 8406 8730
rect 8406 8678 8436 8730
rect 8460 8678 8470 8730
rect 8470 8678 8516 8730
rect 8220 8676 8276 8678
rect 8300 8676 8356 8678
rect 8380 8676 8436 8678
rect 8460 8676 8516 8678
rect 8220 7642 8276 7644
rect 8300 7642 8356 7644
rect 8380 7642 8436 7644
rect 8460 7642 8516 7644
rect 8220 7590 8266 7642
rect 8266 7590 8276 7642
rect 8300 7590 8330 7642
rect 8330 7590 8342 7642
rect 8342 7590 8356 7642
rect 8380 7590 8394 7642
rect 8394 7590 8406 7642
rect 8406 7590 8436 7642
rect 8460 7590 8470 7642
rect 8470 7590 8516 7642
rect 8220 7588 8276 7590
rect 8300 7588 8356 7590
rect 8380 7588 8436 7590
rect 8460 7588 8516 7590
rect 8220 6554 8276 6556
rect 8300 6554 8356 6556
rect 8380 6554 8436 6556
rect 8460 6554 8516 6556
rect 8220 6502 8266 6554
rect 8266 6502 8276 6554
rect 8300 6502 8330 6554
rect 8330 6502 8342 6554
rect 8342 6502 8356 6554
rect 8380 6502 8394 6554
rect 8394 6502 8406 6554
rect 8406 6502 8436 6554
rect 8460 6502 8470 6554
rect 8470 6502 8516 6554
rect 8220 6500 8276 6502
rect 8300 6500 8356 6502
rect 8380 6500 8436 6502
rect 8460 6500 8516 6502
rect 8220 5466 8276 5468
rect 8300 5466 8356 5468
rect 8380 5466 8436 5468
rect 8460 5466 8516 5468
rect 8220 5414 8266 5466
rect 8266 5414 8276 5466
rect 8300 5414 8330 5466
rect 8330 5414 8342 5466
rect 8342 5414 8356 5466
rect 8380 5414 8394 5466
rect 8394 5414 8406 5466
rect 8406 5414 8436 5466
rect 8460 5414 8470 5466
rect 8470 5414 8516 5466
rect 8220 5412 8276 5414
rect 8300 5412 8356 5414
rect 8380 5412 8436 5414
rect 8460 5412 8516 5414
rect 8220 4378 8276 4380
rect 8300 4378 8356 4380
rect 8380 4378 8436 4380
rect 8460 4378 8516 4380
rect 8220 4326 8266 4378
rect 8266 4326 8276 4378
rect 8300 4326 8330 4378
rect 8330 4326 8342 4378
rect 8342 4326 8356 4378
rect 8380 4326 8394 4378
rect 8394 4326 8406 4378
rect 8406 4326 8436 4378
rect 8460 4326 8470 4378
rect 8470 4326 8516 4378
rect 8220 4324 8276 4326
rect 8300 4324 8356 4326
rect 8380 4324 8436 4326
rect 8460 4324 8516 4326
rect 8298 3848 8354 3904
rect 8220 3290 8276 3292
rect 8300 3290 8356 3292
rect 8380 3290 8436 3292
rect 8460 3290 8516 3292
rect 8220 3238 8266 3290
rect 8266 3238 8276 3290
rect 8300 3238 8330 3290
rect 8330 3238 8342 3290
rect 8342 3238 8356 3290
rect 8380 3238 8394 3290
rect 8394 3238 8406 3290
rect 8406 3238 8436 3290
rect 8460 3238 8470 3290
rect 8470 3238 8516 3290
rect 8220 3236 8276 3238
rect 8300 3236 8356 3238
rect 8380 3236 8436 3238
rect 8460 3236 8516 3238
rect 8942 3576 8998 3632
rect 10230 13268 10232 13288
rect 10232 13268 10284 13288
rect 10284 13268 10286 13288
rect 10230 13232 10286 13268
rect 9586 10512 9642 10568
rect 9126 2896 9182 2952
rect 8220 2202 8276 2204
rect 8300 2202 8356 2204
rect 8380 2202 8436 2204
rect 8460 2202 8516 2204
rect 8220 2150 8266 2202
rect 8266 2150 8276 2202
rect 8300 2150 8330 2202
rect 8330 2150 8342 2202
rect 8342 2150 8356 2202
rect 8380 2150 8394 2202
rect 8394 2150 8406 2202
rect 8406 2150 8436 2202
rect 8460 2150 8470 2202
rect 8470 2150 8516 2202
rect 8220 2148 8276 2150
rect 8300 2148 8356 2150
rect 8380 2148 8436 2150
rect 8460 2148 8516 2150
rect 8022 1944 8078 2000
rect 8220 1114 8276 1116
rect 8300 1114 8356 1116
rect 8380 1114 8436 1116
rect 8460 1114 8516 1116
rect 8220 1062 8266 1114
rect 8266 1062 8276 1114
rect 8300 1062 8330 1114
rect 8330 1062 8342 1114
rect 8342 1062 8356 1114
rect 8380 1062 8394 1114
rect 8394 1062 8406 1114
rect 8406 1062 8436 1114
rect 8460 1062 8470 1114
rect 8470 1062 8516 1114
rect 8220 1060 8276 1062
rect 8300 1060 8356 1062
rect 8380 1060 8436 1062
rect 8460 1060 8516 1062
rect 9494 3848 9550 3904
rect 9310 1808 9366 1864
rect 10598 9152 10654 9208
rect 12220 13626 12276 13628
rect 12300 13626 12356 13628
rect 12380 13626 12436 13628
rect 12460 13626 12516 13628
rect 12220 13574 12266 13626
rect 12266 13574 12276 13626
rect 12300 13574 12330 13626
rect 12330 13574 12342 13626
rect 12342 13574 12356 13626
rect 12380 13574 12394 13626
rect 12394 13574 12406 13626
rect 12406 13574 12436 13626
rect 12460 13574 12470 13626
rect 12470 13574 12516 13626
rect 12220 13572 12276 13574
rect 12300 13572 12356 13574
rect 12380 13572 12436 13574
rect 12460 13572 12516 13574
rect 12220 12538 12276 12540
rect 12300 12538 12356 12540
rect 12380 12538 12436 12540
rect 12460 12538 12516 12540
rect 12220 12486 12266 12538
rect 12266 12486 12276 12538
rect 12300 12486 12330 12538
rect 12330 12486 12342 12538
rect 12342 12486 12356 12538
rect 12380 12486 12394 12538
rect 12394 12486 12406 12538
rect 12406 12486 12436 12538
rect 12460 12486 12470 12538
rect 12470 12486 12516 12538
rect 12220 12484 12276 12486
rect 12300 12484 12356 12486
rect 12380 12484 12436 12486
rect 12460 12484 12516 12486
rect 11610 10648 11666 10704
rect 12220 11450 12276 11452
rect 12300 11450 12356 11452
rect 12380 11450 12436 11452
rect 12460 11450 12516 11452
rect 12220 11398 12266 11450
rect 12266 11398 12276 11450
rect 12300 11398 12330 11450
rect 12330 11398 12342 11450
rect 12342 11398 12356 11450
rect 12380 11398 12394 11450
rect 12394 11398 12406 11450
rect 12406 11398 12436 11450
rect 12460 11398 12470 11450
rect 12470 11398 12516 11450
rect 12220 11396 12276 11398
rect 12300 11396 12356 11398
rect 12380 11396 12436 11398
rect 12460 11396 12516 11398
rect 12220 10362 12276 10364
rect 12300 10362 12356 10364
rect 12380 10362 12436 10364
rect 12460 10362 12516 10364
rect 12220 10310 12266 10362
rect 12266 10310 12276 10362
rect 12300 10310 12330 10362
rect 12330 10310 12342 10362
rect 12342 10310 12356 10362
rect 12380 10310 12394 10362
rect 12394 10310 12406 10362
rect 12406 10310 12436 10362
rect 12460 10310 12470 10362
rect 12470 10310 12516 10362
rect 12220 10308 12276 10310
rect 12300 10308 12356 10310
rect 12380 10308 12436 10310
rect 12460 10308 12516 10310
rect 11702 9172 11758 9208
rect 11702 9152 11704 9172
rect 11704 9152 11756 9172
rect 11756 9152 11758 9172
rect 12220 9274 12276 9276
rect 12300 9274 12356 9276
rect 12380 9274 12436 9276
rect 12460 9274 12516 9276
rect 12220 9222 12266 9274
rect 12266 9222 12276 9274
rect 12300 9222 12330 9274
rect 12330 9222 12342 9274
rect 12342 9222 12356 9274
rect 12380 9222 12394 9274
rect 12394 9222 12406 9274
rect 12406 9222 12436 9274
rect 12460 9222 12470 9274
rect 12470 9222 12516 9274
rect 12220 9220 12276 9222
rect 12300 9220 12356 9222
rect 12380 9220 12436 9222
rect 12460 9220 12516 9222
rect 16220 13082 16276 13084
rect 16300 13082 16356 13084
rect 16380 13082 16436 13084
rect 16460 13082 16516 13084
rect 16220 13030 16266 13082
rect 16266 13030 16276 13082
rect 16300 13030 16330 13082
rect 16330 13030 16342 13082
rect 16342 13030 16356 13082
rect 16380 13030 16394 13082
rect 16394 13030 16406 13082
rect 16406 13030 16436 13082
rect 16460 13030 16470 13082
rect 16470 13030 16516 13082
rect 16220 13028 16276 13030
rect 16300 13028 16356 13030
rect 16380 13028 16436 13030
rect 16460 13028 16516 13030
rect 12220 8186 12276 8188
rect 12300 8186 12356 8188
rect 12380 8186 12436 8188
rect 12460 8186 12516 8188
rect 12220 8134 12266 8186
rect 12266 8134 12276 8186
rect 12300 8134 12330 8186
rect 12330 8134 12342 8186
rect 12342 8134 12356 8186
rect 12380 8134 12394 8186
rect 12394 8134 12406 8186
rect 12406 8134 12436 8186
rect 12460 8134 12470 8186
rect 12470 8134 12516 8186
rect 12220 8132 12276 8134
rect 12300 8132 12356 8134
rect 12380 8132 12436 8134
rect 12460 8132 12516 8134
rect 13910 10004 13912 10024
rect 13912 10004 13964 10024
rect 13964 10004 13966 10024
rect 13910 9968 13966 10004
rect 10322 2488 10378 2544
rect 12220 7098 12276 7100
rect 12300 7098 12356 7100
rect 12380 7098 12436 7100
rect 12460 7098 12516 7100
rect 12220 7046 12266 7098
rect 12266 7046 12276 7098
rect 12300 7046 12330 7098
rect 12330 7046 12342 7098
rect 12342 7046 12356 7098
rect 12380 7046 12394 7098
rect 12394 7046 12406 7098
rect 12406 7046 12436 7098
rect 12460 7046 12470 7098
rect 12470 7046 12516 7098
rect 12220 7044 12276 7046
rect 12300 7044 12356 7046
rect 12380 7044 12436 7046
rect 12460 7044 12516 7046
rect 12220 6010 12276 6012
rect 12300 6010 12356 6012
rect 12380 6010 12436 6012
rect 12460 6010 12516 6012
rect 12220 5958 12266 6010
rect 12266 5958 12276 6010
rect 12300 5958 12330 6010
rect 12330 5958 12342 6010
rect 12342 5958 12356 6010
rect 12380 5958 12394 6010
rect 12394 5958 12406 6010
rect 12406 5958 12436 6010
rect 12460 5958 12470 6010
rect 12470 5958 12516 6010
rect 12220 5956 12276 5958
rect 12300 5956 12356 5958
rect 12380 5956 12436 5958
rect 12460 5956 12516 5958
rect 12220 4922 12276 4924
rect 12300 4922 12356 4924
rect 12380 4922 12436 4924
rect 12460 4922 12516 4924
rect 12220 4870 12266 4922
rect 12266 4870 12276 4922
rect 12300 4870 12330 4922
rect 12330 4870 12342 4922
rect 12342 4870 12356 4922
rect 12380 4870 12394 4922
rect 12394 4870 12406 4922
rect 12406 4870 12436 4922
rect 12460 4870 12470 4922
rect 12470 4870 12516 4922
rect 12220 4868 12276 4870
rect 12300 4868 12356 4870
rect 12380 4868 12436 4870
rect 12460 4868 12516 4870
rect 12220 3834 12276 3836
rect 12300 3834 12356 3836
rect 12380 3834 12436 3836
rect 12460 3834 12516 3836
rect 12220 3782 12266 3834
rect 12266 3782 12276 3834
rect 12300 3782 12330 3834
rect 12330 3782 12342 3834
rect 12342 3782 12356 3834
rect 12380 3782 12394 3834
rect 12394 3782 12406 3834
rect 12406 3782 12436 3834
rect 12460 3782 12470 3834
rect 12470 3782 12516 3834
rect 12220 3780 12276 3782
rect 12300 3780 12356 3782
rect 12380 3780 12436 3782
rect 12460 3780 12516 3782
rect 10782 1844 10784 1864
rect 10784 1844 10836 1864
rect 10836 1844 10838 1864
rect 10782 1808 10838 1844
rect 12220 2746 12276 2748
rect 12300 2746 12356 2748
rect 12380 2746 12436 2748
rect 12460 2746 12516 2748
rect 12220 2694 12266 2746
rect 12266 2694 12276 2746
rect 12300 2694 12330 2746
rect 12330 2694 12342 2746
rect 12342 2694 12356 2746
rect 12380 2694 12394 2746
rect 12394 2694 12406 2746
rect 12406 2694 12436 2746
rect 12460 2694 12470 2746
rect 12470 2694 12516 2746
rect 12220 2692 12276 2694
rect 12300 2692 12356 2694
rect 12380 2692 12436 2694
rect 12460 2692 12516 2694
rect 16220 11994 16276 11996
rect 16300 11994 16356 11996
rect 16380 11994 16436 11996
rect 16460 11994 16516 11996
rect 16220 11942 16266 11994
rect 16266 11942 16276 11994
rect 16300 11942 16330 11994
rect 16330 11942 16342 11994
rect 16342 11942 16356 11994
rect 16380 11942 16394 11994
rect 16394 11942 16406 11994
rect 16406 11942 16436 11994
rect 16460 11942 16470 11994
rect 16470 11942 16516 11994
rect 16220 11940 16276 11942
rect 16300 11940 16356 11942
rect 16380 11940 16436 11942
rect 16460 11940 16516 11942
rect 20220 13626 20276 13628
rect 20300 13626 20356 13628
rect 20380 13626 20436 13628
rect 20460 13626 20516 13628
rect 20220 13574 20266 13626
rect 20266 13574 20276 13626
rect 20300 13574 20330 13626
rect 20330 13574 20342 13626
rect 20342 13574 20356 13626
rect 20380 13574 20394 13626
rect 20394 13574 20406 13626
rect 20406 13574 20436 13626
rect 20460 13574 20470 13626
rect 20470 13574 20516 13626
rect 20220 13572 20276 13574
rect 20300 13572 20356 13574
rect 20380 13572 20436 13574
rect 20460 13572 20516 13574
rect 20220 12538 20276 12540
rect 20300 12538 20356 12540
rect 20380 12538 20436 12540
rect 20460 12538 20516 12540
rect 20220 12486 20266 12538
rect 20266 12486 20276 12538
rect 20300 12486 20330 12538
rect 20330 12486 20342 12538
rect 20342 12486 20356 12538
rect 20380 12486 20394 12538
rect 20394 12486 20406 12538
rect 20406 12486 20436 12538
rect 20460 12486 20470 12538
rect 20470 12486 20516 12538
rect 20220 12484 20276 12486
rect 20300 12484 20356 12486
rect 20380 12484 20436 12486
rect 20460 12484 20516 12486
rect 16220 10906 16276 10908
rect 16300 10906 16356 10908
rect 16380 10906 16436 10908
rect 16460 10906 16516 10908
rect 16220 10854 16266 10906
rect 16266 10854 16276 10906
rect 16300 10854 16330 10906
rect 16330 10854 16342 10906
rect 16342 10854 16356 10906
rect 16380 10854 16394 10906
rect 16394 10854 16406 10906
rect 16406 10854 16436 10906
rect 16460 10854 16470 10906
rect 16470 10854 16516 10906
rect 16220 10852 16276 10854
rect 16300 10852 16356 10854
rect 16380 10852 16436 10854
rect 16460 10852 16516 10854
rect 16220 9818 16276 9820
rect 16300 9818 16356 9820
rect 16380 9818 16436 9820
rect 16460 9818 16516 9820
rect 16220 9766 16266 9818
rect 16266 9766 16276 9818
rect 16300 9766 16330 9818
rect 16330 9766 16342 9818
rect 16342 9766 16356 9818
rect 16380 9766 16394 9818
rect 16394 9766 16406 9818
rect 16406 9766 16436 9818
rect 16460 9766 16470 9818
rect 16470 9766 16516 9818
rect 16220 9764 16276 9766
rect 16300 9764 16356 9766
rect 16380 9764 16436 9766
rect 16460 9764 16516 9766
rect 16220 8730 16276 8732
rect 16300 8730 16356 8732
rect 16380 8730 16436 8732
rect 16460 8730 16516 8732
rect 16220 8678 16266 8730
rect 16266 8678 16276 8730
rect 16300 8678 16330 8730
rect 16330 8678 16342 8730
rect 16342 8678 16356 8730
rect 16380 8678 16394 8730
rect 16394 8678 16406 8730
rect 16406 8678 16436 8730
rect 16460 8678 16470 8730
rect 16470 8678 16516 8730
rect 16220 8676 16276 8678
rect 16300 8676 16356 8678
rect 16380 8676 16436 8678
rect 16460 8676 16516 8678
rect 16220 7642 16276 7644
rect 16300 7642 16356 7644
rect 16380 7642 16436 7644
rect 16460 7642 16516 7644
rect 16220 7590 16266 7642
rect 16266 7590 16276 7642
rect 16300 7590 16330 7642
rect 16330 7590 16342 7642
rect 16342 7590 16356 7642
rect 16380 7590 16394 7642
rect 16394 7590 16406 7642
rect 16406 7590 16436 7642
rect 16460 7590 16470 7642
rect 16470 7590 16516 7642
rect 16220 7588 16276 7590
rect 16300 7588 16356 7590
rect 16380 7588 16436 7590
rect 16460 7588 16516 7590
rect 20220 11450 20276 11452
rect 20300 11450 20356 11452
rect 20380 11450 20436 11452
rect 20460 11450 20516 11452
rect 20220 11398 20266 11450
rect 20266 11398 20276 11450
rect 20300 11398 20330 11450
rect 20330 11398 20342 11450
rect 20342 11398 20356 11450
rect 20380 11398 20394 11450
rect 20394 11398 20406 11450
rect 20406 11398 20436 11450
rect 20460 11398 20470 11450
rect 20470 11398 20516 11450
rect 20220 11396 20276 11398
rect 20300 11396 20356 11398
rect 20380 11396 20436 11398
rect 20460 11396 20516 11398
rect 20220 10362 20276 10364
rect 20300 10362 20356 10364
rect 20380 10362 20436 10364
rect 20460 10362 20516 10364
rect 20220 10310 20266 10362
rect 20266 10310 20276 10362
rect 20300 10310 20330 10362
rect 20330 10310 20342 10362
rect 20342 10310 20356 10362
rect 20380 10310 20394 10362
rect 20394 10310 20406 10362
rect 20406 10310 20436 10362
rect 20460 10310 20470 10362
rect 20470 10310 20516 10362
rect 20220 10308 20276 10310
rect 20300 10308 20356 10310
rect 20380 10308 20436 10310
rect 20460 10308 20516 10310
rect 20220 9274 20276 9276
rect 20300 9274 20356 9276
rect 20380 9274 20436 9276
rect 20460 9274 20516 9276
rect 20220 9222 20266 9274
rect 20266 9222 20276 9274
rect 20300 9222 20330 9274
rect 20330 9222 20342 9274
rect 20342 9222 20356 9274
rect 20380 9222 20394 9274
rect 20394 9222 20406 9274
rect 20406 9222 20436 9274
rect 20460 9222 20470 9274
rect 20470 9222 20516 9274
rect 20220 9220 20276 9222
rect 20300 9220 20356 9222
rect 20380 9220 20436 9222
rect 20460 9220 20516 9222
rect 20220 8186 20276 8188
rect 20300 8186 20356 8188
rect 20380 8186 20436 8188
rect 20460 8186 20516 8188
rect 20220 8134 20266 8186
rect 20266 8134 20276 8186
rect 20300 8134 20330 8186
rect 20330 8134 20342 8186
rect 20342 8134 20356 8186
rect 20380 8134 20394 8186
rect 20394 8134 20406 8186
rect 20406 8134 20436 8186
rect 20460 8134 20470 8186
rect 20470 8134 20516 8186
rect 20220 8132 20276 8134
rect 20300 8132 20356 8134
rect 20380 8132 20436 8134
rect 20460 8132 20516 8134
rect 22098 7384 22154 7440
rect 20220 7098 20276 7100
rect 20300 7098 20356 7100
rect 20380 7098 20436 7100
rect 20460 7098 20516 7100
rect 20220 7046 20266 7098
rect 20266 7046 20276 7098
rect 20300 7046 20330 7098
rect 20330 7046 20342 7098
rect 20342 7046 20356 7098
rect 20380 7046 20394 7098
rect 20394 7046 20406 7098
rect 20406 7046 20436 7098
rect 20460 7046 20470 7098
rect 20470 7046 20516 7098
rect 20220 7044 20276 7046
rect 20300 7044 20356 7046
rect 20380 7044 20436 7046
rect 20460 7044 20516 7046
rect 16220 6554 16276 6556
rect 16300 6554 16356 6556
rect 16380 6554 16436 6556
rect 16460 6554 16516 6556
rect 16220 6502 16266 6554
rect 16266 6502 16276 6554
rect 16300 6502 16330 6554
rect 16330 6502 16342 6554
rect 16342 6502 16356 6554
rect 16380 6502 16394 6554
rect 16394 6502 16406 6554
rect 16406 6502 16436 6554
rect 16460 6502 16470 6554
rect 16470 6502 16516 6554
rect 16220 6500 16276 6502
rect 16300 6500 16356 6502
rect 16380 6500 16436 6502
rect 16460 6500 16516 6502
rect 20220 6010 20276 6012
rect 20300 6010 20356 6012
rect 20380 6010 20436 6012
rect 20460 6010 20516 6012
rect 20220 5958 20266 6010
rect 20266 5958 20276 6010
rect 20300 5958 20330 6010
rect 20330 5958 20342 6010
rect 20342 5958 20356 6010
rect 20380 5958 20394 6010
rect 20394 5958 20406 6010
rect 20406 5958 20436 6010
rect 20460 5958 20470 6010
rect 20470 5958 20516 6010
rect 20220 5956 20276 5958
rect 20300 5956 20356 5958
rect 20380 5956 20436 5958
rect 20460 5956 20516 5958
rect 16220 5466 16276 5468
rect 16300 5466 16356 5468
rect 16380 5466 16436 5468
rect 16460 5466 16516 5468
rect 16220 5414 16266 5466
rect 16266 5414 16276 5466
rect 16300 5414 16330 5466
rect 16330 5414 16342 5466
rect 16342 5414 16356 5466
rect 16380 5414 16394 5466
rect 16394 5414 16406 5466
rect 16406 5414 16436 5466
rect 16460 5414 16470 5466
rect 16470 5414 16516 5466
rect 16220 5412 16276 5414
rect 16300 5412 16356 5414
rect 16380 5412 16436 5414
rect 16460 5412 16516 5414
rect 11978 2524 11980 2544
rect 11980 2524 12032 2544
rect 12032 2524 12034 2544
rect 11978 2488 12034 2524
rect 12346 2488 12402 2544
rect 12714 2488 12770 2544
rect 11242 1556 11298 1592
rect 11242 1536 11244 1556
rect 11244 1536 11296 1556
rect 11296 1536 11298 1556
rect 12220 1658 12276 1660
rect 12300 1658 12356 1660
rect 12380 1658 12436 1660
rect 12460 1658 12516 1660
rect 12220 1606 12266 1658
rect 12266 1606 12276 1658
rect 12300 1606 12330 1658
rect 12330 1606 12342 1658
rect 12342 1606 12356 1658
rect 12380 1606 12394 1658
rect 12394 1606 12406 1658
rect 12406 1606 12436 1658
rect 12460 1606 12470 1658
rect 12470 1606 12516 1658
rect 12220 1604 12276 1606
rect 12300 1604 12356 1606
rect 12380 1604 12436 1606
rect 12460 1604 12516 1606
rect 20220 4922 20276 4924
rect 20300 4922 20356 4924
rect 20380 4922 20436 4924
rect 20460 4922 20516 4924
rect 20220 4870 20266 4922
rect 20266 4870 20276 4922
rect 20300 4870 20330 4922
rect 20330 4870 20342 4922
rect 20342 4870 20356 4922
rect 20380 4870 20394 4922
rect 20394 4870 20406 4922
rect 20406 4870 20436 4922
rect 20460 4870 20470 4922
rect 20470 4870 20516 4922
rect 20220 4868 20276 4870
rect 20300 4868 20356 4870
rect 20380 4868 20436 4870
rect 20460 4868 20516 4870
rect 16220 4378 16276 4380
rect 16300 4378 16356 4380
rect 16380 4378 16436 4380
rect 16460 4378 16516 4380
rect 16220 4326 16266 4378
rect 16266 4326 16276 4378
rect 16300 4326 16330 4378
rect 16330 4326 16342 4378
rect 16342 4326 16356 4378
rect 16380 4326 16394 4378
rect 16394 4326 16406 4378
rect 16406 4326 16436 4378
rect 16460 4326 16470 4378
rect 16470 4326 16516 4378
rect 16220 4324 16276 4326
rect 16300 4324 16356 4326
rect 16380 4324 16436 4326
rect 16460 4324 16516 4326
rect 20220 3834 20276 3836
rect 20300 3834 20356 3836
rect 20380 3834 20436 3836
rect 20460 3834 20516 3836
rect 20220 3782 20266 3834
rect 20266 3782 20276 3834
rect 20300 3782 20330 3834
rect 20330 3782 20342 3834
rect 20342 3782 20356 3834
rect 20380 3782 20394 3834
rect 20394 3782 20406 3834
rect 20406 3782 20436 3834
rect 20460 3782 20470 3834
rect 20470 3782 20516 3834
rect 20220 3780 20276 3782
rect 20300 3780 20356 3782
rect 20380 3780 20436 3782
rect 20460 3780 20516 3782
rect 14002 2896 14058 2952
rect 14094 2388 14096 2408
rect 14096 2388 14148 2408
rect 14148 2388 14150 2408
rect 14094 2352 14150 2388
rect 16220 3290 16276 3292
rect 16300 3290 16356 3292
rect 16380 3290 16436 3292
rect 16460 3290 16516 3292
rect 16220 3238 16266 3290
rect 16266 3238 16276 3290
rect 16300 3238 16330 3290
rect 16330 3238 16342 3290
rect 16342 3238 16356 3290
rect 16380 3238 16394 3290
rect 16394 3238 16406 3290
rect 16406 3238 16436 3290
rect 16460 3238 16470 3290
rect 16470 3238 16516 3290
rect 16220 3236 16276 3238
rect 16300 3236 16356 3238
rect 16380 3236 16436 3238
rect 16460 3236 16516 3238
rect 20220 2746 20276 2748
rect 20300 2746 20356 2748
rect 20380 2746 20436 2748
rect 20460 2746 20516 2748
rect 20220 2694 20266 2746
rect 20266 2694 20276 2746
rect 20300 2694 20330 2746
rect 20330 2694 20342 2746
rect 20342 2694 20356 2746
rect 20380 2694 20394 2746
rect 20394 2694 20406 2746
rect 20406 2694 20436 2746
rect 20460 2694 20470 2746
rect 20470 2694 20516 2746
rect 20220 2692 20276 2694
rect 20300 2692 20356 2694
rect 20380 2692 20436 2694
rect 20460 2692 20516 2694
rect 22098 2488 22154 2544
rect 16220 2202 16276 2204
rect 16300 2202 16356 2204
rect 16380 2202 16436 2204
rect 16460 2202 16516 2204
rect 16220 2150 16266 2202
rect 16266 2150 16276 2202
rect 16300 2150 16330 2202
rect 16330 2150 16342 2202
rect 16342 2150 16356 2202
rect 16380 2150 16394 2202
rect 16394 2150 16406 2202
rect 16406 2150 16436 2202
rect 16460 2150 16470 2202
rect 16470 2150 16516 2202
rect 16220 2148 16276 2150
rect 16300 2148 16356 2150
rect 16380 2148 16436 2150
rect 16460 2148 16516 2150
rect 20258 1964 20314 2000
rect 20258 1944 20260 1964
rect 20260 1944 20312 1964
rect 20312 1944 20314 1964
rect 16220 1114 16276 1116
rect 16300 1114 16356 1116
rect 16380 1114 16436 1116
rect 16460 1114 16516 1116
rect 16220 1062 16266 1114
rect 16266 1062 16276 1114
rect 16300 1062 16330 1114
rect 16330 1062 16342 1114
rect 16342 1062 16356 1114
rect 16380 1062 16394 1114
rect 16394 1062 16406 1114
rect 16406 1062 16436 1114
rect 16460 1062 16470 1114
rect 16470 1062 16516 1114
rect 16220 1060 16276 1062
rect 16300 1060 16356 1062
rect 16380 1060 16436 1062
rect 16460 1060 16516 1062
rect 20220 1658 20276 1660
rect 20300 1658 20356 1660
rect 20380 1658 20436 1660
rect 20460 1658 20516 1660
rect 20220 1606 20266 1658
rect 20266 1606 20276 1658
rect 20300 1606 20330 1658
rect 20330 1606 20342 1658
rect 20342 1606 20356 1658
rect 20380 1606 20394 1658
rect 20394 1606 20406 1658
rect 20406 1606 20436 1658
rect 20460 1606 20470 1658
rect 20470 1606 20516 1658
rect 20220 1604 20276 1606
rect 20300 1604 20356 1606
rect 20380 1604 20436 1606
rect 20460 1604 20516 1606
<< metal3 >>
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 12210 13632 12526 13633
rect 12210 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12526 13632
rect 12210 13567 12526 13568
rect 20210 13632 20526 13633
rect 20210 13568 20216 13632
rect 20280 13568 20296 13632
rect 20360 13568 20376 13632
rect 20440 13568 20456 13632
rect 20520 13568 20526 13632
rect 20210 13567 20526 13568
rect 10225 13290 10291 13293
rect 2730 13288 10291 13290
rect 2730 13232 10230 13288
rect 10286 13232 10291 13288
rect 2730 13230 10291 13232
rect 0 13154 800 13184
rect 2730 13154 2790 13230
rect 10225 13227 10291 13230
rect 0 13094 2790 13154
rect 0 13064 800 13094
rect 8210 13088 8526 13089
rect 8210 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8526 13088
rect 8210 13023 8526 13024
rect 16210 13088 16526 13089
rect 16210 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16526 13088
rect 16210 13023 16526 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 12210 12544 12526 12545
rect 12210 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12526 12544
rect 12210 12479 12526 12480
rect 20210 12544 20526 12545
rect 20210 12480 20216 12544
rect 20280 12480 20296 12544
rect 20360 12480 20376 12544
rect 20440 12480 20456 12544
rect 20520 12480 20526 12544
rect 20210 12479 20526 12480
rect 0 12338 800 12368
rect 5533 12338 5599 12341
rect 0 12336 5599 12338
rect 0 12280 5538 12336
rect 5594 12280 5599 12336
rect 0 12278 5599 12280
rect 0 12248 800 12278
rect 5533 12275 5599 12278
rect 23200 12248 24000 12368
rect 8210 12000 8526 12001
rect 8210 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8526 12000
rect 8210 11935 8526 11936
rect 16210 12000 16526 12001
rect 16210 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16526 12000
rect 16210 11935 16526 11936
rect 0 11522 800 11552
rect 1761 11522 1827 11525
rect 0 11520 1827 11522
rect 0 11464 1766 11520
rect 1822 11464 1827 11520
rect 0 11462 1827 11464
rect 0 11432 800 11462
rect 1761 11459 1827 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 12210 11456 12526 11457
rect 12210 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12526 11456
rect 12210 11391 12526 11392
rect 20210 11456 20526 11457
rect 20210 11392 20216 11456
rect 20280 11392 20296 11456
rect 20360 11392 20376 11456
rect 20440 11392 20456 11456
rect 20520 11392 20526 11456
rect 20210 11391 20526 11392
rect 8210 10912 8526 10913
rect 8210 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8526 10912
rect 8210 10847 8526 10848
rect 16210 10912 16526 10913
rect 16210 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16526 10912
rect 16210 10847 16526 10848
rect 0 10706 800 10736
rect 11605 10706 11671 10709
rect 0 10704 11671 10706
rect 0 10648 11610 10704
rect 11666 10648 11671 10704
rect 0 10646 11671 10648
rect 0 10616 800 10646
rect 11605 10643 11671 10646
rect 7833 10570 7899 10573
rect 9581 10570 9647 10573
rect 7833 10568 9647 10570
rect 7833 10512 7838 10568
rect 7894 10512 9586 10568
rect 9642 10512 9647 10568
rect 7833 10510 9647 10512
rect 7833 10507 7899 10510
rect 9581 10507 9647 10510
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 12210 10368 12526 10369
rect 12210 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12526 10368
rect 12210 10303 12526 10304
rect 20210 10368 20526 10369
rect 20210 10304 20216 10368
rect 20280 10304 20296 10368
rect 20360 10304 20376 10368
rect 20440 10304 20456 10368
rect 20520 10304 20526 10368
rect 20210 10303 20526 10304
rect 13905 10026 13971 10029
rect 2730 10024 13971 10026
rect 2730 9968 13910 10024
rect 13966 9968 13971 10024
rect 2730 9966 13971 9968
rect 0 9890 800 9920
rect 2730 9890 2790 9966
rect 13905 9963 13971 9966
rect 0 9830 2790 9890
rect 5441 9890 5507 9893
rect 7005 9890 7071 9893
rect 7833 9890 7899 9893
rect 5441 9888 7899 9890
rect 5441 9832 5446 9888
rect 5502 9832 7010 9888
rect 7066 9832 7838 9888
rect 7894 9832 7899 9888
rect 5441 9830 7899 9832
rect 0 9800 800 9830
rect 5441 9827 5507 9830
rect 7005 9827 7071 9830
rect 7833 9827 7899 9830
rect 8210 9824 8526 9825
rect 8210 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8526 9824
rect 8210 9759 8526 9760
rect 16210 9824 16526 9825
rect 16210 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16526 9824
rect 16210 9759 16526 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 12210 9280 12526 9281
rect 12210 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12526 9280
rect 12210 9215 12526 9216
rect 20210 9280 20526 9281
rect 20210 9216 20216 9280
rect 20280 9216 20296 9280
rect 20360 9216 20376 9280
rect 20440 9216 20456 9280
rect 20520 9216 20526 9280
rect 20210 9215 20526 9216
rect 10593 9210 10659 9213
rect 11697 9210 11763 9213
rect 10593 9208 11763 9210
rect 10593 9152 10598 9208
rect 10654 9152 11702 9208
rect 11758 9152 11763 9208
rect 10593 9150 11763 9152
rect 10593 9147 10659 9150
rect 11697 9147 11763 9150
rect 0 9074 800 9104
rect 6453 9074 6519 9077
rect 0 9072 6519 9074
rect 0 9016 6458 9072
rect 6514 9016 6519 9072
rect 0 9014 6519 9016
rect 0 8984 800 9014
rect 6453 9011 6519 9014
rect 8210 8736 8526 8737
rect 8210 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8526 8736
rect 8210 8671 8526 8672
rect 16210 8736 16526 8737
rect 16210 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16526 8736
rect 16210 8671 16526 8672
rect 0 8258 800 8288
rect 1577 8258 1643 8261
rect 0 8256 1643 8258
rect 0 8200 1582 8256
rect 1638 8200 1643 8256
rect 0 8198 1643 8200
rect 0 8168 800 8198
rect 1577 8195 1643 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 12210 8192 12526 8193
rect 12210 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12526 8192
rect 12210 8127 12526 8128
rect 20210 8192 20526 8193
rect 20210 8128 20216 8192
rect 20280 8128 20296 8192
rect 20360 8128 20376 8192
rect 20440 8128 20456 8192
rect 20520 8128 20526 8192
rect 20210 8127 20526 8128
rect 8210 7648 8526 7649
rect 8210 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8526 7648
rect 8210 7583 8526 7584
rect 16210 7648 16526 7649
rect 16210 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16526 7648
rect 16210 7583 16526 7584
rect 0 7442 800 7472
rect 7005 7442 7071 7445
rect 0 7440 7071 7442
rect 0 7384 7010 7440
rect 7066 7384 7071 7440
rect 0 7382 7071 7384
rect 0 7352 800 7382
rect 7005 7379 7071 7382
rect 22093 7442 22159 7445
rect 23200 7442 24000 7472
rect 22093 7440 24000 7442
rect 22093 7384 22098 7440
rect 22154 7384 24000 7440
rect 22093 7382 24000 7384
rect 22093 7379 22159 7382
rect 23200 7352 24000 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 12210 7104 12526 7105
rect 12210 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12526 7104
rect 12210 7039 12526 7040
rect 20210 7104 20526 7105
rect 20210 7040 20216 7104
rect 20280 7040 20296 7104
rect 20360 7040 20376 7104
rect 20440 7040 20456 7104
rect 20520 7040 20526 7104
rect 20210 7039 20526 7040
rect 0 6626 800 6656
rect 6177 6626 6243 6629
rect 0 6624 6243 6626
rect 0 6568 6182 6624
rect 6238 6568 6243 6624
rect 0 6566 6243 6568
rect 0 6536 800 6566
rect 6177 6563 6243 6566
rect 8210 6560 8526 6561
rect 8210 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8526 6560
rect 8210 6495 8526 6496
rect 16210 6560 16526 6561
rect 16210 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16526 6560
rect 16210 6495 16526 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 12210 6016 12526 6017
rect 12210 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12526 6016
rect 12210 5951 12526 5952
rect 20210 6016 20526 6017
rect 20210 5952 20216 6016
rect 20280 5952 20296 6016
rect 20360 5952 20376 6016
rect 20440 5952 20456 6016
rect 20520 5952 20526 6016
rect 20210 5951 20526 5952
rect 0 5810 800 5840
rect 1301 5810 1367 5813
rect 0 5808 1367 5810
rect 0 5752 1306 5808
rect 1362 5752 1367 5808
rect 0 5750 1367 5752
rect 0 5720 800 5750
rect 1301 5747 1367 5750
rect 6177 5810 6243 5813
rect 7373 5810 7439 5813
rect 6177 5808 7439 5810
rect 6177 5752 6182 5808
rect 6238 5752 7378 5808
rect 7434 5752 7439 5808
rect 6177 5750 7439 5752
rect 6177 5747 6243 5750
rect 7373 5747 7439 5750
rect 8210 5472 8526 5473
rect 8210 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8526 5472
rect 8210 5407 8526 5408
rect 16210 5472 16526 5473
rect 16210 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16526 5472
rect 16210 5407 16526 5408
rect 0 4994 800 5024
rect 0 4934 2790 4994
rect 0 4904 800 4934
rect 2730 4722 2790 4934
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 12210 4928 12526 4929
rect 12210 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12526 4928
rect 12210 4863 12526 4864
rect 20210 4928 20526 4929
rect 20210 4864 20216 4928
rect 20280 4864 20296 4928
rect 20360 4864 20376 4928
rect 20440 4864 20456 4928
rect 20520 4864 20526 4928
rect 20210 4863 20526 4864
rect 4705 4722 4771 4725
rect 2730 4720 4771 4722
rect 2730 4664 4710 4720
rect 4766 4664 4771 4720
rect 2730 4662 4771 4664
rect 4705 4659 4771 4662
rect 8210 4384 8526 4385
rect 8210 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8526 4384
rect 8210 4319 8526 4320
rect 16210 4384 16526 4385
rect 16210 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16526 4384
rect 16210 4319 16526 4320
rect 0 4178 800 4208
rect 2405 4178 2471 4181
rect 0 4176 2471 4178
rect 0 4120 2410 4176
rect 2466 4120 2471 4176
rect 0 4118 2471 4120
rect 0 4088 800 4118
rect 2405 4115 2471 4118
rect 3877 4042 3943 4045
rect 5901 4042 5967 4045
rect 3877 4040 5967 4042
rect 3877 3984 3882 4040
rect 3938 3984 5906 4040
rect 5962 3984 5967 4040
rect 3877 3982 5967 3984
rect 3877 3979 3943 3982
rect 5901 3979 5967 3982
rect 4797 3906 4863 3909
rect 8293 3906 8359 3909
rect 9489 3906 9555 3909
rect 4797 3904 9555 3906
rect 4797 3848 4802 3904
rect 4858 3848 8298 3904
rect 8354 3848 9494 3904
rect 9550 3848 9555 3904
rect 4797 3846 9555 3848
rect 4797 3843 4863 3846
rect 8293 3843 8359 3846
rect 9489 3843 9555 3846
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 12210 3840 12526 3841
rect 12210 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12526 3840
rect 12210 3775 12526 3776
rect 20210 3840 20526 3841
rect 20210 3776 20216 3840
rect 20280 3776 20296 3840
rect 20360 3776 20376 3840
rect 20440 3776 20456 3840
rect 20520 3776 20526 3840
rect 20210 3775 20526 3776
rect 2405 3634 2471 3637
rect 8937 3634 9003 3637
rect 2405 3632 9003 3634
rect 2405 3576 2410 3632
rect 2466 3576 8942 3632
rect 8998 3576 9003 3632
rect 2405 3574 9003 3576
rect 2405 3571 2471 3574
rect 8937 3571 9003 3574
rect 4521 3498 4587 3501
rect 6729 3498 6795 3501
rect 4521 3496 6795 3498
rect 4521 3440 4526 3496
rect 4582 3440 6734 3496
rect 6790 3440 6795 3496
rect 4521 3438 6795 3440
rect 4521 3435 4587 3438
rect 6729 3435 6795 3438
rect 0 3362 800 3392
rect 1301 3362 1367 3365
rect 0 3360 1367 3362
rect 0 3304 1306 3360
rect 1362 3304 1367 3360
rect 0 3302 1367 3304
rect 0 3272 800 3302
rect 1301 3299 1367 3302
rect 8210 3296 8526 3297
rect 8210 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8526 3296
rect 8210 3231 8526 3232
rect 16210 3296 16526 3297
rect 16210 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16526 3296
rect 16210 3231 16526 3232
rect 3049 2954 3115 2957
rect 5809 2954 5875 2957
rect 3049 2952 5875 2954
rect 3049 2896 3054 2952
rect 3110 2896 5814 2952
rect 5870 2896 5875 2952
rect 3049 2894 5875 2896
rect 3049 2891 3115 2894
rect 5809 2891 5875 2894
rect 9121 2954 9187 2957
rect 13997 2954 14063 2957
rect 9121 2952 14063 2954
rect 9121 2896 9126 2952
rect 9182 2896 14002 2952
rect 14058 2896 14063 2952
rect 9121 2894 14063 2896
rect 9121 2891 9187 2894
rect 13997 2891 14063 2894
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 12210 2752 12526 2753
rect 12210 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12526 2752
rect 12210 2687 12526 2688
rect 20210 2752 20526 2753
rect 20210 2688 20216 2752
rect 20280 2688 20296 2752
rect 20360 2688 20376 2752
rect 20440 2688 20456 2752
rect 20520 2688 20526 2752
rect 20210 2687 20526 2688
rect 0 2546 800 2576
rect 1761 2546 1827 2549
rect 0 2544 1827 2546
rect 0 2488 1766 2544
rect 1822 2488 1827 2544
rect 0 2486 1827 2488
rect 0 2456 800 2486
rect 1761 2483 1827 2486
rect 10317 2546 10383 2549
rect 11973 2546 12039 2549
rect 10317 2544 12039 2546
rect 10317 2488 10322 2544
rect 10378 2488 11978 2544
rect 12034 2488 12039 2544
rect 10317 2486 12039 2488
rect 10317 2483 10383 2486
rect 11973 2483 12039 2486
rect 12341 2546 12407 2549
rect 12709 2546 12775 2549
rect 12341 2544 12775 2546
rect 12341 2488 12346 2544
rect 12402 2488 12714 2544
rect 12770 2488 12775 2544
rect 12341 2486 12775 2488
rect 12341 2483 12407 2486
rect 12709 2483 12775 2486
rect 22093 2546 22159 2549
rect 23200 2546 24000 2576
rect 22093 2544 24000 2546
rect 22093 2488 22098 2544
rect 22154 2488 24000 2544
rect 22093 2486 24000 2488
rect 22093 2483 22159 2486
rect 23200 2456 24000 2486
rect 2589 2410 2655 2413
rect 14089 2410 14155 2413
rect 2589 2408 14155 2410
rect 2589 2352 2594 2408
rect 2650 2352 14094 2408
rect 14150 2352 14155 2408
rect 2589 2350 14155 2352
rect 2589 2347 2655 2350
rect 14089 2347 14155 2350
rect 8210 2208 8526 2209
rect 8210 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8526 2208
rect 8210 2143 8526 2144
rect 16210 2208 16526 2209
rect 16210 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16526 2208
rect 16210 2143 16526 2144
rect 3693 2002 3759 2005
rect 5993 2002 6059 2005
rect 3693 2000 6059 2002
rect 3693 1944 3698 2000
rect 3754 1944 5998 2000
rect 6054 1944 6059 2000
rect 3693 1942 6059 1944
rect 3693 1939 3759 1942
rect 5993 1939 6059 1942
rect 8017 2002 8083 2005
rect 20253 2002 20319 2005
rect 8017 2000 20319 2002
rect 8017 1944 8022 2000
rect 8078 1944 20258 2000
rect 20314 1944 20319 2000
rect 8017 1942 20319 1944
rect 8017 1939 8083 1942
rect 20253 1939 20319 1942
rect 6361 1866 6427 1869
rect 6637 1866 6703 1869
rect 2730 1864 6703 1866
rect 2730 1808 6366 1864
rect 6422 1808 6642 1864
rect 6698 1808 6703 1864
rect 2730 1806 6703 1808
rect 0 1730 800 1760
rect 2730 1730 2790 1806
rect 6361 1803 6427 1806
rect 6637 1803 6703 1806
rect 6821 1866 6887 1869
rect 9305 1866 9371 1869
rect 10777 1866 10843 1869
rect 6821 1864 10843 1866
rect 6821 1808 6826 1864
rect 6882 1808 9310 1864
rect 9366 1808 10782 1864
rect 10838 1808 10843 1864
rect 6821 1806 10843 1808
rect 6821 1803 6887 1806
rect 9305 1803 9371 1806
rect 10777 1803 10843 1806
rect 0 1670 2790 1730
rect 0 1640 800 1670
rect 4210 1664 4526 1665
rect 4210 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4526 1664
rect 4210 1599 4526 1600
rect 12210 1664 12526 1665
rect 12210 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12526 1664
rect 12210 1599 12526 1600
rect 20210 1664 20526 1665
rect 20210 1600 20216 1664
rect 20280 1600 20296 1664
rect 20360 1600 20376 1664
rect 20440 1600 20456 1664
rect 20520 1600 20526 1664
rect 20210 1599 20526 1600
rect 5073 1594 5139 1597
rect 11237 1594 11303 1597
rect 5073 1592 11303 1594
rect 5073 1536 5078 1592
rect 5134 1536 11242 1592
rect 11298 1536 11303 1592
rect 5073 1534 11303 1536
rect 5073 1531 5139 1534
rect 11237 1531 11303 1534
rect 8210 1120 8526 1121
rect 8210 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8526 1120
rect 8210 1055 8526 1056
rect 16210 1120 16526 1121
rect 16210 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16526 1120
rect 16210 1055 16526 1056
<< via3 >>
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 12216 13628 12280 13632
rect 12216 13572 12220 13628
rect 12220 13572 12276 13628
rect 12276 13572 12280 13628
rect 12216 13568 12280 13572
rect 12296 13628 12360 13632
rect 12296 13572 12300 13628
rect 12300 13572 12356 13628
rect 12356 13572 12360 13628
rect 12296 13568 12360 13572
rect 12376 13628 12440 13632
rect 12376 13572 12380 13628
rect 12380 13572 12436 13628
rect 12436 13572 12440 13628
rect 12376 13568 12440 13572
rect 12456 13628 12520 13632
rect 12456 13572 12460 13628
rect 12460 13572 12516 13628
rect 12516 13572 12520 13628
rect 12456 13568 12520 13572
rect 20216 13628 20280 13632
rect 20216 13572 20220 13628
rect 20220 13572 20276 13628
rect 20276 13572 20280 13628
rect 20216 13568 20280 13572
rect 20296 13628 20360 13632
rect 20296 13572 20300 13628
rect 20300 13572 20356 13628
rect 20356 13572 20360 13628
rect 20296 13568 20360 13572
rect 20376 13628 20440 13632
rect 20376 13572 20380 13628
rect 20380 13572 20436 13628
rect 20436 13572 20440 13628
rect 20376 13568 20440 13572
rect 20456 13628 20520 13632
rect 20456 13572 20460 13628
rect 20460 13572 20516 13628
rect 20516 13572 20520 13628
rect 20456 13568 20520 13572
rect 8216 13084 8280 13088
rect 8216 13028 8220 13084
rect 8220 13028 8276 13084
rect 8276 13028 8280 13084
rect 8216 13024 8280 13028
rect 8296 13084 8360 13088
rect 8296 13028 8300 13084
rect 8300 13028 8356 13084
rect 8356 13028 8360 13084
rect 8296 13024 8360 13028
rect 8376 13084 8440 13088
rect 8376 13028 8380 13084
rect 8380 13028 8436 13084
rect 8436 13028 8440 13084
rect 8376 13024 8440 13028
rect 8456 13084 8520 13088
rect 8456 13028 8460 13084
rect 8460 13028 8516 13084
rect 8516 13028 8520 13084
rect 8456 13024 8520 13028
rect 16216 13084 16280 13088
rect 16216 13028 16220 13084
rect 16220 13028 16276 13084
rect 16276 13028 16280 13084
rect 16216 13024 16280 13028
rect 16296 13084 16360 13088
rect 16296 13028 16300 13084
rect 16300 13028 16356 13084
rect 16356 13028 16360 13084
rect 16296 13024 16360 13028
rect 16376 13084 16440 13088
rect 16376 13028 16380 13084
rect 16380 13028 16436 13084
rect 16436 13028 16440 13084
rect 16376 13024 16440 13028
rect 16456 13084 16520 13088
rect 16456 13028 16460 13084
rect 16460 13028 16516 13084
rect 16516 13028 16520 13084
rect 16456 13024 16520 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 12216 12540 12280 12544
rect 12216 12484 12220 12540
rect 12220 12484 12276 12540
rect 12276 12484 12280 12540
rect 12216 12480 12280 12484
rect 12296 12540 12360 12544
rect 12296 12484 12300 12540
rect 12300 12484 12356 12540
rect 12356 12484 12360 12540
rect 12296 12480 12360 12484
rect 12376 12540 12440 12544
rect 12376 12484 12380 12540
rect 12380 12484 12436 12540
rect 12436 12484 12440 12540
rect 12376 12480 12440 12484
rect 12456 12540 12520 12544
rect 12456 12484 12460 12540
rect 12460 12484 12516 12540
rect 12516 12484 12520 12540
rect 12456 12480 12520 12484
rect 20216 12540 20280 12544
rect 20216 12484 20220 12540
rect 20220 12484 20276 12540
rect 20276 12484 20280 12540
rect 20216 12480 20280 12484
rect 20296 12540 20360 12544
rect 20296 12484 20300 12540
rect 20300 12484 20356 12540
rect 20356 12484 20360 12540
rect 20296 12480 20360 12484
rect 20376 12540 20440 12544
rect 20376 12484 20380 12540
rect 20380 12484 20436 12540
rect 20436 12484 20440 12540
rect 20376 12480 20440 12484
rect 20456 12540 20520 12544
rect 20456 12484 20460 12540
rect 20460 12484 20516 12540
rect 20516 12484 20520 12540
rect 20456 12480 20520 12484
rect 8216 11996 8280 12000
rect 8216 11940 8220 11996
rect 8220 11940 8276 11996
rect 8276 11940 8280 11996
rect 8216 11936 8280 11940
rect 8296 11996 8360 12000
rect 8296 11940 8300 11996
rect 8300 11940 8356 11996
rect 8356 11940 8360 11996
rect 8296 11936 8360 11940
rect 8376 11996 8440 12000
rect 8376 11940 8380 11996
rect 8380 11940 8436 11996
rect 8436 11940 8440 11996
rect 8376 11936 8440 11940
rect 8456 11996 8520 12000
rect 8456 11940 8460 11996
rect 8460 11940 8516 11996
rect 8516 11940 8520 11996
rect 8456 11936 8520 11940
rect 16216 11996 16280 12000
rect 16216 11940 16220 11996
rect 16220 11940 16276 11996
rect 16276 11940 16280 11996
rect 16216 11936 16280 11940
rect 16296 11996 16360 12000
rect 16296 11940 16300 11996
rect 16300 11940 16356 11996
rect 16356 11940 16360 11996
rect 16296 11936 16360 11940
rect 16376 11996 16440 12000
rect 16376 11940 16380 11996
rect 16380 11940 16436 11996
rect 16436 11940 16440 11996
rect 16376 11936 16440 11940
rect 16456 11996 16520 12000
rect 16456 11940 16460 11996
rect 16460 11940 16516 11996
rect 16516 11940 16520 11996
rect 16456 11936 16520 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 12216 11452 12280 11456
rect 12216 11396 12220 11452
rect 12220 11396 12276 11452
rect 12276 11396 12280 11452
rect 12216 11392 12280 11396
rect 12296 11452 12360 11456
rect 12296 11396 12300 11452
rect 12300 11396 12356 11452
rect 12356 11396 12360 11452
rect 12296 11392 12360 11396
rect 12376 11452 12440 11456
rect 12376 11396 12380 11452
rect 12380 11396 12436 11452
rect 12436 11396 12440 11452
rect 12376 11392 12440 11396
rect 12456 11452 12520 11456
rect 12456 11396 12460 11452
rect 12460 11396 12516 11452
rect 12516 11396 12520 11452
rect 12456 11392 12520 11396
rect 20216 11452 20280 11456
rect 20216 11396 20220 11452
rect 20220 11396 20276 11452
rect 20276 11396 20280 11452
rect 20216 11392 20280 11396
rect 20296 11452 20360 11456
rect 20296 11396 20300 11452
rect 20300 11396 20356 11452
rect 20356 11396 20360 11452
rect 20296 11392 20360 11396
rect 20376 11452 20440 11456
rect 20376 11396 20380 11452
rect 20380 11396 20436 11452
rect 20436 11396 20440 11452
rect 20376 11392 20440 11396
rect 20456 11452 20520 11456
rect 20456 11396 20460 11452
rect 20460 11396 20516 11452
rect 20516 11396 20520 11452
rect 20456 11392 20520 11396
rect 8216 10908 8280 10912
rect 8216 10852 8220 10908
rect 8220 10852 8276 10908
rect 8276 10852 8280 10908
rect 8216 10848 8280 10852
rect 8296 10908 8360 10912
rect 8296 10852 8300 10908
rect 8300 10852 8356 10908
rect 8356 10852 8360 10908
rect 8296 10848 8360 10852
rect 8376 10908 8440 10912
rect 8376 10852 8380 10908
rect 8380 10852 8436 10908
rect 8436 10852 8440 10908
rect 8376 10848 8440 10852
rect 8456 10908 8520 10912
rect 8456 10852 8460 10908
rect 8460 10852 8516 10908
rect 8516 10852 8520 10908
rect 8456 10848 8520 10852
rect 16216 10908 16280 10912
rect 16216 10852 16220 10908
rect 16220 10852 16276 10908
rect 16276 10852 16280 10908
rect 16216 10848 16280 10852
rect 16296 10908 16360 10912
rect 16296 10852 16300 10908
rect 16300 10852 16356 10908
rect 16356 10852 16360 10908
rect 16296 10848 16360 10852
rect 16376 10908 16440 10912
rect 16376 10852 16380 10908
rect 16380 10852 16436 10908
rect 16436 10852 16440 10908
rect 16376 10848 16440 10852
rect 16456 10908 16520 10912
rect 16456 10852 16460 10908
rect 16460 10852 16516 10908
rect 16516 10852 16520 10908
rect 16456 10848 16520 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 12216 10364 12280 10368
rect 12216 10308 12220 10364
rect 12220 10308 12276 10364
rect 12276 10308 12280 10364
rect 12216 10304 12280 10308
rect 12296 10364 12360 10368
rect 12296 10308 12300 10364
rect 12300 10308 12356 10364
rect 12356 10308 12360 10364
rect 12296 10304 12360 10308
rect 12376 10364 12440 10368
rect 12376 10308 12380 10364
rect 12380 10308 12436 10364
rect 12436 10308 12440 10364
rect 12376 10304 12440 10308
rect 12456 10364 12520 10368
rect 12456 10308 12460 10364
rect 12460 10308 12516 10364
rect 12516 10308 12520 10364
rect 12456 10304 12520 10308
rect 20216 10364 20280 10368
rect 20216 10308 20220 10364
rect 20220 10308 20276 10364
rect 20276 10308 20280 10364
rect 20216 10304 20280 10308
rect 20296 10364 20360 10368
rect 20296 10308 20300 10364
rect 20300 10308 20356 10364
rect 20356 10308 20360 10364
rect 20296 10304 20360 10308
rect 20376 10364 20440 10368
rect 20376 10308 20380 10364
rect 20380 10308 20436 10364
rect 20436 10308 20440 10364
rect 20376 10304 20440 10308
rect 20456 10364 20520 10368
rect 20456 10308 20460 10364
rect 20460 10308 20516 10364
rect 20516 10308 20520 10364
rect 20456 10304 20520 10308
rect 8216 9820 8280 9824
rect 8216 9764 8220 9820
rect 8220 9764 8276 9820
rect 8276 9764 8280 9820
rect 8216 9760 8280 9764
rect 8296 9820 8360 9824
rect 8296 9764 8300 9820
rect 8300 9764 8356 9820
rect 8356 9764 8360 9820
rect 8296 9760 8360 9764
rect 8376 9820 8440 9824
rect 8376 9764 8380 9820
rect 8380 9764 8436 9820
rect 8436 9764 8440 9820
rect 8376 9760 8440 9764
rect 8456 9820 8520 9824
rect 8456 9764 8460 9820
rect 8460 9764 8516 9820
rect 8516 9764 8520 9820
rect 8456 9760 8520 9764
rect 16216 9820 16280 9824
rect 16216 9764 16220 9820
rect 16220 9764 16276 9820
rect 16276 9764 16280 9820
rect 16216 9760 16280 9764
rect 16296 9820 16360 9824
rect 16296 9764 16300 9820
rect 16300 9764 16356 9820
rect 16356 9764 16360 9820
rect 16296 9760 16360 9764
rect 16376 9820 16440 9824
rect 16376 9764 16380 9820
rect 16380 9764 16436 9820
rect 16436 9764 16440 9820
rect 16376 9760 16440 9764
rect 16456 9820 16520 9824
rect 16456 9764 16460 9820
rect 16460 9764 16516 9820
rect 16516 9764 16520 9820
rect 16456 9760 16520 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 12216 9276 12280 9280
rect 12216 9220 12220 9276
rect 12220 9220 12276 9276
rect 12276 9220 12280 9276
rect 12216 9216 12280 9220
rect 12296 9276 12360 9280
rect 12296 9220 12300 9276
rect 12300 9220 12356 9276
rect 12356 9220 12360 9276
rect 12296 9216 12360 9220
rect 12376 9276 12440 9280
rect 12376 9220 12380 9276
rect 12380 9220 12436 9276
rect 12436 9220 12440 9276
rect 12376 9216 12440 9220
rect 12456 9276 12520 9280
rect 12456 9220 12460 9276
rect 12460 9220 12516 9276
rect 12516 9220 12520 9276
rect 12456 9216 12520 9220
rect 20216 9276 20280 9280
rect 20216 9220 20220 9276
rect 20220 9220 20276 9276
rect 20276 9220 20280 9276
rect 20216 9216 20280 9220
rect 20296 9276 20360 9280
rect 20296 9220 20300 9276
rect 20300 9220 20356 9276
rect 20356 9220 20360 9276
rect 20296 9216 20360 9220
rect 20376 9276 20440 9280
rect 20376 9220 20380 9276
rect 20380 9220 20436 9276
rect 20436 9220 20440 9276
rect 20376 9216 20440 9220
rect 20456 9276 20520 9280
rect 20456 9220 20460 9276
rect 20460 9220 20516 9276
rect 20516 9220 20520 9276
rect 20456 9216 20520 9220
rect 8216 8732 8280 8736
rect 8216 8676 8220 8732
rect 8220 8676 8276 8732
rect 8276 8676 8280 8732
rect 8216 8672 8280 8676
rect 8296 8732 8360 8736
rect 8296 8676 8300 8732
rect 8300 8676 8356 8732
rect 8356 8676 8360 8732
rect 8296 8672 8360 8676
rect 8376 8732 8440 8736
rect 8376 8676 8380 8732
rect 8380 8676 8436 8732
rect 8436 8676 8440 8732
rect 8376 8672 8440 8676
rect 8456 8732 8520 8736
rect 8456 8676 8460 8732
rect 8460 8676 8516 8732
rect 8516 8676 8520 8732
rect 8456 8672 8520 8676
rect 16216 8732 16280 8736
rect 16216 8676 16220 8732
rect 16220 8676 16276 8732
rect 16276 8676 16280 8732
rect 16216 8672 16280 8676
rect 16296 8732 16360 8736
rect 16296 8676 16300 8732
rect 16300 8676 16356 8732
rect 16356 8676 16360 8732
rect 16296 8672 16360 8676
rect 16376 8732 16440 8736
rect 16376 8676 16380 8732
rect 16380 8676 16436 8732
rect 16436 8676 16440 8732
rect 16376 8672 16440 8676
rect 16456 8732 16520 8736
rect 16456 8676 16460 8732
rect 16460 8676 16516 8732
rect 16516 8676 16520 8732
rect 16456 8672 16520 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 12216 8188 12280 8192
rect 12216 8132 12220 8188
rect 12220 8132 12276 8188
rect 12276 8132 12280 8188
rect 12216 8128 12280 8132
rect 12296 8188 12360 8192
rect 12296 8132 12300 8188
rect 12300 8132 12356 8188
rect 12356 8132 12360 8188
rect 12296 8128 12360 8132
rect 12376 8188 12440 8192
rect 12376 8132 12380 8188
rect 12380 8132 12436 8188
rect 12436 8132 12440 8188
rect 12376 8128 12440 8132
rect 12456 8188 12520 8192
rect 12456 8132 12460 8188
rect 12460 8132 12516 8188
rect 12516 8132 12520 8188
rect 12456 8128 12520 8132
rect 20216 8188 20280 8192
rect 20216 8132 20220 8188
rect 20220 8132 20276 8188
rect 20276 8132 20280 8188
rect 20216 8128 20280 8132
rect 20296 8188 20360 8192
rect 20296 8132 20300 8188
rect 20300 8132 20356 8188
rect 20356 8132 20360 8188
rect 20296 8128 20360 8132
rect 20376 8188 20440 8192
rect 20376 8132 20380 8188
rect 20380 8132 20436 8188
rect 20436 8132 20440 8188
rect 20376 8128 20440 8132
rect 20456 8188 20520 8192
rect 20456 8132 20460 8188
rect 20460 8132 20516 8188
rect 20516 8132 20520 8188
rect 20456 8128 20520 8132
rect 8216 7644 8280 7648
rect 8216 7588 8220 7644
rect 8220 7588 8276 7644
rect 8276 7588 8280 7644
rect 8216 7584 8280 7588
rect 8296 7644 8360 7648
rect 8296 7588 8300 7644
rect 8300 7588 8356 7644
rect 8356 7588 8360 7644
rect 8296 7584 8360 7588
rect 8376 7644 8440 7648
rect 8376 7588 8380 7644
rect 8380 7588 8436 7644
rect 8436 7588 8440 7644
rect 8376 7584 8440 7588
rect 8456 7644 8520 7648
rect 8456 7588 8460 7644
rect 8460 7588 8516 7644
rect 8516 7588 8520 7644
rect 8456 7584 8520 7588
rect 16216 7644 16280 7648
rect 16216 7588 16220 7644
rect 16220 7588 16276 7644
rect 16276 7588 16280 7644
rect 16216 7584 16280 7588
rect 16296 7644 16360 7648
rect 16296 7588 16300 7644
rect 16300 7588 16356 7644
rect 16356 7588 16360 7644
rect 16296 7584 16360 7588
rect 16376 7644 16440 7648
rect 16376 7588 16380 7644
rect 16380 7588 16436 7644
rect 16436 7588 16440 7644
rect 16376 7584 16440 7588
rect 16456 7644 16520 7648
rect 16456 7588 16460 7644
rect 16460 7588 16516 7644
rect 16516 7588 16520 7644
rect 16456 7584 16520 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 12216 7100 12280 7104
rect 12216 7044 12220 7100
rect 12220 7044 12276 7100
rect 12276 7044 12280 7100
rect 12216 7040 12280 7044
rect 12296 7100 12360 7104
rect 12296 7044 12300 7100
rect 12300 7044 12356 7100
rect 12356 7044 12360 7100
rect 12296 7040 12360 7044
rect 12376 7100 12440 7104
rect 12376 7044 12380 7100
rect 12380 7044 12436 7100
rect 12436 7044 12440 7100
rect 12376 7040 12440 7044
rect 12456 7100 12520 7104
rect 12456 7044 12460 7100
rect 12460 7044 12516 7100
rect 12516 7044 12520 7100
rect 12456 7040 12520 7044
rect 20216 7100 20280 7104
rect 20216 7044 20220 7100
rect 20220 7044 20276 7100
rect 20276 7044 20280 7100
rect 20216 7040 20280 7044
rect 20296 7100 20360 7104
rect 20296 7044 20300 7100
rect 20300 7044 20356 7100
rect 20356 7044 20360 7100
rect 20296 7040 20360 7044
rect 20376 7100 20440 7104
rect 20376 7044 20380 7100
rect 20380 7044 20436 7100
rect 20436 7044 20440 7100
rect 20376 7040 20440 7044
rect 20456 7100 20520 7104
rect 20456 7044 20460 7100
rect 20460 7044 20516 7100
rect 20516 7044 20520 7100
rect 20456 7040 20520 7044
rect 8216 6556 8280 6560
rect 8216 6500 8220 6556
rect 8220 6500 8276 6556
rect 8276 6500 8280 6556
rect 8216 6496 8280 6500
rect 8296 6556 8360 6560
rect 8296 6500 8300 6556
rect 8300 6500 8356 6556
rect 8356 6500 8360 6556
rect 8296 6496 8360 6500
rect 8376 6556 8440 6560
rect 8376 6500 8380 6556
rect 8380 6500 8436 6556
rect 8436 6500 8440 6556
rect 8376 6496 8440 6500
rect 8456 6556 8520 6560
rect 8456 6500 8460 6556
rect 8460 6500 8516 6556
rect 8516 6500 8520 6556
rect 8456 6496 8520 6500
rect 16216 6556 16280 6560
rect 16216 6500 16220 6556
rect 16220 6500 16276 6556
rect 16276 6500 16280 6556
rect 16216 6496 16280 6500
rect 16296 6556 16360 6560
rect 16296 6500 16300 6556
rect 16300 6500 16356 6556
rect 16356 6500 16360 6556
rect 16296 6496 16360 6500
rect 16376 6556 16440 6560
rect 16376 6500 16380 6556
rect 16380 6500 16436 6556
rect 16436 6500 16440 6556
rect 16376 6496 16440 6500
rect 16456 6556 16520 6560
rect 16456 6500 16460 6556
rect 16460 6500 16516 6556
rect 16516 6500 16520 6556
rect 16456 6496 16520 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 12216 6012 12280 6016
rect 12216 5956 12220 6012
rect 12220 5956 12276 6012
rect 12276 5956 12280 6012
rect 12216 5952 12280 5956
rect 12296 6012 12360 6016
rect 12296 5956 12300 6012
rect 12300 5956 12356 6012
rect 12356 5956 12360 6012
rect 12296 5952 12360 5956
rect 12376 6012 12440 6016
rect 12376 5956 12380 6012
rect 12380 5956 12436 6012
rect 12436 5956 12440 6012
rect 12376 5952 12440 5956
rect 12456 6012 12520 6016
rect 12456 5956 12460 6012
rect 12460 5956 12516 6012
rect 12516 5956 12520 6012
rect 12456 5952 12520 5956
rect 20216 6012 20280 6016
rect 20216 5956 20220 6012
rect 20220 5956 20276 6012
rect 20276 5956 20280 6012
rect 20216 5952 20280 5956
rect 20296 6012 20360 6016
rect 20296 5956 20300 6012
rect 20300 5956 20356 6012
rect 20356 5956 20360 6012
rect 20296 5952 20360 5956
rect 20376 6012 20440 6016
rect 20376 5956 20380 6012
rect 20380 5956 20436 6012
rect 20436 5956 20440 6012
rect 20376 5952 20440 5956
rect 20456 6012 20520 6016
rect 20456 5956 20460 6012
rect 20460 5956 20516 6012
rect 20516 5956 20520 6012
rect 20456 5952 20520 5956
rect 8216 5468 8280 5472
rect 8216 5412 8220 5468
rect 8220 5412 8276 5468
rect 8276 5412 8280 5468
rect 8216 5408 8280 5412
rect 8296 5468 8360 5472
rect 8296 5412 8300 5468
rect 8300 5412 8356 5468
rect 8356 5412 8360 5468
rect 8296 5408 8360 5412
rect 8376 5468 8440 5472
rect 8376 5412 8380 5468
rect 8380 5412 8436 5468
rect 8436 5412 8440 5468
rect 8376 5408 8440 5412
rect 8456 5468 8520 5472
rect 8456 5412 8460 5468
rect 8460 5412 8516 5468
rect 8516 5412 8520 5468
rect 8456 5408 8520 5412
rect 16216 5468 16280 5472
rect 16216 5412 16220 5468
rect 16220 5412 16276 5468
rect 16276 5412 16280 5468
rect 16216 5408 16280 5412
rect 16296 5468 16360 5472
rect 16296 5412 16300 5468
rect 16300 5412 16356 5468
rect 16356 5412 16360 5468
rect 16296 5408 16360 5412
rect 16376 5468 16440 5472
rect 16376 5412 16380 5468
rect 16380 5412 16436 5468
rect 16436 5412 16440 5468
rect 16376 5408 16440 5412
rect 16456 5468 16520 5472
rect 16456 5412 16460 5468
rect 16460 5412 16516 5468
rect 16516 5412 16520 5468
rect 16456 5408 16520 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 12216 4924 12280 4928
rect 12216 4868 12220 4924
rect 12220 4868 12276 4924
rect 12276 4868 12280 4924
rect 12216 4864 12280 4868
rect 12296 4924 12360 4928
rect 12296 4868 12300 4924
rect 12300 4868 12356 4924
rect 12356 4868 12360 4924
rect 12296 4864 12360 4868
rect 12376 4924 12440 4928
rect 12376 4868 12380 4924
rect 12380 4868 12436 4924
rect 12436 4868 12440 4924
rect 12376 4864 12440 4868
rect 12456 4924 12520 4928
rect 12456 4868 12460 4924
rect 12460 4868 12516 4924
rect 12516 4868 12520 4924
rect 12456 4864 12520 4868
rect 20216 4924 20280 4928
rect 20216 4868 20220 4924
rect 20220 4868 20276 4924
rect 20276 4868 20280 4924
rect 20216 4864 20280 4868
rect 20296 4924 20360 4928
rect 20296 4868 20300 4924
rect 20300 4868 20356 4924
rect 20356 4868 20360 4924
rect 20296 4864 20360 4868
rect 20376 4924 20440 4928
rect 20376 4868 20380 4924
rect 20380 4868 20436 4924
rect 20436 4868 20440 4924
rect 20376 4864 20440 4868
rect 20456 4924 20520 4928
rect 20456 4868 20460 4924
rect 20460 4868 20516 4924
rect 20516 4868 20520 4924
rect 20456 4864 20520 4868
rect 8216 4380 8280 4384
rect 8216 4324 8220 4380
rect 8220 4324 8276 4380
rect 8276 4324 8280 4380
rect 8216 4320 8280 4324
rect 8296 4380 8360 4384
rect 8296 4324 8300 4380
rect 8300 4324 8356 4380
rect 8356 4324 8360 4380
rect 8296 4320 8360 4324
rect 8376 4380 8440 4384
rect 8376 4324 8380 4380
rect 8380 4324 8436 4380
rect 8436 4324 8440 4380
rect 8376 4320 8440 4324
rect 8456 4380 8520 4384
rect 8456 4324 8460 4380
rect 8460 4324 8516 4380
rect 8516 4324 8520 4380
rect 8456 4320 8520 4324
rect 16216 4380 16280 4384
rect 16216 4324 16220 4380
rect 16220 4324 16276 4380
rect 16276 4324 16280 4380
rect 16216 4320 16280 4324
rect 16296 4380 16360 4384
rect 16296 4324 16300 4380
rect 16300 4324 16356 4380
rect 16356 4324 16360 4380
rect 16296 4320 16360 4324
rect 16376 4380 16440 4384
rect 16376 4324 16380 4380
rect 16380 4324 16436 4380
rect 16436 4324 16440 4380
rect 16376 4320 16440 4324
rect 16456 4380 16520 4384
rect 16456 4324 16460 4380
rect 16460 4324 16516 4380
rect 16516 4324 16520 4380
rect 16456 4320 16520 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 12216 3836 12280 3840
rect 12216 3780 12220 3836
rect 12220 3780 12276 3836
rect 12276 3780 12280 3836
rect 12216 3776 12280 3780
rect 12296 3836 12360 3840
rect 12296 3780 12300 3836
rect 12300 3780 12356 3836
rect 12356 3780 12360 3836
rect 12296 3776 12360 3780
rect 12376 3836 12440 3840
rect 12376 3780 12380 3836
rect 12380 3780 12436 3836
rect 12436 3780 12440 3836
rect 12376 3776 12440 3780
rect 12456 3836 12520 3840
rect 12456 3780 12460 3836
rect 12460 3780 12516 3836
rect 12516 3780 12520 3836
rect 12456 3776 12520 3780
rect 20216 3836 20280 3840
rect 20216 3780 20220 3836
rect 20220 3780 20276 3836
rect 20276 3780 20280 3836
rect 20216 3776 20280 3780
rect 20296 3836 20360 3840
rect 20296 3780 20300 3836
rect 20300 3780 20356 3836
rect 20356 3780 20360 3836
rect 20296 3776 20360 3780
rect 20376 3836 20440 3840
rect 20376 3780 20380 3836
rect 20380 3780 20436 3836
rect 20436 3780 20440 3836
rect 20376 3776 20440 3780
rect 20456 3836 20520 3840
rect 20456 3780 20460 3836
rect 20460 3780 20516 3836
rect 20516 3780 20520 3836
rect 20456 3776 20520 3780
rect 8216 3292 8280 3296
rect 8216 3236 8220 3292
rect 8220 3236 8276 3292
rect 8276 3236 8280 3292
rect 8216 3232 8280 3236
rect 8296 3292 8360 3296
rect 8296 3236 8300 3292
rect 8300 3236 8356 3292
rect 8356 3236 8360 3292
rect 8296 3232 8360 3236
rect 8376 3292 8440 3296
rect 8376 3236 8380 3292
rect 8380 3236 8436 3292
rect 8436 3236 8440 3292
rect 8376 3232 8440 3236
rect 8456 3292 8520 3296
rect 8456 3236 8460 3292
rect 8460 3236 8516 3292
rect 8516 3236 8520 3292
rect 8456 3232 8520 3236
rect 16216 3292 16280 3296
rect 16216 3236 16220 3292
rect 16220 3236 16276 3292
rect 16276 3236 16280 3292
rect 16216 3232 16280 3236
rect 16296 3292 16360 3296
rect 16296 3236 16300 3292
rect 16300 3236 16356 3292
rect 16356 3236 16360 3292
rect 16296 3232 16360 3236
rect 16376 3292 16440 3296
rect 16376 3236 16380 3292
rect 16380 3236 16436 3292
rect 16436 3236 16440 3292
rect 16376 3232 16440 3236
rect 16456 3292 16520 3296
rect 16456 3236 16460 3292
rect 16460 3236 16516 3292
rect 16516 3236 16520 3292
rect 16456 3232 16520 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 12216 2748 12280 2752
rect 12216 2692 12220 2748
rect 12220 2692 12276 2748
rect 12276 2692 12280 2748
rect 12216 2688 12280 2692
rect 12296 2748 12360 2752
rect 12296 2692 12300 2748
rect 12300 2692 12356 2748
rect 12356 2692 12360 2748
rect 12296 2688 12360 2692
rect 12376 2748 12440 2752
rect 12376 2692 12380 2748
rect 12380 2692 12436 2748
rect 12436 2692 12440 2748
rect 12376 2688 12440 2692
rect 12456 2748 12520 2752
rect 12456 2692 12460 2748
rect 12460 2692 12516 2748
rect 12516 2692 12520 2748
rect 12456 2688 12520 2692
rect 20216 2748 20280 2752
rect 20216 2692 20220 2748
rect 20220 2692 20276 2748
rect 20276 2692 20280 2748
rect 20216 2688 20280 2692
rect 20296 2748 20360 2752
rect 20296 2692 20300 2748
rect 20300 2692 20356 2748
rect 20356 2692 20360 2748
rect 20296 2688 20360 2692
rect 20376 2748 20440 2752
rect 20376 2692 20380 2748
rect 20380 2692 20436 2748
rect 20436 2692 20440 2748
rect 20376 2688 20440 2692
rect 20456 2748 20520 2752
rect 20456 2692 20460 2748
rect 20460 2692 20516 2748
rect 20516 2692 20520 2748
rect 20456 2688 20520 2692
rect 8216 2204 8280 2208
rect 8216 2148 8220 2204
rect 8220 2148 8276 2204
rect 8276 2148 8280 2204
rect 8216 2144 8280 2148
rect 8296 2204 8360 2208
rect 8296 2148 8300 2204
rect 8300 2148 8356 2204
rect 8356 2148 8360 2204
rect 8296 2144 8360 2148
rect 8376 2204 8440 2208
rect 8376 2148 8380 2204
rect 8380 2148 8436 2204
rect 8436 2148 8440 2204
rect 8376 2144 8440 2148
rect 8456 2204 8520 2208
rect 8456 2148 8460 2204
rect 8460 2148 8516 2204
rect 8516 2148 8520 2204
rect 8456 2144 8520 2148
rect 16216 2204 16280 2208
rect 16216 2148 16220 2204
rect 16220 2148 16276 2204
rect 16276 2148 16280 2204
rect 16216 2144 16280 2148
rect 16296 2204 16360 2208
rect 16296 2148 16300 2204
rect 16300 2148 16356 2204
rect 16356 2148 16360 2204
rect 16296 2144 16360 2148
rect 16376 2204 16440 2208
rect 16376 2148 16380 2204
rect 16380 2148 16436 2204
rect 16436 2148 16440 2204
rect 16376 2144 16440 2148
rect 16456 2204 16520 2208
rect 16456 2148 16460 2204
rect 16460 2148 16516 2204
rect 16516 2148 16520 2204
rect 16456 2144 16520 2148
rect 4216 1660 4280 1664
rect 4216 1604 4220 1660
rect 4220 1604 4276 1660
rect 4276 1604 4280 1660
rect 4216 1600 4280 1604
rect 4296 1660 4360 1664
rect 4296 1604 4300 1660
rect 4300 1604 4356 1660
rect 4356 1604 4360 1660
rect 4296 1600 4360 1604
rect 4376 1660 4440 1664
rect 4376 1604 4380 1660
rect 4380 1604 4436 1660
rect 4436 1604 4440 1660
rect 4376 1600 4440 1604
rect 4456 1660 4520 1664
rect 4456 1604 4460 1660
rect 4460 1604 4516 1660
rect 4516 1604 4520 1660
rect 4456 1600 4520 1604
rect 12216 1660 12280 1664
rect 12216 1604 12220 1660
rect 12220 1604 12276 1660
rect 12276 1604 12280 1660
rect 12216 1600 12280 1604
rect 12296 1660 12360 1664
rect 12296 1604 12300 1660
rect 12300 1604 12356 1660
rect 12356 1604 12360 1660
rect 12296 1600 12360 1604
rect 12376 1660 12440 1664
rect 12376 1604 12380 1660
rect 12380 1604 12436 1660
rect 12436 1604 12440 1660
rect 12376 1600 12440 1604
rect 12456 1660 12520 1664
rect 12456 1604 12460 1660
rect 12460 1604 12516 1660
rect 12516 1604 12520 1660
rect 12456 1600 12520 1604
rect 20216 1660 20280 1664
rect 20216 1604 20220 1660
rect 20220 1604 20276 1660
rect 20276 1604 20280 1660
rect 20216 1600 20280 1604
rect 20296 1660 20360 1664
rect 20296 1604 20300 1660
rect 20300 1604 20356 1660
rect 20356 1604 20360 1660
rect 20296 1600 20360 1604
rect 20376 1660 20440 1664
rect 20376 1604 20380 1660
rect 20380 1604 20436 1660
rect 20436 1604 20440 1660
rect 20376 1600 20440 1604
rect 20456 1660 20520 1664
rect 20456 1604 20460 1660
rect 20460 1604 20516 1660
rect 20516 1604 20520 1660
rect 20456 1600 20520 1604
rect 8216 1116 8280 1120
rect 8216 1060 8220 1116
rect 8220 1060 8276 1116
rect 8276 1060 8280 1116
rect 8216 1056 8280 1060
rect 8296 1116 8360 1120
rect 8296 1060 8300 1116
rect 8300 1060 8356 1116
rect 8356 1060 8360 1116
rect 8296 1056 8360 1060
rect 8376 1116 8440 1120
rect 8376 1060 8380 1116
rect 8380 1060 8436 1116
rect 8436 1060 8440 1116
rect 8376 1056 8440 1060
rect 8456 1116 8520 1120
rect 8456 1060 8460 1116
rect 8460 1060 8516 1116
rect 8516 1060 8520 1116
rect 8456 1056 8520 1060
rect 16216 1116 16280 1120
rect 16216 1060 16220 1116
rect 16220 1060 16276 1116
rect 16276 1060 16280 1116
rect 16216 1056 16280 1060
rect 16296 1116 16360 1120
rect 16296 1060 16300 1116
rect 16300 1060 16356 1116
rect 16356 1060 16360 1116
rect 16296 1056 16360 1060
rect 16376 1116 16440 1120
rect 16376 1060 16380 1116
rect 16380 1060 16436 1116
rect 16436 1060 16440 1116
rect 16376 1056 16440 1060
rect 16456 1116 16520 1120
rect 16456 1060 16460 1116
rect 16460 1060 16516 1116
rect 16516 1060 16520 1116
rect 16456 1056 16520 1060
<< metal4 >>
rect 4208 13632 4528 13648
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 1664 4528 2688
rect 4208 1600 4216 1664
rect 4280 1600 4296 1664
rect 4360 1600 4376 1664
rect 4440 1600 4456 1664
rect 4520 1600 4528 1664
rect 4208 1040 4528 1600
rect 8208 13088 8528 13648
rect 8208 13024 8216 13088
rect 8280 13024 8296 13088
rect 8360 13024 8376 13088
rect 8440 13024 8456 13088
rect 8520 13024 8528 13088
rect 8208 12000 8528 13024
rect 8208 11936 8216 12000
rect 8280 11936 8296 12000
rect 8360 11936 8376 12000
rect 8440 11936 8456 12000
rect 8520 11936 8528 12000
rect 8208 10912 8528 11936
rect 8208 10848 8216 10912
rect 8280 10848 8296 10912
rect 8360 10848 8376 10912
rect 8440 10848 8456 10912
rect 8520 10848 8528 10912
rect 8208 9824 8528 10848
rect 8208 9760 8216 9824
rect 8280 9760 8296 9824
rect 8360 9760 8376 9824
rect 8440 9760 8456 9824
rect 8520 9760 8528 9824
rect 8208 8736 8528 9760
rect 8208 8672 8216 8736
rect 8280 8672 8296 8736
rect 8360 8672 8376 8736
rect 8440 8672 8456 8736
rect 8520 8672 8528 8736
rect 8208 7648 8528 8672
rect 8208 7584 8216 7648
rect 8280 7584 8296 7648
rect 8360 7584 8376 7648
rect 8440 7584 8456 7648
rect 8520 7584 8528 7648
rect 8208 6560 8528 7584
rect 8208 6496 8216 6560
rect 8280 6496 8296 6560
rect 8360 6496 8376 6560
rect 8440 6496 8456 6560
rect 8520 6496 8528 6560
rect 8208 5472 8528 6496
rect 8208 5408 8216 5472
rect 8280 5408 8296 5472
rect 8360 5408 8376 5472
rect 8440 5408 8456 5472
rect 8520 5408 8528 5472
rect 8208 4384 8528 5408
rect 8208 4320 8216 4384
rect 8280 4320 8296 4384
rect 8360 4320 8376 4384
rect 8440 4320 8456 4384
rect 8520 4320 8528 4384
rect 8208 3296 8528 4320
rect 8208 3232 8216 3296
rect 8280 3232 8296 3296
rect 8360 3232 8376 3296
rect 8440 3232 8456 3296
rect 8520 3232 8528 3296
rect 8208 2208 8528 3232
rect 8208 2144 8216 2208
rect 8280 2144 8296 2208
rect 8360 2144 8376 2208
rect 8440 2144 8456 2208
rect 8520 2144 8528 2208
rect 8208 1120 8528 2144
rect 8208 1056 8216 1120
rect 8280 1056 8296 1120
rect 8360 1056 8376 1120
rect 8440 1056 8456 1120
rect 8520 1056 8528 1120
rect 8208 1040 8528 1056
rect 12208 13632 12528 13648
rect 12208 13568 12216 13632
rect 12280 13568 12296 13632
rect 12360 13568 12376 13632
rect 12440 13568 12456 13632
rect 12520 13568 12528 13632
rect 12208 12544 12528 13568
rect 12208 12480 12216 12544
rect 12280 12480 12296 12544
rect 12360 12480 12376 12544
rect 12440 12480 12456 12544
rect 12520 12480 12528 12544
rect 12208 11456 12528 12480
rect 12208 11392 12216 11456
rect 12280 11392 12296 11456
rect 12360 11392 12376 11456
rect 12440 11392 12456 11456
rect 12520 11392 12528 11456
rect 12208 10368 12528 11392
rect 12208 10304 12216 10368
rect 12280 10304 12296 10368
rect 12360 10304 12376 10368
rect 12440 10304 12456 10368
rect 12520 10304 12528 10368
rect 12208 9280 12528 10304
rect 12208 9216 12216 9280
rect 12280 9216 12296 9280
rect 12360 9216 12376 9280
rect 12440 9216 12456 9280
rect 12520 9216 12528 9280
rect 12208 8192 12528 9216
rect 12208 8128 12216 8192
rect 12280 8128 12296 8192
rect 12360 8128 12376 8192
rect 12440 8128 12456 8192
rect 12520 8128 12528 8192
rect 12208 7104 12528 8128
rect 12208 7040 12216 7104
rect 12280 7040 12296 7104
rect 12360 7040 12376 7104
rect 12440 7040 12456 7104
rect 12520 7040 12528 7104
rect 12208 6016 12528 7040
rect 12208 5952 12216 6016
rect 12280 5952 12296 6016
rect 12360 5952 12376 6016
rect 12440 5952 12456 6016
rect 12520 5952 12528 6016
rect 12208 4928 12528 5952
rect 12208 4864 12216 4928
rect 12280 4864 12296 4928
rect 12360 4864 12376 4928
rect 12440 4864 12456 4928
rect 12520 4864 12528 4928
rect 12208 3840 12528 4864
rect 12208 3776 12216 3840
rect 12280 3776 12296 3840
rect 12360 3776 12376 3840
rect 12440 3776 12456 3840
rect 12520 3776 12528 3840
rect 12208 2752 12528 3776
rect 12208 2688 12216 2752
rect 12280 2688 12296 2752
rect 12360 2688 12376 2752
rect 12440 2688 12456 2752
rect 12520 2688 12528 2752
rect 12208 1664 12528 2688
rect 12208 1600 12216 1664
rect 12280 1600 12296 1664
rect 12360 1600 12376 1664
rect 12440 1600 12456 1664
rect 12520 1600 12528 1664
rect 12208 1040 12528 1600
rect 16208 13088 16528 13648
rect 16208 13024 16216 13088
rect 16280 13024 16296 13088
rect 16360 13024 16376 13088
rect 16440 13024 16456 13088
rect 16520 13024 16528 13088
rect 16208 12000 16528 13024
rect 16208 11936 16216 12000
rect 16280 11936 16296 12000
rect 16360 11936 16376 12000
rect 16440 11936 16456 12000
rect 16520 11936 16528 12000
rect 16208 10912 16528 11936
rect 16208 10848 16216 10912
rect 16280 10848 16296 10912
rect 16360 10848 16376 10912
rect 16440 10848 16456 10912
rect 16520 10848 16528 10912
rect 16208 9824 16528 10848
rect 16208 9760 16216 9824
rect 16280 9760 16296 9824
rect 16360 9760 16376 9824
rect 16440 9760 16456 9824
rect 16520 9760 16528 9824
rect 16208 8736 16528 9760
rect 16208 8672 16216 8736
rect 16280 8672 16296 8736
rect 16360 8672 16376 8736
rect 16440 8672 16456 8736
rect 16520 8672 16528 8736
rect 16208 7648 16528 8672
rect 16208 7584 16216 7648
rect 16280 7584 16296 7648
rect 16360 7584 16376 7648
rect 16440 7584 16456 7648
rect 16520 7584 16528 7648
rect 16208 6560 16528 7584
rect 16208 6496 16216 6560
rect 16280 6496 16296 6560
rect 16360 6496 16376 6560
rect 16440 6496 16456 6560
rect 16520 6496 16528 6560
rect 16208 5472 16528 6496
rect 16208 5408 16216 5472
rect 16280 5408 16296 5472
rect 16360 5408 16376 5472
rect 16440 5408 16456 5472
rect 16520 5408 16528 5472
rect 16208 4384 16528 5408
rect 16208 4320 16216 4384
rect 16280 4320 16296 4384
rect 16360 4320 16376 4384
rect 16440 4320 16456 4384
rect 16520 4320 16528 4384
rect 16208 3296 16528 4320
rect 16208 3232 16216 3296
rect 16280 3232 16296 3296
rect 16360 3232 16376 3296
rect 16440 3232 16456 3296
rect 16520 3232 16528 3296
rect 16208 2208 16528 3232
rect 16208 2144 16216 2208
rect 16280 2144 16296 2208
rect 16360 2144 16376 2208
rect 16440 2144 16456 2208
rect 16520 2144 16528 2208
rect 16208 1120 16528 2144
rect 16208 1056 16216 1120
rect 16280 1056 16296 1120
rect 16360 1056 16376 1120
rect 16440 1056 16456 1120
rect 16520 1056 16528 1120
rect 16208 1040 16528 1056
rect 20208 13632 20528 13648
rect 20208 13568 20216 13632
rect 20280 13568 20296 13632
rect 20360 13568 20376 13632
rect 20440 13568 20456 13632
rect 20520 13568 20528 13632
rect 20208 12544 20528 13568
rect 20208 12480 20216 12544
rect 20280 12480 20296 12544
rect 20360 12480 20376 12544
rect 20440 12480 20456 12544
rect 20520 12480 20528 12544
rect 20208 11456 20528 12480
rect 20208 11392 20216 11456
rect 20280 11392 20296 11456
rect 20360 11392 20376 11456
rect 20440 11392 20456 11456
rect 20520 11392 20528 11456
rect 20208 10368 20528 11392
rect 20208 10304 20216 10368
rect 20280 10304 20296 10368
rect 20360 10304 20376 10368
rect 20440 10304 20456 10368
rect 20520 10304 20528 10368
rect 20208 9280 20528 10304
rect 20208 9216 20216 9280
rect 20280 9216 20296 9280
rect 20360 9216 20376 9280
rect 20440 9216 20456 9280
rect 20520 9216 20528 9280
rect 20208 8192 20528 9216
rect 20208 8128 20216 8192
rect 20280 8128 20296 8192
rect 20360 8128 20376 8192
rect 20440 8128 20456 8192
rect 20520 8128 20528 8192
rect 20208 7104 20528 8128
rect 20208 7040 20216 7104
rect 20280 7040 20296 7104
rect 20360 7040 20376 7104
rect 20440 7040 20456 7104
rect 20520 7040 20528 7104
rect 20208 6016 20528 7040
rect 20208 5952 20216 6016
rect 20280 5952 20296 6016
rect 20360 5952 20376 6016
rect 20440 5952 20456 6016
rect 20520 5952 20528 6016
rect 20208 4928 20528 5952
rect 20208 4864 20216 4928
rect 20280 4864 20296 4928
rect 20360 4864 20376 4928
rect 20440 4864 20456 4928
rect 20520 4864 20528 4928
rect 20208 3840 20528 4864
rect 20208 3776 20216 3840
rect 20280 3776 20296 3840
rect 20360 3776 20376 3840
rect 20440 3776 20456 3840
rect 20520 3776 20528 3840
rect 20208 2752 20528 3776
rect 20208 2688 20216 2752
rect 20280 2688 20296 2752
rect 20360 2688 20376 2752
rect 20440 2688 20456 2752
rect 20520 2688 20528 2752
rect 20208 1664 20528 2688
rect 20208 1600 20216 1664
rect 20280 1600 20296 1664
rect 20360 1600 20376 1664
rect 20440 1600 20456 1664
rect 20520 1600 20528 1664
rect 20208 1040 20528 1600
use sky130_fd_sc_hd__xnor2_2  _096_
timestamp 21601
transform -1 0 7544 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _097_
timestamp 21601
transform -1 0 10120 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_2  _098_
timestamp 21601
transform 1 0 12144 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _099_
timestamp 21601
transform 1 0 12236 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _100_
timestamp 21601
transform -1 0 11316 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _101_
timestamp 21601
transform -1 0 15272 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _102_
timestamp 21601
transform -1 0 21712 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _103_
timestamp 21601
transform -1 0 5888 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_2  _104_
timestamp 21601
transform -1 0 7084 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _105_
timestamp 21601
transform 1 0 6624 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _106_
timestamp 21601
transform -1 0 6256 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _107_
timestamp 21601
transform -1 0 8464 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _108_
timestamp 1562557784
transform -1 0 3680 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _109_
timestamp 1562557784
transform -1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _110_
timestamp 21601
transform -1 0 4508 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _111_
timestamp 1562557784
transform -1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _112_
timestamp 1562557784
transform 1 0 7820 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _113_
timestamp 21601
transform -1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _114_
timestamp 21601
transform 1 0 2852 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _115_
timestamp 21601
transform 1 0 3588 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _116_
timestamp 21601
transform 1 0 4140 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _117_
timestamp 21601
transform 1 0 3956 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _118_
timestamp 1562557784
transform 1 0 4048 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _119_
timestamp 1562557784
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1562557784
transform -1 0 4232 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _121_
timestamp 21601
transform -1 0 11132 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _122_
timestamp 1562557784
transform -1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _123_
timestamp 21601
transform 1 0 9752 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _124_
timestamp 21601
transform 1 0 5520 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _125_
timestamp 21601
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _126_
timestamp 21601
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _127_
timestamp 21601
transform 1 0 10488 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _128_
timestamp 21601
transform 1 0 11500 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _129_
timestamp 1562557784
transform -1 0 1748 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _130_
timestamp 21601
transform 1 0 6900 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _131_
timestamp 21601
transform -1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _132_
timestamp 21601
transform 1 0 2484 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _133_
timestamp 21601
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _134_
timestamp 21601
transform 1 0 4784 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _135_
timestamp 1562557784
transform 1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136_
timestamp 1562557784
transform -1 0 7728 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _137_
timestamp 1562557784
transform -1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _138_
timestamp 1562557784
transform -1 0 5152 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _139_
timestamp 1562557784
transform 1 0 7268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _140_
timestamp 1562557784
transform 1 0 10304 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _141_
timestamp 1562557784
transform 1 0 11592 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142_
timestamp 1562557784
transform -1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1562557784
transform -1 0 14352 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _144_
timestamp 1562557784
transform 1 0 1472 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _145_
timestamp 1562557784
transform 1 0 3312 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _146_
timestamp 1562557784
transform 1 0 8924 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _147_
timestamp 1562557784
transform 1 0 11040 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148_
timestamp 1562557784
transform -1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _149_
timestamp 1562557784
transform 1 0 14536 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _150_
timestamp 1562557784
transform 1 0 12696 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _151_
timestamp 1562557784
transform 1 0 17572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _152_
timestamp 1562557784
transform -1 0 15548 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _153_
timestamp 1562557784
transform 1 0 11132 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154_
timestamp 1562557784
transform -1 0 3588 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _155_
timestamp 1562557784
transform 1 0 5244 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _156_
timestamp 1562557784
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _157_
timestamp 1562557784
transform -1 0 15824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _158_
timestamp 21601
transform -1 0 12052 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_2  _159_
timestamp 21601
transform 1 0 9016 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _160_
timestamp 1562557784
transform -1 0 12420 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _161_
timestamp 21601
transform -1 0 15272 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _162_
timestamp 1562557784
transform 1 0 12972 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _163_
timestamp 21601
transform 1 0 12420 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _164_
timestamp 1562557784
transform 1 0 16100 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _165_
timestamp 21601
transform -1 0 12788 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _166_
timestamp 21601
transform -1 0 12144 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _167_
timestamp 21601
transform -1 0 9476 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _168_
timestamp 21601
transform 1 0 9752 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _169_
timestamp 21601
transform -1 0 11408 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _170_
timestamp 21601
transform -1 0 12052 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _171_
timestamp 21601
transform -1 0 13432 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _172_
timestamp 21601
transform 1 0 13432 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _173_
timestamp 21601
transform 1 0 15364 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _174_
timestamp 21601
transform 1 0 6348 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _175_
timestamp 21601
transform -1 0 6808 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _176_
timestamp 21601
transform -1 0 4140 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _177_
timestamp 1562557784
transform 1 0 3496 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _178_
timestamp 21601
transform -1 0 2116 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _179_
timestamp 21601
transform 1 0 5704 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _180_
timestamp 21601
transform -1 0 3496 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _181_
timestamp 1562557784
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _182_
timestamp 21601
transform -1 0 2116 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _183_
timestamp 21601
transform 1 0 5796 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _184_
timestamp 21601
transform -1 0 2576 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _185_
timestamp 1562557784
transform 1 0 1472 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _186_
timestamp 21601
transform 1 0 2944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _187_
timestamp 1562557784
transform -1 0 5980 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _188_
timestamp 21601
transform -1 0 1840 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _189_
timestamp 21601
transform 1 0 3772 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _190_
timestamp 21601
transform 1 0 7084 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _191_
timestamp 1562557784
transform -1 0 6716 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _192_
timestamp 21601
transform 1 0 8188 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _193_
timestamp 21601
transform -1 0 6532 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _194_
timestamp 21601
transform -1 0 10120 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _195_
timestamp 21601
transform 1 0 10120 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _196_
timestamp 21601
transform -1 0 10120 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _197_
timestamp 1562557784
transform 1 0 10580 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _198_
timestamp 21601
transform 1 0 8280 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _199_
timestamp 21601
transform -1 0 7176 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _200_
timestamp 21601
transform -1 0 8096 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_2  _201_
timestamp 21601
transform -1 0 2760 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _202_
timestamp 21601
transform 1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _203_
timestamp 21601
transform 1 0 6348 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _204_
timestamp 1562557784
transform 1 0 10304 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _205_
timestamp 21601
transform -1 0 9568 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _206_
timestamp 21601
transform 1 0 4508 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _207_
timestamp 21601
transform -1 0 8740 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1562557784
transform -1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _209_
timestamp 21601
transform -1 0 2024 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _210_
timestamp 21601
transform 1 0 2484 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _211_
timestamp 21601
transform 1 0 9660 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _212_
timestamp 1562557784
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _213_
timestamp 21601
transform 1 0 13156 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _214_
timestamp 21601
transform -1 0 11960 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _215_
timestamp 21601
transform 1 0 12696 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _216_
timestamp 21601
transform 1 0 10488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _217_
timestamp 1562557784
transform 1 0 15364 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _218_
timestamp 21601
transform 1 0 11500 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _219_
timestamp 21601
transform -1 0 6900 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _220_
timestamp 21601
transform -1 0 16376 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _221_
timestamp 21601
transform 1 0 16652 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _222_
timestamp 21601
transform -1 0 16560 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _223_
timestamp 1562557784
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _224_
timestamp 21601
transform 1 0 15732 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _225_
timestamp 21601
transform -1 0 13984 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _226_
timestamp 21601
transform -1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _227_
timestamp 21601
transform 1 0 11776 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _228_
timestamp 21601
transform -1 0 11132 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _229_
timestamp 21601
transform -1 0 10672 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _230_
timestamp 21601
transform 1 0 3772 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _231_
timestamp 1562557784
transform -1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _232_
timestamp 21601
transform -1 0 2208 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _233_
timestamp 21601
transform -1 0 3220 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _234_
timestamp 21601
transform 1 0 8188 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _235_
timestamp 21601
transform -1 0 6808 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _236_
timestamp 21601
transform -1 0 6256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _237_
timestamp 1562557784
transform 1 0 6532 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _238_
timestamp 21601
transform -1 0 6256 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _239_
timestamp 21601
transform -1 0 5612 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_2  _240_
timestamp 21601
transform 1 0 6808 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _241_
timestamp 21601
transform 1 0 1564 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_2  _242_
timestamp 21601
transform 1 0 3772 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _243_
timestamp 21601
transform 1 0 3864 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _244_
timestamp 21601
transform -1 0 4968 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _245_
timestamp 21601
transform 1 0 14076 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _246_
timestamp 21601
transform 1 0 19780 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _247_
timestamp 21601
transform 1 0 20240 0 1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _248_
timestamp 21601
transform 1 0 9476 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _249_
timestamp 21601
transform 1 0 11500 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _250_
timestamp 21601
transform -1 0 13984 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _251_
timestamp 21601
transform 1 0 12052 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _252_
timestamp 21601
transform 1 0 11776 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _253_
timestamp 21601
transform 1 0 13340 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _254_
timestamp 21601
transform 1 0 10120 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _255_
timestamp 21601
transform -1 0 8740 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _256_
timestamp 21601
transform -1 0 11408 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _257_
timestamp 21601
transform 1 0 7544 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _258_
timestamp 21601
transform 1 0 6900 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _259_
timestamp 21601
transform 1 0 10672 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _260_
timestamp 21601
transform 1 0 14076 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _261_
timestamp 21601
transform 1 0 11868 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _262_
timestamp 21601
transform 1 0 12052 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _263_
timestamp 21601
transform 1 0 12052 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _264_
timestamp 21601
transform 1 0 16008 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _265_
timestamp 21601
transform 1 0 14076 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _266_
timestamp 21601
transform 1 0 13432 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _267_
timestamp 21601
transform -1 0 5704 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _268_
timestamp 21601
transform 1 0 2116 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _269_
timestamp 21601
transform 1 0 4324 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _270_
timestamp 21601
transform -1 0 3312 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _271_
timestamp 21601
transform 1 0 1748 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _272_
timestamp 21601
transform 1 0 1748 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _273_
timestamp 21601
transform 1 0 3864 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _274_
timestamp 21601
transform -1 0 3404 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _275_
timestamp 21601
transform 1 0 1748 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _276_
timestamp 21601
transform 1 0 1748 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _277_
timestamp 21601
transform 1 0 3772 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _278_
timestamp 21601
transform -1 0 3312 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _279_
timestamp 21601
transform 1 0 1380 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _280_
timestamp 21601
transform 1 0 4416 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _281_
timestamp 21601
transform 1 0 1748 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _282_
timestamp 21601
transform 1 0 3588 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _283_
timestamp 21601
transform 1 0 8372 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _284_
timestamp 21601
transform 1 0 7084 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _285_
timestamp 21601
transform 1 0 9200 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _286_
timestamp 21601
transform 1 0 5980 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _287_
timestamp 21601
transform 1 0 9384 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _288_
timestamp 21601
transform 1 0 11592 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _289_
timestamp 21601
transform 1 0 10120 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _290_
timestamp 21601
transform 1 0 10396 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _291_
timestamp 21601
transform 1 0 8188 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _292_
timestamp 21601
transform 1 0 6440 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _293_
timestamp 21601
transform -1 0 11500 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _294_
timestamp 21601
transform 1 0 6348 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _295_
timestamp 21601
transform 1 0 1748 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _296_
timestamp 21601
transform 1 0 3772 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _297_
timestamp 21601
transform 1 0 4324 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _298_
timestamp 21601
transform 1 0 5336 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _299_
timestamp 21601
transform 1 0 7452 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _300_
timestamp 21601
transform 1 0 3864 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _301_
timestamp 21601
transform 1 0 6440 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _302_
timestamp 21601
transform 1 0 4968 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _303_
timestamp 21601
transform 1 0 4324 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _304_
timestamp 21601
transform 1 0 6900 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _305_
timestamp 21601
transform -1 0 10304 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _306_
timestamp 21601
transform 1 0 9476 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _307_
timestamp 21601
transform 1 0 6440 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _308_
timestamp 21601
transform 1 0 1748 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _309_
timestamp 21601
transform 1 0 3680 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _310_
timestamp 21601
transform 1 0 3956 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _311_
timestamp 21601
transform 1 0 2024 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _312_
timestamp 21601
transform -1 0 11224 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _313_
timestamp 21601
transform -1 0 16100 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _314_
timestamp 21601
transform 1 0 11224 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _315_
timestamp 21601
transform 1 0 13064 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _316_
timestamp 21601
transform 1 0 9476 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _317_
timestamp 21601
transform 1 0 8924 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _318_
timestamp 21601
transform -1 0 13432 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _319_
timestamp 21601
transform 1 0 6900 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _320_
timestamp 21601
transform 1 0 15640 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _321_
timestamp 21601
transform -1 0 19504 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _322_
timestamp 21601
transform 1 0 14536 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _323_
timestamp 21601
transform 1 0 16652 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _324_
timestamp 21601
transform 1 0 16192 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _325_
timestamp 21601
transform 1 0 14260 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _326_
timestamp 21601
transform -1 0 18860 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _327_
timestamp 21601
transform 1 0 13156 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _328_
timestamp 21601
transform 1 0 11500 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _329_
timestamp 21601
transform 1 0 6348 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _330_
timestamp 21601
transform 1 0 8464 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _331_
timestamp 21601
transform 1 0 11316 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _332_
timestamp 21601
transform 1 0 12972 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _333_
timestamp 21601
transform -1 0 10856 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _334_
timestamp 21601
transform 1 0 11500 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _335_
timestamp 21601
transform 1 0 10856 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _336_
timestamp 21601
transform 1 0 9476 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _337_
timestamp 21601
transform 1 0 1748 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _338_
timestamp 21601
transform 1 0 2208 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _339_
timestamp 21601
transform 1 0 3312 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _340_
timestamp 21601
transform -1 0 3312 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _341_
timestamp 21601
transform 1 0 6900 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _342_
timestamp 21601
transform 1 0 6256 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _343_
timestamp 21601
transform -1 0 9660 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _344_
timestamp 21601
transform 1 0 4968 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _345_
timestamp 21601
transform 1 0 6808 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _346_
timestamp 21601
transform 1 0 4324 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _347_
timestamp 21601
transform 1 0 7636 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _348_
timestamp 21601
transform -1 0 6256 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _349_
timestamp 21601
transform 1 0 7544 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _350_
timestamp 21601
transform 1 0 1932 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _351_
timestamp 21601
transform -1 0 3680 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _352_
timestamp 21601
transform 1 0 4140 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _353_
timestamp 21601
transform 1 0 5520 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _354_
timestamp 1562557784
transform 1 0 10580 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _355_
timestamp 21601
transform -1 0 22172 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_12  _356_
timestamp 21601
transform 1 0 16744 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  _357_
timestamp 21601
transform 1 0 21068 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  _358_
timestamp 21601
transform 1 0 18584 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  _359_
timestamp 21601
transform 1 0 20240 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  _360_
timestamp 21601
transform 1 0 14904 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  _361_
timestamp 21601
transform 1 0 14076 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__clkbuf_8  clk_div1_delay.dly_clkbuf
timestamp 21601
transform 1 0 16652 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[1\].dlygen
timestamp 21601
transform -1 0 13800 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[2\].dlygen
timestamp 21601
transform 1 0 13432 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[3\].dlygen
timestamp 21601
transform 1 0 14168 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[4\].dlygen
timestamp 21601
transform -1 0 14812 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[5\].dlygen
timestamp 21601
transform 1 0 14904 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[6\].dlygen
timestamp 21601
transform -1 0 15548 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[7\].dlygen
timestamp 21601
transform 1 0 15640 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  clk_div1_delay.gen_dlygen\[8\].dlygen
timestamp 21601
transform -1 0 16284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  fanout1
timestamp 21601
transform -1 0 6808 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  fanout2
timestamp 21601
transform 1 0 12604 0 1 2176
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_1  fanout3
timestamp 21601
transform -1 0 10672 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  fanout4
timestamp 21601
transform 1 0 10396 0 -1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_12  fanout5
timestamp 21601
transform 1 0 13708 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  fanout6
timestamp 21601
transform 1 0 15088 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  fanout7
timestamp 21601
transform -1 0 13892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24
timestamp 21601
transform 1 0 3312 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 21601
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 21601
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 21601
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_134
timestamp 21601
transform 1 0 13432 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 21601
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_149
timestamp 21601
transform 1 0 14812 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 21601
transform 1 0 15088 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_155
timestamp 21601
transform 1 0 15364 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_158
timestamp 21601
transform 1 0 15640 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_161
timestamp 21601
transform 1 0 15916 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_164
timestamp 21601
transform 1 0 16192 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 21601
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 21601
transform 1 0 16652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_172
timestamp 21601
transform 1 0 16928 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_175
timestamp 21601
transform 1 0 17204 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_178
timestamp 21601
transform 1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_181
timestamp 21601
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_184
timestamp 21601
transform 1 0 18032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 21601
transform 1 0 18308 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_190
timestamp 21601
transform 1 0 18584 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_193
timestamp 21601
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_197
timestamp 21601
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_200
timestamp 21601
transform 1 0 19504 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_203
timestamp 21601
transform 1 0 19780 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_206
timestamp 21601
transform 1 0 20056 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_209
timestamp 21601
transform 1 0 20332 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_212
timestamp 21601
transform 1 0 20608 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_215
timestamp 21601
transform 1 0 20884 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 21601
transform 1 0 21160 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 21601
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_225
timestamp 21601
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_228
timestamp 21601
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_231
timestamp 21601
transform 1 0 22356 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 21601
transform 1 0 1380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_65
timestamp 21601
transform 1 0 7084 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_148
timestamp 21601
transform 1 0 14720 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 21601
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 21601
transform 1 0 16652 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_186
timestamp 21601
transform 1 0 18216 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 21601
transform 1 0 18492 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_206
timestamp 21601
transform 1 0 20056 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_229
timestamp 21601
transform 1 0 22172 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_232
timestamp 21601
transform 1 0 22448 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_3
timestamp 21601
transform 1 0 1380 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 21601
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_62
timestamp 21601
transform 1 0 6808 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 21601
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 21601
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_157
timestamp 21601
transform 1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_160
timestamp 21601
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_163
timestamp 21601
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_166
timestamp 21601
transform 1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_169
timestamp 21601
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_172
timestamp 21601
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_175
timestamp 21601
transform 1 0 17204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_178
timestamp 21601
transform 1 0 17480 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_181
timestamp 21601
transform 1 0 17756 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_184
timestamp 21601
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_187
timestamp 21601
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_190
timestamp 21601
transform 1 0 18584 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_193
timestamp 21601
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_197
timestamp 21601
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_200
timestamp 21601
transform 1 0 19504 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_203
timestamp 21601
transform 1 0 19780 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_206
timestamp 21601
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_209
timestamp 21601
transform 1 0 20332 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_212
timestamp 21601
transform 1 0 20608 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_215
timestamp 21601
transform 1 0 20884 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_3
timestamp 21601
transform 1 0 1380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_33
timestamp 21601
transform 1 0 4140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 21601
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_106
timestamp 21601
transform 1 0 10856 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 21601
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_154
timestamp 21601
transform 1 0 15272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_157
timestamp 21601
transform 1 0 15548 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_160
timestamp 21601
transform 1 0 15824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_163
timestamp 21601
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_166
timestamp 21601
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_169
timestamp 21601
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_172
timestamp 21601
transform 1 0 16928 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_175
timestamp 21601
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_178
timestamp 21601
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_181
timestamp 21601
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_184
timestamp 21601
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_187
timestamp 21601
transform 1 0 18308 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_190
timestamp 21601
transform 1 0 18584 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_193
timestamp 21601
transform 1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_196
timestamp 21601
transform 1 0 19136 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_199
timestamp 21601
transform 1 0 19412 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_202
timestamp 21601
transform 1 0 19688 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_205
timestamp 21601
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_208
timestamp 21601
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_211
timestamp 21601
transform 1 0 20516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_214
timestamp 21601
transform 1 0 20792 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_217
timestamp 21601
transform 1 0 21068 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_220
timestamp 21601
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 21601
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_225
timestamp 21601
transform 1 0 21804 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_228
timestamp 21601
transform 1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 21601
transform 1 0 22356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 21601
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_90
timestamp 21601
transform 1 0 9384 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_162
timestamp 21601
transform 1 0 16008 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_165
timestamp 21601
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_168
timestamp 21601
transform 1 0 16560 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_171
timestamp 21601
transform 1 0 16836 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_174
timestamp 21601
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_177
timestamp 21601
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_180
timestamp 21601
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_183
timestamp 21601
transform 1 0 17940 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_186
timestamp 21601
transform 1 0 18216 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_189
timestamp 21601
transform 1 0 18492 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_192
timestamp 21601
transform 1 0 18768 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 21601
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_197
timestamp 21601
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_200
timestamp 21601
transform 1 0 19504 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_203
timestamp 21601
transform 1 0 19780 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_206
timestamp 21601
transform 1 0 20056 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_209
timestamp 21601
transform 1 0 20332 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_212
timestamp 21601
transform 1 0 20608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_215
timestamp 21601
transform 1 0 20884 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_218
timestamp 21601
transform 1 0 21160 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp 21601
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_224
timestamp 21601
transform 1 0 21712 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_227
timestamp 21601
transform 1 0 21988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_230
timestamp 21601
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 21601
transform 1 0 1380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_29
timestamp 21601
transform 1 0 3772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_57
timestamp 21601
transform 1 0 6348 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_103
timestamp 21601
transform 1 0 10580 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_106
timestamp 21601
transform 1 0 10856 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_109
timestamp 21601
transform 1 0 11132 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_113
timestamp 21601
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_153
timestamp 21601
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_156
timestamp 21601
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_159
timestamp 21601
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_162
timestamp 21601
transform 1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_165
timestamp 21601
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_169
timestamp 21601
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_172
timestamp 21601
transform 1 0 16928 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_175
timestamp 21601
transform 1 0 17204 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_178
timestamp 21601
transform 1 0 17480 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_181
timestamp 21601
transform 1 0 17756 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_184
timestamp 21601
transform 1 0 18032 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_187
timestamp 21601
transform 1 0 18308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_190
timestamp 21601
transform 1 0 18584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_193
timestamp 21601
transform 1 0 18860 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_196
timestamp 21601
transform 1 0 19136 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_199
timestamp 21601
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_202
timestamp 21601
transform 1 0 19688 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_205
timestamp 21601
transform 1 0 19964 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_208
timestamp 21601
transform 1 0 20240 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_211
timestamp 21601
transform 1 0 20516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_214
timestamp 21601
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_217
timestamp 21601
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_220
timestamp 21601
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 21601
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 21601
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_228
timestamp 21601
transform 1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_231
timestamp 21601
transform 1 0 22356 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_3
timestamp 21601
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_6
timestamp 21601
transform 1 0 1656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_74
timestamp 21601
transform 1 0 7912 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 21601
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_95
timestamp 21601
transform 1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_144
timestamp 21601
transform 1 0 14352 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_147
timestamp 21601
transform 1 0 14628 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 21601
transform 1 0 14904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_153
timestamp 21601
transform 1 0 15180 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_156
timestamp 21601
transform 1 0 15456 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_159
timestamp 21601
transform 1 0 15732 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_162
timestamp 21601
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_165
timestamp 21601
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_168
timestamp 21601
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_171
timestamp 21601
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_174
timestamp 21601
transform 1 0 17112 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_177
timestamp 21601
transform 1 0 17388 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_180
timestamp 21601
transform 1 0 17664 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_183
timestamp 21601
transform 1 0 17940 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_186
timestamp 21601
transform 1 0 18216 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_189
timestamp 21601
transform 1 0 18492 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_192
timestamp 21601
transform 1 0 18768 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 21601
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_197
timestamp 21601
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_200
timestamp 21601
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_203
timestamp 21601
transform 1 0 19780 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_206
timestamp 21601
transform 1 0 20056 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_209
timestamp 21601
transform 1 0 20332 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_212
timestamp 21601
transform 1 0 20608 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_215
timestamp 21601
transform 1 0 20884 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_218
timestamp 21601
transform 1 0 21160 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_221
timestamp 21601
transform 1 0 21436 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_224
timestamp 21601
transform 1 0 21712 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_227
timestamp 21601
transform 1 0 21988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_230
timestamp 21601
transform 1 0 22264 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_64
timestamp 21601
transform 1 0 6992 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_86
timestamp 21601
transform 1 0 9016 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_109
timestamp 21601
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_131
timestamp 21601
transform 1 0 13156 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_154
timestamp 21601
transform 1 0 15272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_157
timestamp 21601
transform 1 0 15548 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_160
timestamp 21601
transform 1 0 15824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_163
timestamp 21601
transform 1 0 16100 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_166
timestamp 21601
transform 1 0 16376 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 21601
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_172
timestamp 21601
transform 1 0 16928 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_175
timestamp 21601
transform 1 0 17204 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_178
timestamp 21601
transform 1 0 17480 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_181
timestamp 21601
transform 1 0 17756 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_184
timestamp 21601
transform 1 0 18032 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_187
timestamp 21601
transform 1 0 18308 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_190
timestamp 21601
transform 1 0 18584 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_193
timestamp 21601
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_196
timestamp 21601
transform 1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_199
timestamp 21601
transform 1 0 19412 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_202
timestamp 21601
transform 1 0 19688 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_205
timestamp 21601
transform 1 0 19964 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_208
timestamp 21601
transform 1 0 20240 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_211
timestamp 21601
transform 1 0 20516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_214
timestamp 21601
transform 1 0 20792 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_217
timestamp 21601
transform 1 0 21068 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_220
timestamp 21601
transform 1 0 21344 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 21601
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 21601
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_228
timestamp 21601
transform 1 0 22080 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_231
timestamp 21601
transform 1 0 22356 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_3
timestamp 21601
transform 1 0 1380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_6
timestamp 21601
transform 1 0 1656 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_29
timestamp 21601
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_52
timestamp 21601
transform 1 0 5888 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_76
timestamp 21601
transform 1 0 8096 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_88
timestamp 21601
transform 1 0 9200 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_98
timestamp 21601
transform 1 0 10120 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_127
timestamp 21601
transform 1 0 12788 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_132
timestamp 21601
transform 1 0 13248 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_135
timestamp 21601
transform 1 0 13524 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_138
timestamp 21601
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_149
timestamp 21601
transform 1 0 14812 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_152
timestamp 21601
transform 1 0 15088 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_155
timestamp 21601
transform 1 0 15364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_158
timestamp 21601
transform 1 0 15640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_161
timestamp 21601
transform 1 0 15916 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_164
timestamp 21601
transform 1 0 16192 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_167
timestamp 21601
transform 1 0 16468 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_170
timestamp 21601
transform 1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_173
timestamp 21601
transform 1 0 17020 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_176
timestamp 21601
transform 1 0 17296 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_179
timestamp 21601
transform 1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_182
timestamp 21601
transform 1 0 17848 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_185
timestamp 21601
transform 1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_188
timestamp 21601
transform 1 0 18400 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_191
timestamp 21601
transform 1 0 18676 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_194
timestamp 21601
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_197
timestamp 21601
transform 1 0 19228 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_200
timestamp 21601
transform 1 0 19504 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_203
timestamp 21601
transform 1 0 19780 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_206
timestamp 21601
transform 1 0 20056 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_209
timestamp 21601
transform 1 0 20332 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_212
timestamp 21601
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_215
timestamp 21601
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_218
timestamp 21601
transform 1 0 21160 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_221
timestamp 21601
transform 1 0 21436 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_224
timestamp 21601
transform 1 0 21712 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_227
timestamp 21601
transform 1 0 21988 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_230
timestamp 21601
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 21601
transform 1 0 3588 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_50
timestamp 21601
transform 1 0 5704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_57
timestamp 21601
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_67
timestamp 21601
transform 1 0 7268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 21601
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_113
timestamp 21601
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_135
timestamp 21601
transform 1 0 13524 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_138
timestamp 21601
transform 1 0 13800 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_141
timestamp 21601
transform 1 0 14076 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_144
timestamp 21601
transform 1 0 14352 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_147
timestamp 21601
transform 1 0 14628 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_150
timestamp 21601
transform 1 0 14904 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_153
timestamp 21601
transform 1 0 15180 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_156
timestamp 21601
transform 1 0 15456 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_159
timestamp 21601
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_162
timestamp 21601
transform 1 0 16008 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_165
timestamp 21601
transform 1 0 16284 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_169
timestamp 21601
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_172
timestamp 21601
transform 1 0 16928 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_175
timestamp 21601
transform 1 0 17204 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_178
timestamp 21601
transform 1 0 17480 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_181
timestamp 21601
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_184
timestamp 21601
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_187
timestamp 21601
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_190
timestamp 21601
transform 1 0 18584 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_193
timestamp 21601
transform 1 0 18860 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_196
timestamp 21601
transform 1 0 19136 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_199
timestamp 21601
transform 1 0 19412 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_202
timestamp 21601
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_205
timestamp 21601
transform 1 0 19964 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_208
timestamp 21601
transform 1 0 20240 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_211
timestamp 21601
transform 1 0 20516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_214
timestamp 21601
transform 1 0 20792 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_217
timestamp 21601
transform 1 0 21068 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_220
timestamp 21601
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 21601
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_9_225
timestamp 21601
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_228
timestamp 21601
transform 1 0 22080 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_231
timestamp 21601
transform 1 0 22356 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 21601
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_6
timestamp 21601
transform 1 0 1656 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 21601
transform 1 0 3772 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_32
timestamp 21601
transform 1 0 4048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_44
timestamp 21601
transform 1 0 5152 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_80
timestamp 21601
transform 1 0 8464 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 21601
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_85
timestamp 21601
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_183
timestamp 21601
transform 1 0 17940 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_186
timestamp 21601
transform 1 0 18216 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_189
timestamp 21601
transform 1 0 18492 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_192
timestamp 21601
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 21601
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 21601
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_200
timestamp 21601
transform 1 0 19504 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_203
timestamp 21601
transform 1 0 19780 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_206
timestamp 21601
transform 1 0 20056 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_209
timestamp 21601
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_212
timestamp 21601
transform 1 0 20608 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_215
timestamp 21601
transform 1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_218
timestamp 21601
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_221
timestamp 21601
transform 1 0 21436 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_224
timestamp 21601
transform 1 0 21712 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_227
timestamp 21601
transform 1 0 21988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_230
timestamp 21601
transform 1 0 22264 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_48
timestamp 21601
transform 1 0 5520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_51
timestamp 21601
transform 1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_54
timestamp 21601
transform 1 0 6072 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 21601
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_66
timestamp 21601
transform 1 0 7176 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_76
timestamp 21601
transform 1 0 8096 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_106
timestamp 21601
transform 1 0 10856 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 21601
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_113
timestamp 21601
transform 1 0 11500 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_116
timestamp 21601
transform 1 0 11776 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_119
timestamp 21601
transform 1 0 12052 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_122
timestamp 21601
transform 1 0 12328 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_125
timestamp 21601
transform 1 0 12604 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 21601
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_169
timestamp 21601
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_172
timestamp 21601
transform 1 0 16928 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_175
timestamp 21601
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_178
timestamp 21601
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_181
timestamp 21601
transform 1 0 17756 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_184
timestamp 21601
transform 1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_187
timestamp 21601
transform 1 0 18308 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_190
timestamp 21601
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_193
timestamp 21601
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_196
timestamp 21601
transform 1 0 19136 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_199
timestamp 21601
transform 1 0 19412 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_202
timestamp 21601
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_205
timestamp 21601
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_208
timestamp 21601
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_211
timestamp 21601
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_214
timestamp 21601
transform 1 0 20792 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_217
timestamp 21601
transform 1 0 21068 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_220
timestamp 21601
transform 1 0 21344 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 21601
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_225
timestamp 21601
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_228
timestamp 21601
transform 1 0 22080 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_231
timestamp 21601
transform 1 0 22356 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 21601
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_57
timestamp 21601
transform 1 0 6348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_79
timestamp 21601
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_82
timestamp 21601
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_85
timestamp 21601
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_88
timestamp 21601
transform 1 0 9200 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_91
timestamp 21601
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 21601
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_144
timestamp 21601
transform 1 0 14352 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_167
timestamp 21601
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_170
timestamp 21601
transform 1 0 16744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_173
timestamp 21601
transform 1 0 17020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_176
timestamp 21601
transform 1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_179
timestamp 21601
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_182
timestamp 21601
transform 1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_185
timestamp 21601
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_188
timestamp 21601
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_191
timestamp 21601
transform 1 0 18676 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 21601
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 21601
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_200
timestamp 21601
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_203
timestamp 21601
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_206
timestamp 21601
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_209
timestamp 21601
transform 1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_212
timestamp 21601
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_215
timestamp 21601
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_218
timestamp 21601
transform 1 0 21160 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_221
timestamp 21601
transform 1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_224
timestamp 21601
transform 1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_227
timestamp 21601
transform 1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_230
timestamp 21601
transform 1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 21601
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_6
timestamp 21601
transform 1 0 1656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_49
timestamp 21601
transform 1 0 5612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_52
timestamp 21601
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 21601
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_88
timestamp 21601
transform 1 0 9200 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_150
timestamp 21601
transform 1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_153
timestamp 21601
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_156
timestamp 21601
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_159
timestamp 21601
transform 1 0 15732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_190
timestamp 21601
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_193
timestamp 21601
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_196
timestamp 21601
transform 1 0 19136 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_199
timestamp 21601
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_202
timestamp 21601
transform 1 0 19688 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_205
timestamp 21601
transform 1 0 19964 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_208
timestamp 21601
transform 1 0 20240 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_211
timestamp 21601
transform 1 0 20516 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_214
timestamp 21601
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_217
timestamp 21601
transform 1 0 21068 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_220
timestamp 21601
transform 1 0 21344 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 21601
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_225
timestamp 21601
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_228
timestamp 21601
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_231
timestamp 21601
transform 1 0 22356 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_3
timestamp 21601
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_6
timestamp 21601
transform 1 0 1656 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_29
timestamp 21601
transform 1 0 3772 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_52
timestamp 21601
transform 1 0 5888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_55
timestamp 21601
transform 1 0 6164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_132
timestamp 21601
transform 1 0 13248 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_135
timestamp 21601
transform 1 0 13524 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 21601
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_157
timestamp 21601
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_182
timestamp 21601
transform 1 0 17848 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_185
timestamp 21601
transform 1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_188
timestamp 21601
transform 1 0 18400 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_191
timestamp 21601
transform 1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 21601
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_197
timestamp 21601
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_200
timestamp 21601
transform 1 0 19504 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_203
timestamp 21601
transform 1 0 19780 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_206
timestamp 21601
transform 1 0 20056 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_209
timestamp 21601
transform 1 0 20332 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_212
timestamp 21601
transform 1 0 20608 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_215
timestamp 21601
transform 1 0 20884 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_218
timestamp 21601
transform 1 0 21160 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_221
timestamp 21601
transform 1 0 21436 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_224
timestamp 21601
transform 1 0 21712 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_227
timestamp 21601
transform 1 0 21988 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_230
timestamp 21601
transform 1 0 22264 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_37
timestamp 21601
transform 1 0 4508 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_40
timestamp 21601
transform 1 0 4784 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_43
timestamp 21601
transform 1 0 5060 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_46
timestamp 21601
transform 1 0 5336 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_78
timestamp 21601
transform 1 0 8280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_128
timestamp 21601
transform 1 0 12880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_158
timestamp 21601
transform 1 0 15640 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_166
timestamp 21601
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_174
timestamp 21601
transform 1 0 17112 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_177
timestamp 21601
transform 1 0 17388 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_200
timestamp 21601
transform 1 0 19504 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_203
timestamp 21601
transform 1 0 19780 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_206
timestamp 21601
transform 1 0 20056 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_209
timestamp 21601
transform 1 0 20332 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_212
timestamp 21601
transform 1 0 20608 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_215
timestamp 21601
transform 1 0 20884 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_218
timestamp 21601
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_221
timestamp 21601
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_225
timestamp 21601
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_228
timestamp 21601
transform 1 0 22080 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp 21601
transform 1 0 22356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 21601
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_6
timestamp 21601
transform 1 0 1656 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_23
timestamp 21601
transform 1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 21601
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_37
timestamp 21601
transform 1 0 4508 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 21601
transform 1 0 7728 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_81
timestamp 21601
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_98
timestamp 21601
transform 1 0 10120 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_101
timestamp 21601
transform 1 0 10396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_110
timestamp 21601
transform 1 0 11224 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_134
timestamp 21601
transform 1 0 13432 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_141
timestamp 21601
transform 1 0 14076 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_185
timestamp 21601
transform 1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_188
timestamp 21601
transform 1 0 18400 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_191
timestamp 21601
transform 1 0 18676 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_194
timestamp 21601
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 21601
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_200
timestamp 21601
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_203
timestamp 21601
transform 1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_206
timestamp 21601
transform 1 0 20056 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_209
timestamp 21601
transform 1 0 20332 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_212
timestamp 21601
transform 1 0 20608 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_215
timestamp 21601
transform 1 0 20884 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_218
timestamp 21601
transform 1 0 21160 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_221
timestamp 21601
transform 1 0 21436 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_224
timestamp 21601
transform 1 0 21712 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_227
timestamp 21601
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_230
timestamp 21601
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 21601
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_30
timestamp 21601
transform 1 0 3864 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 21601
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 21601
transform 1 0 7544 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_93
timestamp 21601
transform 1 0 9660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_110
timestamp 21601
transform 1 0 11224 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_121
timestamp 21601
transform 1 0 12236 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_124
timestamp 21601
transform 1 0 12512 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_127
timestamp 21601
transform 1 0 12788 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 21601
transform 1 0 16376 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_193
timestamp 21601
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_196
timestamp 21601
transform 1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_199
timestamp 21601
transform 1 0 19412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_202
timestamp 21601
transform 1 0 19688 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_205
timestamp 21601
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_208
timestamp 21601
transform 1 0 20240 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_211
timestamp 21601
transform 1 0 20516 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_214
timestamp 21601
transform 1 0 20792 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_217
timestamp 21601
transform 1 0 21068 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_220
timestamp 21601
transform 1 0 21344 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 21601
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_225
timestamp 21601
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_228
timestamp 21601
transform 1 0 22080 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_231
timestamp 21601
transform 1 0 22356 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 21601
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_6
timestamp 21601
transform 1 0 1656 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_29
timestamp 21601
transform 1 0 3772 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_88
timestamp 21601
transform 1 0 9200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 21601
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_141
timestamp 21601
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_171
timestamp 21601
transform 1 0 16836 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_174
timestamp 21601
transform 1 0 17112 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_177
timestamp 21601
transform 1 0 17388 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_180
timestamp 21601
transform 1 0 17664 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_183
timestamp 21601
transform 1 0 17940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_186
timestamp 21601
transform 1 0 18216 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_189
timestamp 21601
transform 1 0 18492 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_192
timestamp 21601
transform 1 0 18768 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 21601
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 21601
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_200
timestamp 21601
transform 1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_203
timestamp 21601
transform 1 0 19780 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_206
timestamp 21601
transform 1 0 20056 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_209
timestamp 21601
transform 1 0 20332 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_212
timestamp 21601
transform 1 0 20608 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_215
timestamp 21601
transform 1 0 20884 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_218
timestamp 21601
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_221
timestamp 21601
transform 1 0 21436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_224
timestamp 21601
transform 1 0 21712 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_227
timestamp 21601
transform 1 0 21988 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_230
timestamp 21601
transform 1 0 22264 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_3
timestamp 21601
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_23
timestamp 21601
transform 1 0 3220 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_62
timestamp 21601
transform 1 0 6808 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_92
timestamp 21601
transform 1 0 9568 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_118
timestamp 21601
transform 1 0 11960 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_121
timestamp 21601
transform 1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_124
timestamp 21601
transform 1 0 12512 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_133
timestamp 21601
transform 1 0 13340 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_136
timestamp 21601
transform 1 0 13616 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_160
timestamp 21601
transform 1 0 15824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_163
timestamp 21601
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 21601
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_201
timestamp 21601
transform 1 0 19596 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_204
timestamp 21601
transform 1 0 19872 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_207
timestamp 21601
transform 1 0 20148 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_210
timestamp 21601
transform 1 0 20424 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_213
timestamp 21601
transform 1 0 20700 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_217
timestamp 21601
transform 1 0 21068 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_220
timestamp 21601
transform 1 0 21344 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 21601
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_225
timestamp 21601
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_228
timestamp 21601
transform 1 0 22080 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_231
timestamp 21601
transform 1 0 22356 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 21601
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_127
timestamp 21601
transform 1 0 12788 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 21601
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_178
timestamp 21601
transform 1 0 17480 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_231
timestamp 21601
transform 1 0 22356 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_3
timestamp 21601
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_33
timestamp 21601
transform 1 0 4140 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_57
timestamp 21601
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 21601
transform 1 0 16376 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_202
timestamp 21601
transform 1 0 19688 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 21601
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_37
timestamp 21601
transform 1 0 4508 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_40
timestamp 21601
transform 1 0 4784 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_57
timestamp 21601
transform 1 0 6348 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_60
timestamp 21601
transform 1 0 6624 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 21601
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_85
timestamp 21601
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_88
timestamp 21601
transform 1 0 9200 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_91
timestamp 21601
transform 1 0 9476 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_94
timestamp 21601
transform 1 0 9752 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_113
timestamp 21601
transform 1 0 11500 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_124
timestamp 21601
transform 1 0 12512 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_127
timestamp 21601
transform 1 0 12788 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_130
timestamp 21601
transform 1 0 13064 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_133
timestamp 21601
transform 1 0 13340 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_136
timestamp 21601
transform 1 0 13616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 21601
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_165
timestamp 21601
transform 1 0 16284 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 21601
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_205
timestamp 21601
transform 1 0 19964 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_208
timestamp 21601
transform 1 0 20240 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_225
timestamp 21601
transform 1 0 21804 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_228
timestamp 21601
transform 1 0 22080 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_231
timestamp 21601
transform 1 0 22356 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 21601
transform -1 0 14812 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 21601
transform -1 0 14720 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 21601
transform -1 0 22540 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 21601
transform -1 0 14812 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 21601
transform -1 0 14536 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  pclk_div_skewed_delay.dly_clkbuf
timestamp 21601
transform -1 0 18676 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  pclk_div_skewed_delay.gen_dlygen\[1\].dlygen
timestamp 21601
transform 1 0 16008 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  pclk_div_skewed_delay.gen_dlygen\[2\].dlygen
timestamp 21601
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  pclk_div_skewed_delay.gen_dlygen\[3\].dlygen
timestamp 21601
transform 1 0 16744 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  pclk_div_skewed_delay.gen_dlygen\[4\].dlygen
timestamp 21601
transform 1 0 17388 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  pclk_div_skewed_delay.gen_dlygen\[5\].dlygen
timestamp 21601
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_23
timestamp 21601
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 21601
transform -1 0 22816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_24
timestamp 21601
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 21601
transform -1 0 22816 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_25
timestamp 21601
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 21601
transform -1 0 22816 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_26
timestamp 21601
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 21601
transform -1 0 22816 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_27
timestamp 21601
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 21601
transform -1 0 22816 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_28
timestamp 21601
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 21601
transform -1 0 22816 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_29
timestamp 21601
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 21601
transform -1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_30
timestamp 21601
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 21601
transform -1 0 22816 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_31
timestamp 21601
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 21601
transform -1 0 22816 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_32
timestamp 21601
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 21601
transform -1 0 22816 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_33
timestamp 21601
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 21601
transform -1 0 22816 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_34
timestamp 21601
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 21601
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_35
timestamp 21601
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 21601
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_36
timestamp 21601
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 21601
transform -1 0 22816 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_37
timestamp 21601
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 21601
transform -1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_38
timestamp 21601
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 21601
transform -1 0 22816 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_39
timestamp 21601
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 21601
transform -1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_40
timestamp 21601
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 21601
transform -1 0 22816 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_41
timestamp 21601
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 21601
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_42
timestamp 21601
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 21601
transform -1 0 22816 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_43
timestamp 21601
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 21601
transform -1 0 22816 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_44
timestamp 21601
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 21601
transform -1 0 22816 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_45
timestamp 21601
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 21601
transform -1 0 22816 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_46
timestamp 21601
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_47
timestamp 21601
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_48
timestamp 21601
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_49
timestamp 21601
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_50
timestamp 21601
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_51
timestamp 21601
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_52
timestamp 21601
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_53
timestamp 21601
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_54
timestamp 21601
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_55
timestamp 21601
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_56
timestamp 21601
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_57
timestamp 21601
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_58
timestamp 21601
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_59
timestamp 21601
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_60
timestamp 21601
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_61
timestamp 21601
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_62
timestamp 21601
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_63
timestamp 21601
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_64
timestamp 21601
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_65
timestamp 21601
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_66
timestamp 21601
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_67
timestamp 21601
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_68
timestamp 21601
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_69
timestamp 21601
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_70
timestamp 21601
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_71
timestamp 21601
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_72
timestamp 21601
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_73
timestamp 21601
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_74
timestamp 21601
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_75
timestamp 21601
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_76
timestamp 21601
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_77
timestamp 21601
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_78
timestamp 21601
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_79
timestamp 21601
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_80
timestamp 21601
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_81
timestamp 21601
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_82
timestamp 21601
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_83
timestamp 21601
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_84
timestamp 21601
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_85
timestamp 21601
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_86
timestamp 21601
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_87
timestamp 21601
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_88
timestamp 21601
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_89
timestamp 21601
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_90
timestamp 21601
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_91
timestamp 21601
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_92
timestamp 21601
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_93
timestamp 21601
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_94
timestamp 21601
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_95
timestamp 21601
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_96
timestamp 21601
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_97
timestamp 21601
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_98
timestamp 21601
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_99
timestamp 21601
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_100
timestamp 21601
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 21601
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_102
timestamp 21601
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_103
timestamp 21601
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 21601
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_105
timestamp 21601
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_106
timestamp 21601
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 21601
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_108
timestamp 21601
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp 21601
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 21601
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_111
timestamp 21601
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp 21601
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_113
timestamp 21601
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_114
timestamp 21601
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp 21601
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_116
timestamp 21601
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_117
timestamp 21601
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp 21601
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_119
timestamp 21601
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_120
timestamp 21601
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_121
timestamp 21601
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_122
timestamp 21601
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_123
timestamp 21601
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_124
timestamp 21601
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_125
timestamp 21601
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_126
timestamp 21601
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_127
timestamp 21601
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_128
timestamp 21601
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_129
timestamp 21601
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_130
timestamp 21601
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_131
timestamp 21601
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_132
timestamp 21601
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_133
timestamp 21601
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_134
timestamp 21601
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_135
timestamp 21601
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_136
timestamp 21601
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_137
timestamp 21601
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_138
timestamp 21601
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_139
timestamp 21601
transform 1 0 6256 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_140
timestamp 21601
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_141
timestamp 21601
transform 1 0 11408 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_142
timestamp 21601
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_143
timestamp 21601
transform 1 0 16560 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_144
timestamp 21601
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_145
timestamp 21601
transform 1 0 21712 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  usb_clk_delayed.dly_clkbuf
timestamp 21601
transform -1 0 19688 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[1\].dlygen
timestamp 21601
transform 1 0 13800 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[2\].dlygen
timestamp 21601
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[3\].dlygen
timestamp 21601
transform 1 0 16100 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[4\].dlygen
timestamp 21601
transform 1 0 16652 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[5\].dlygen
timestamp 21601
transform 1 0 17388 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[6\].dlygen
timestamp 21601
transform 1 0 18124 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[7\].dlygen
timestamp 21601
transform -1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[8\].dlygen
timestamp 21601
transform 1 0 18400 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  usb_clk_delayed.gen_dlygen\[9\].dlygen
timestamp 21601
transform 1 0 18860 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_8  user_clk_delay.dly_clkbuf
timestamp 21601
transform 1 0 19228 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkdlybuf4s18_2  user_clk_delay.gen_dlygen\[1\].dlygen
timestamp 21601
transform 1 0 19228 0 1 13056
box -38 -48 774 592
<< labels >>
flabel metal4 s 8208 1040 8528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16208 1040 16528 13648 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 1040 4528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 12208 1040 12528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 20208 1040 20528 13648 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 16486 14200 16542 15000 0 FreeSans 224 90 0 0 clk
port 2 nsew signal output
flabel metal2 s 21638 14200 21694 15000 0 FreeSans 224 90 0 0 clk_mon
port 3 nsew signal output
flabel metal2 s 10046 14200 10102 15000 0 FreeSans 224 90 0 0 clk_mon_sel[0]
port 4 nsew signal input
flabel metal2 s 11334 14200 11390 15000 0 FreeSans 224 90 0 0 clk_mon_sel[1]
port 5 nsew signal input
flabel metal2 s 12622 14200 12678 15000 0 FreeSans 224 90 0 0 clk_mon_sel[2]
port 6 nsew signal input
flabel metal2 s 1030 14200 1086 15000 0 FreeSans 224 90 0 0 clk_mux1_out
port 7 nsew signal output
flabel metal3 s 23200 7352 24000 7472 0 FreeSans 480 0 0 0 dll_clk
port 8 nsew signal input
flabel metal3 s 23200 12248 24000 12368 0 FreeSans 480 0 0 0 dll_clk90
port 9 nsew signal input
flabel metal3 s 23200 2456 24000 2576 0 FreeSans 480 0 0 0 hkrst_n
port 10 nsew signal input
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 hsxo
port 11 nsew signal input
flabel metal2 s 4894 14200 4950 15000 0 FreeSans 224 90 0 0 hsxo_en
port 12 nsew signal input
flabel metal2 s 17498 0 17554 800 0 FreeSans 224 90 0 0 hsxo_en_tf
port 13 nsew signal output
flabel metal2 s 8758 14200 8814 15000 0 FreeSans 224 90 0 0 hsxo_standby
port 14 nsew signal input
flabel metal2 s 23018 0 23074 800 0 FreeSans 224 90 0 0 hsxo_standby_tf
port 15 nsew signal output
flabel metal2 s 8298 0 8354 800 0 FreeSans 224 90 0 0 lsxo
port 16 nsew signal input
flabel metal2 s 6182 14200 6238 15000 0 FreeSans 224 90 0 0 lsxo_en
port 17 nsew signal input
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 lsxo_en_tf
port 18 nsew signal output
flabel metal2 s 7470 14200 7526 15000 0 FreeSans 224 90 0 0 lsxo_standby
port 19 nsew signal input
flabel metal2 s 21178 0 21234 800 0 FreeSans 224 90 0 0 lsxo_standby_tf
port 20 nsew signal output
flabel metal2 s 17774 14200 17830 15000 0 FreeSans 224 90 0 0 pclk
port 21 nsew signal output
flabel metal2 s 11978 0 12034 800 0 FreeSans 224 90 0 0 por_n
port 22 nsew signal input
flabel metal2 s 4618 0 4674 800 0 FreeSans 224 90 0 0 rcosc_16m
port 23 nsew signal input
flabel metal2 s 3606 14200 3662 15000 0 FreeSans 224 90 0 0 rcosc_16m_en
port 24 nsew signal input
flabel metal2 s 15658 0 15714 800 0 FreeSans 224 90 0 0 rcosc_16m_en_tf
port 25 nsew signal output
flabel metal2 s 2778 0 2834 800 0 FreeSans 224 90 0 0 rcosc_500k
port 26 nsew signal input
flabel metal2 s 2318 14200 2374 15000 0 FreeSans 224 90 0 0 rcosc_500k_en
port 27 nsew signal input
flabel metal2 s 13818 0 13874 800 0 FreeSans 224 90 0 0 rcosc_500k_en_tf
port 28 nsew signal output
flabel metal2 s 22926 14200 22982 15000 0 FreeSans 224 90 0 0 rst_n
port 29 nsew signal output
flabel metal3 s 0 6536 800 6656 0 FreeSans 480 0 0 0 sel_clkdiv0[0]
port 30 nsew signal input
flabel metal3 s 0 7352 800 7472 0 FreeSans 480 0 0 0 sel_clkdiv0[1]
port 31 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 sel_clkdiv0[2]
port 32 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 sel_clkdiv1[0]
port 33 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 sel_clkdiv1[1]
port 34 nsew signal input
flabel metal3 s 0 10616 800 10736 0 FreeSans 480 0 0 0 sel_clkdiv1[2]
port 35 nsew signal input
flabel metal3 s 0 11432 800 11552 0 FreeSans 480 0 0 0 sel_clkdiv2[0]
port 36 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 sel_clkdiv2[1]
port 37 nsew signal input
flabel metal3 s 0 13064 800 13184 0 FreeSans 480 0 0 0 sel_clkdiv2[2]
port 38 nsew signal input
flabel metal3 s 0 1640 800 1760 0 FreeSans 480 0 0 0 sel_mux0
port 39 nsew signal input
flabel metal3 s 0 2456 800 2576 0 FreeSans 480 0 0 0 sel_mux1
port 40 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 sel_mux2
port 41 nsew signal input
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 sel_mux3
port 42 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 sel_mux4
port 43 nsew signal input
flabel metal3 s 0 5720 800 5840 0 FreeSans 480 0 0 0 sel_mux5
port 44 nsew signal input
flabel metal2 s 19062 14200 19118 15000 0 FreeSans 224 90 0 0 usb_clk
port 45 nsew signal output
flabel metal2 s 20350 14200 20406 15000 0 FreeSans 224 90 0 0 user_clk
port 46 nsew signal output
flabel metal2 s 13910 14200 13966 15000 0 FreeSans 224 90 0 0 user_dly_sel[0]
port 47 nsew signal input
flabel metal2 s 15198 14200 15254 15000 0 FreeSans 224 90 0 0 user_dly_sel[1]
port 48 nsew signal input
flabel metal2 s 938 0 994 800 0 FreeSans 224 90 0 0 xclk
port 49 nsew signal input
flabel metal2 s 10138 0 10194 800 0 FreeSans 224 90 0 0 xrst_n
port 50 nsew signal input
rlabel metal1 11960 13056 11960 13056 0 VGND
rlabel metal1 11960 13600 11960 13600 0 VPWR
rlabel metal2 5566 6562 5566 6562 0 CLKDIV_0.CLK_DIV_MUX.clk0
rlabel metal1 8786 5678 8786 5678 0 CLKDIV_0.CLK_DIV_MUX.clk1
rlabel metal1 9841 6766 9841 6766 0 CLKDIV_0.CLK_DIV_MUX.clk2
rlabel metal1 9890 6664 9890 6664 0 CLKDIV_0.CLK_DIV_MUX.clk3
rlabel metal2 7498 7072 7498 7072 0 CLKDIV_0.CLK_DIV_MUX.clko
rlabel metal2 7774 4930 7774 4930 0 CLKDIV_0.CLK_DIV_MUX.m1.Q1a
rlabel metal1 8556 5610 8556 5610 0 CLKDIV_0.CLK_DIV_MUX.m1.Q1b
rlabel metal1 10120 4250 10120 4250 0 CLKDIV_0.CLK_DIV_MUX.m1.Q2a
rlabel metal2 7130 5882 7130 5882 0 CLKDIV_0.CLK_DIV_MUX.m1.Q2b
rlabel metal2 6302 5100 6302 5100 0 CLKDIV_0.CLK_DIV_MUX.m1.q1a_in
rlabel metal2 8694 4794 8694 4794 0 CLKDIV_0.CLK_DIV_MUX.m1.q2a_in
rlabel metal1 12098 5882 12098 5882 0 CLKDIV_0.CLK_DIV_MUX.m2.Q1a
rlabel metal2 10074 5916 10074 5916 0 CLKDIV_0.CLK_DIV_MUX.m2.Q1b
rlabel metal1 11316 6426 11316 6426 0 CLKDIV_0.CLK_DIV_MUX.m2.Q2a
rlabel metal2 10074 6596 10074 6596 0 CLKDIV_0.CLK_DIV_MUX.m2.Q2b
rlabel metal2 10718 6426 10718 6426 0 CLKDIV_0.CLK_DIV_MUX.m2.q1a_in
rlabel metal1 9706 5882 9706 5882 0 CLKDIV_0.CLK_DIV_MUX.m2.q2a_in
rlabel metal1 7452 7922 7452 7922 0 CLKDIV_0.CLK_DIV_MUX.m3.Q1a
rlabel metal1 8280 8058 8280 8058 0 CLKDIV_0.CLK_DIV_MUX.m3.Q1b
rlabel metal1 10074 7514 10074 7514 0 CLKDIV_0.CLK_DIV_MUX.m3.Q2a
rlabel metal2 8050 7548 8050 7548 0 CLKDIV_0.CLK_DIV_MUX.m3.Q2b
rlabel metal1 6808 7514 6808 7514 0 CLKDIV_0.CLK_DIV_MUX.m3.q1a_in
rlabel metal1 8648 7446 8648 7446 0 CLKDIV_0.CLK_DIV_MUX.m3.q2a_in
rlabel metal2 2070 7650 2070 7650 0 CLKDIV_0.DIV_BYPASS_MUX.Q1a
rlabel metal1 3312 8058 3312 8058 0 CLKDIV_0.DIV_BYPASS_MUX.Q1b
rlabel metal1 5060 7514 5060 7514 0 CLKDIV_0.DIV_BYPASS_MUX.Q2a
rlabel metal1 1794 6324 1794 6324 0 CLKDIV_0.DIV_BYPASS_MUX.Q2b
rlabel metal1 3312 7378 3312 7378 0 CLKDIV_0.DIV_BYPASS_MUX.clk1
rlabel metal2 1702 6868 1702 6868 0 CLKDIV_0.DIV_BYPASS_MUX.q1a_in
rlabel metal2 3910 7582 3910 7582 0 CLKDIV_0.DIV_BYPASS_MUX.q2a_in
rlabel metal2 12650 9044 12650 9044 0 CLKDIV_1.CLK_DIV_MUX.clk0
rlabel metal1 10304 9962 10304 9962 0 CLKDIV_1.CLK_DIV_MUX.clk1
rlabel metal1 16698 8500 16698 8500 0 CLKDIV_1.CLK_DIV_MUX.clk2
rlabel metal2 15502 8772 15502 8772 0 CLKDIV_1.CLK_DIV_MUX.clk3
rlabel metal1 13662 10030 13662 10030 0 CLKDIV_1.CLK_DIV_MUX.clko
rlabel metal1 8970 9010 8970 9010 0 CLKDIV_1.CLK_DIV_MUX.m1.Q1a
rlabel metal2 10718 8704 10718 8704 0 CLKDIV_1.CLK_DIV_MUX.m1.Q1b
rlabel metal2 11730 8126 11730 8126 0 CLKDIV_1.CLK_DIV_MUX.m1.Q2a
rlabel metal2 10534 9690 10534 9690 0 CLKDIV_1.CLK_DIV_MUX.m1.Q2b
rlabel metal1 6624 9078 6624 9078 0 CLKDIV_1.CLK_DIV_MUX.m1.q1a_in
rlabel metal1 10396 8398 10396 8398 0 CLKDIV_1.CLK_DIV_MUX.m1.q2a_in
rlabel metal2 18446 9044 18446 9044 0 CLKDIV_1.CLK_DIV_MUX.m2.Q1a
rlabel metal1 16330 9418 16330 9418 0 CLKDIV_1.CLK_DIV_MUX.m2.Q1b
rlabel metal1 14996 7786 14996 7786 0 CLKDIV_1.CLK_DIV_MUX.m2.Q2a
rlabel metal1 16560 8466 16560 8466 0 CLKDIV_1.CLK_DIV_MUX.m2.Q2b
rlabel metal2 16974 8908 16974 8908 0 CLKDIV_1.CLK_DIV_MUX.m2.q1a_in
rlabel metal1 15916 8874 15916 8874 0 CLKDIV_1.CLK_DIV_MUX.m2.q2a_in
rlabel metal1 14904 9486 14904 9486 0 CLKDIV_1.CLK_DIV_MUX.m3.Q1a
rlabel metal2 15778 10404 15778 10404 0 CLKDIV_1.CLK_DIV_MUX.m3.Q1b
rlabel metal2 17986 10404 17986 10404 0 CLKDIV_1.CLK_DIV_MUX.m3.Q2a
rlabel metal2 15686 10438 15686 10438 0 CLKDIV_1.CLK_DIV_MUX.m3.Q2b
rlabel metal1 13524 9622 13524 9622 0 CLKDIV_1.CLK_DIV_MUX.m3.q1a_in
rlabel metal2 16514 10268 16514 10268 0 CLKDIV_1.CLK_DIV_MUX.m3.q2a_in
rlabel metal1 11454 11186 11454 11186 0 CLKDIV_1.DIV_BYPASS_MUX.Q1a
rlabel metal1 12880 11322 12880 11322 0 CLKDIV_1.DIV_BYPASS_MUX.Q1b
rlabel metal1 15318 10778 15318 10778 0 CLKDIV_1.DIV_BYPASS_MUX.Q2a
rlabel via1 13572 11118 13572 11118 0 CLKDIV_1.DIV_BYPASS_MUX.Q2b
rlabel metal1 13156 11050 13156 11050 0 CLKDIV_1.DIV_BYPASS_MUX.clk0
rlabel metal2 13478 11390 13478 11390 0 CLKDIV_1.DIV_BYPASS_MUX.clk1
rlabel metal2 13754 11764 13754 11764 0 CLKDIV_1.DIV_BYPASS_MUX.clko
rlabel metal2 10902 11390 10902 11390 0 CLKDIV_1.DIV_BYPASS_MUX.q1a_in
rlabel metal2 13386 11118 13386 11118 0 CLKDIV_1.DIV_BYPASS_MUX.q2a_in
rlabel metal2 1702 11186 1702 11186 0 CLKDIV_2.CLK_DIV_MUX.clk0
rlabel metal1 2346 11771 2346 11771 0 CLKDIV_2.CLK_DIV_MUX.clk1
rlabel metal1 4370 11118 4370 11118 0 CLKDIV_2.CLK_DIV_MUX.clk2
rlabel metal2 6946 11390 6946 11390 0 CLKDIV_2.CLK_DIV_MUX.clk3
rlabel metal1 7774 12750 7774 12750 0 CLKDIV_2.CLK_DIV_MUX.clko
rlabel metal1 2024 12886 2024 12886 0 CLKDIV_2.CLK_DIV_MUX.m1.Q1a
rlabel metal1 2162 12682 2162 12682 0 CLKDIV_2.CLK_DIV_MUX.m1.Q1b
rlabel metal2 3634 11934 3634 11934 0 CLKDIV_2.CLK_DIV_MUX.m1.Q2a
rlabel metal1 3772 13294 3772 13294 0 CLKDIV_2.CLK_DIV_MUX.m1.Q2b
rlabel metal1 2944 11866 2944 11866 0 CLKDIV_2.CLK_DIV_MUX.m1.q1a_in
rlabel metal2 2070 12376 2070 12376 0 CLKDIV_2.CLK_DIV_MUX.m1.q2a_in
rlabel metal1 6670 11322 6670 11322 0 CLKDIV_2.CLK_DIV_MUX.m2.Q1a
rlabel metal1 7452 12070 7452 12070 0 CLKDIV_2.CLK_DIV_MUX.m2.Q1b
rlabel metal1 9016 10574 9016 10574 0 CLKDIV_2.CLK_DIV_MUX.m2.Q2a
rlabel metal1 6394 11730 6394 11730 0 CLKDIV_2.CLK_DIV_MUX.m2.Q2b
rlabel metal1 5888 11186 5888 11186 0 CLKDIV_2.CLK_DIV_MUX.m2.q1a_in
rlabel metal1 7951 11322 7951 11322 0 CLKDIV_2.CLK_DIV_MUX.m2.q2a_in
rlabel metal1 4554 12410 4554 12410 0 CLKDIV_2.CLK_DIV_MUX.m3.Q1a
rlabel metal2 6118 13090 6118 13090 0 CLKDIV_2.CLK_DIV_MUX.m3.Q1b
rlabel metal1 8280 11662 8280 11662 0 CLKDIV_2.CLK_DIV_MUX.m3.Q2a
rlabel metal1 6900 12818 6900 12818 0 CLKDIV_2.CLK_DIV_MUX.m3.Q2b
rlabel metal1 5566 13158 5566 13158 0 CLKDIV_2.CLK_DIV_MUX.m3.q1a_in
rlabel metal1 7130 13192 7130 13192 0 CLKDIV_2.CLK_DIV_MUX.m3.q2a_in
rlabel metal1 11178 12104 11178 12104 0 CLKDIV_2.DIV_BYPASS_MUX.Q1a
rlabel metal1 10672 13226 10672 13226 0 CLKDIV_2.DIV_BYPASS_MUX.Q1b
rlabel metal1 11546 12750 11546 12750 0 CLKDIV_2.DIV_BYPASS_MUX.Q2a
rlabel metal2 13294 13124 13294 13124 0 CLKDIV_2.DIV_BYPASS_MUX.Q2b
rlabel metal1 9430 12750 9430 12750 0 CLKDIV_2.DIV_BYPASS_MUX.clk1
rlabel metal1 19274 13362 19274 13362 0 CLKDIV_2.DIV_BYPASS_MUX.clko
rlabel metal1 10672 13158 10672 13158 0 CLKDIV_2.DIV_BYPASS_MUX.q1a_in
rlabel metal2 9798 13022 9798 13022 0 CLKDIV_2.DIV_BYPASS_MUX.q2a_in
rlabel metal1 1978 1530 1978 1530 0 CLKMUX_0.Q1a
rlabel metal1 3956 2074 3956 2074 0 CLKMUX_0.Q1b
rlabel metal1 4278 1530 4278 1530 0 CLKMUX_0.Q2a
rlabel metal1 6072 1870 6072 1870 0 CLKMUX_0.Q2b
rlabel metal1 5980 1258 5980 1258 0 CLKMUX_0.q1a_in
rlabel metal1 5529 1530 5529 1530 0 CLKMUX_0.q2a_in
rlabel metal1 1840 2958 1840 2958 0 CLKMUX_1.Q1a
rlabel metal1 2070 1972 2070 1972 0 CLKMUX_1.Q1b
rlabel metal1 4186 2312 4186 2312 0 CLKMUX_1.Q2a
rlabel metal1 5888 2278 5888 2278 0 CLKMUX_1.Q2b
rlabel metal3 4462 2924 4462 2924 0 CLKMUX_1.q1a_in
rlabel metal1 1840 2074 1840 2074 0 CLKMUX_1.q2a_in
rlabel metal1 1794 5338 1794 5338 0 CLKMUX_2.Q1a
rlabel via1 2159 6290 2159 6290 0 CLKMUX_2.Q1b
rlabel metal1 4002 4658 4002 4658 0 CLKMUX_2.Q2a
rlabel metal2 2346 5916 2346 5916 0 CLKMUX_2.Q2b
rlabel metal1 4462 4250 4462 4250 0 CLKMUX_2.q1a_in
rlabel metal1 1840 4250 1840 4250 0 CLKMUX_2.q2a_in
rlabel metal1 6762 3128 6762 3128 0 CLKMUX_3.Q1a
rlabel via1 6764 1938 6764 1938 0 CLKMUX_3.Q1b
rlabel metal2 5290 3672 5290 3672 0 CLKMUX_3.Q2a
rlabel metal1 6762 3604 6762 3604 0 CLKMUX_3.Q2b
rlabel metal1 5520 2958 5520 2958 0 CLKMUX_3.q1a_in
rlabel metal1 2254 4046 2254 4046 0 CLKMUX_3.q2a_in
rlabel metal1 9062 2958 9062 2958 0 CLKMUX_4.Q1a
rlabel metal1 8970 4590 8970 4590 0 CLKMUX_4.Q1b
rlabel metal1 9246 3570 9246 3570 0 CLKMUX_4.Q2a
rlabel metal1 8211 4590 8211 4590 0 CLKMUX_4.Q2b
rlabel metal1 2714 9928 2714 9928 0 CLKMUX_4.clko
rlabel metal1 4830 3672 4830 3672 0 CLKMUX_4.q1a_in
rlabel metal1 7222 3400 7222 3400 0 CLKMUX_4.q2a_in
rlabel metal1 3956 8534 3956 8534 0 CLKMUX_5.Q1a
rlabel metal1 5198 9554 5198 9554 0 CLKMUX_5.Q1b
rlabel metal1 3910 8874 3910 8874 0 CLKMUX_5.Q2a
rlabel via1 6006 9554 6006 9554 0 CLKMUX_5.Q2b
rlabel metal1 2484 8602 2484 8602 0 CLKMUX_5.q1a_in
rlabel metal1 1784 9146 1784 9146 0 CLKMUX_5.q2a_in
rlabel metal1 12558 2618 12558 2618 0 CLK_MON_MUX_0.m1.Q1a
rlabel metal1 14142 3026 14142 3026 0 CLK_MON_MUX_0.m1.Q1b
rlabel metal1 14398 3400 14398 3400 0 CLK_MON_MUX_0.m1.Q2a
rlabel metal1 15226 3094 15226 3094 0 CLK_MON_MUX_0.m1.Q2b
rlabel metal1 11040 2482 11040 2482 0 CLK_MON_MUX_0.m1.q1a_in
rlabel metal1 12374 3400 12374 3400 0 CLK_MON_MUX_0.m1.q2a_in
rlabel metal1 7406 1530 7406 1530 0 CLK_MON_MUX_0.m2.Q1a
rlabel via1 9432 2414 9432 2414 0 CLK_MON_MUX_0.m2.Q1b
rlabel metal1 9896 1530 9896 1530 0 CLK_MON_MUX_0.m2.Q2a
rlabel metal1 9338 1360 9338 1360 0 CLK_MON_MUX_0.m2.Q2b
rlabel metal1 8740 1258 8740 1258 0 CLK_MON_MUX_0.m2.q1a_in
rlabel metal1 10258 2516 10258 2516 0 CLK_MON_MUX_0.m2.q2a_in
rlabel metal1 13754 4794 13754 4794 0 CLK_MON_MUX_0.m3.Q1a
rlabel metal1 12466 5270 12466 5270 0 CLK_MON_MUX_0.m3.Q1b
rlabel metal2 12098 4318 12098 4318 0 CLK_MON_MUX_0.m3.Q2a
rlabel metal1 13156 5270 13156 5270 0 CLK_MON_MUX_0.m3.Q2b
rlabel metal2 12742 5168 12742 5168 0 CLK_MON_MUX_0.m3.q1a_in
rlabel metal1 11040 4658 11040 4658 0 CLK_MON_MUX_0.m3.q2a_in
rlabel metal1 16090 6970 16090 6970 0 CLK_MON_MUX_1.Q1a
rlabel metal2 15410 7140 15410 7140 0 CLK_MON_MUX_1.Q1b
rlabel metal1 14398 6664 14398 6664 0 CLK_MON_MUX_1.Q2a
rlabel metal2 15686 7548 15686 7548 0 CLK_MON_MUX_1.Q2b
rlabel metal1 19826 12852 19826 12852 0 CLK_MON_MUX_1.clko
rlabel metal2 13754 7582 13754 7582 0 CLK_MON_MUX_1.q1a_in
rlabel metal2 12926 7072 12926 7072 0 CLK_MON_MUX_1.q2a_in
rlabel metal2 14674 1530 14674 1530 0 RST_SYNC.delay\[0\]
rlabel metal1 13938 1190 13938 1190 0 RST_SYNC.delay\[1\]
rlabel via1 12558 1275 12558 1275 0 RST_SYNC.rst_n_in
rlabel metal1 15042 11866 15042 11866 0 _000_
rlabel metal2 11822 4556 11822 4556 0 _001_
rlabel metal1 13248 5202 13248 5202 0 _002_
rlabel metal2 16054 7004 16054 7004 0 _003_
rlabel metal1 3772 2482 3772 2482 0 _004_
rlabel metal2 3818 4828 3818 4828 0 _005_
rlabel metal1 1702 7854 1702 7854 0 _006_
rlabel metal1 5428 3570 5428 3570 0 _007_
rlabel metal1 6532 7514 6532 7514 0 _008_
rlabel metal1 11086 7514 11086 7514 0 _009_
rlabel metal1 10258 3060 10258 3060 0 _010_
rlabel metal1 11086 11866 11086 11866 0 _011_
rlabel metal2 15502 9758 15502 9758 0 _012_
rlabel metal1 18814 10710 18814 10710 0 _013_
rlabel metal2 4370 12988 4370 12988 0 _014_
rlabel metal1 7176 12614 7176 12614 0 _015_
rlabel metal2 4094 6494 4094 6494 0 _016_
rlabel metal1 4692 5270 4692 5270 0 _017_
rlabel metal1 5750 6358 5750 6358 0 _018_
rlabel metal2 7774 6494 7774 6494 0 _019_
rlabel metal1 6946 9486 6946 9486 0 _020_
rlabel metal2 8786 9792 8786 9792 0 _021_
rlabel metal1 11178 8840 11178 8840 0 _022_
rlabel metal2 13294 8670 13294 8670 0 _023_
rlabel metal1 2024 10710 2024 10710 0 _024_
rlabel metal2 2714 11424 2714 11424 0 _025_
rlabel metal1 4508 10710 4508 10710 0 _026_
rlabel metal2 5842 10336 5842 10336 0 _027_
rlabel metal1 20470 12750 20470 12750 0 _028_
rlabel metal1 20608 13226 20608 13226 0 _029_
rlabel metal2 13386 3774 13386 3774 0 _030_
rlabel metal1 12834 5168 12834 5168 0 _031_
rlabel metal1 10902 1190 10902 1190 0 _032_
rlabel metal1 7498 1870 7498 1870 0 _033_
rlabel metal2 14122 4012 14122 4012 0 _034_
rlabel metal1 11822 2958 11822 2958 0 _035_
rlabel metal2 14122 7276 14122 7276 0 _036_
rlabel metal2 13478 6154 13478 6154 0 _037_
rlabel metal2 2162 2108 2162 2108 0 _038_
rlabel metal1 3818 1258 3818 1258 0 _039_
rlabel metal1 2668 2482 2668 2482 0 _040_
rlabel metal1 1702 3570 1702 3570 0 _041_
rlabel metal2 3358 4182 3358 4182 0 _042_
rlabel metal1 2254 5746 2254 5746 0 _043_
rlabel metal1 1748 6154 1748 6154 0 _044_
rlabel metal1 3818 7514 3818 7514 0 _045_
rlabel metal2 7130 5372 7130 5372 0 _046_
rlabel metal1 9154 5202 9154 5202 0 _047_
rlabel metal1 11408 6290 11408 6290 0 _048_
rlabel metal1 8694 6766 8694 6766 0 _049_
rlabel metal2 9522 7140 9522 7140 0 _050_
rlabel via1 7679 7378 7679 7378 0 _051_
rlabel metal1 1840 8330 1840 8330 0 _052_
rlabel metal1 3818 6188 3818 6188 0 _053_
rlabel metal1 4370 5100 4370 5100 0 _054_
rlabel metal1 5198 6834 5198 6834 0 _055_
rlabel metal1 7498 6188 7498 6188 0 _056_
rlabel metal1 6164 1938 6164 1938 0 _057_
rlabel metal1 5336 2074 5336 2074 0 _058_
rlabel metal1 9522 3468 9522 3468 0 _059_
rlabel metal1 8648 4522 8648 4522 0 _060_
rlabel metal2 3726 8942 3726 8942 0 _061_
rlabel metal2 4002 9180 4002 9180 0 _062_
rlabel metal2 11178 11356 11178 11356 0 _063_
rlabel metal2 16054 11356 16054 11356 0 _064_
rlabel metal1 9016 8466 9016 8466 0 _065_
rlabel metal2 13386 8092 13386 8092 0 _066_
rlabel metal1 18584 9146 18584 9146 0 _067_
rlabel metal1 15180 8942 15180 8942 0 _068_
rlabel metal1 16100 10030 16100 10030 0 _069_
rlabel metal1 15364 9554 15364 9554 0 _070_
rlabel metal2 11546 10268 11546 10268 0 _071_
rlabel metal1 6256 9486 6256 9486 0 _072_
rlabel metal2 8510 9622 8510 9622 0 _073_
rlabel metal2 11362 9180 11362 9180 0 _074_
rlabel metal2 13018 9452 13018 9452 0 _075_
rlabel metal1 12006 10438 12006 10438 0 _076_
rlabel metal2 11546 12988 11546 12988 0 _077_
rlabel metal1 1932 12410 1932 12410 0 _078_
rlabel metal1 3404 13158 3404 13158 0 _079_
rlabel metal1 5842 11866 5842 11866 0 _080_
rlabel metal2 9062 10880 9062 10880 0 _081_
rlabel metal1 6486 12818 6486 12818 0 _082_
rlabel metal1 4738 13294 4738 13294 0 _083_
rlabel metal1 7544 12750 7544 12750 0 _084_
rlabel metal2 1978 10404 1978 10404 0 _085_
rlabel metal2 3634 10676 3634 10676 0 _086_
rlabel via1 4186 10557 4186 10557 0 _087_
rlabel metal1 5566 10132 5566 10132 0 _088_
rlabel metal1 4922 11084 4922 11084 0 _089_
rlabel metal1 4508 11186 4508 11186 0 _090_
rlabel metal1 12558 8364 12558 8364 0 _091_
rlabel metal2 11086 9180 11086 9180 0 _092_
rlabel metal1 6808 5814 6808 5814 0 _093_
rlabel metal1 6026 6324 6026 6324 0 _094_
rlabel metal1 10166 1870 10166 1870 0 _095_
rlabel metal2 16054 13583 16054 13583 0 clk
rlabel metal1 13340 12410 13340 12410 0 clk_div1_delay.dly\[1\]
rlabel metal1 14122 12818 14122 12818 0 clk_div1_delay.dly\[2\]
rlabel metal2 14766 13124 14766 13124 0 clk_div1_delay.dly\[3\]
rlabel metal1 14904 12818 14904 12818 0 clk_div1_delay.dly\[4\]
rlabel metal2 15502 13124 15502 13124 0 clk_div1_delay.dly\[5\]
rlabel metal1 15640 12818 15640 12818 0 clk_div1_delay.dly\[6\]
rlabel metal1 16192 12954 16192 12954 0 clk_div1_delay.dly\[7\]
rlabel metal2 16698 13022 16698 13022 0 clk_div1_delay.dly\[8\]
rlabel metal1 21482 13253 21482 13253 0 clk_mon
rlabel metal1 21988 12750 21988 12750 0 clk_mon_div\[0\]
rlabel metal1 9936 2550 9936 2550 0 clk_mon_sel[0]
rlabel metal1 12466 5712 12466 5712 0 clk_mon_sel[1]
rlabel metal2 12749 14348 12749 14348 0 clk_mon_sel[2]
rlabel metal1 2530 6256 2530 6256 0 clk_mux1_out
rlabel metal2 2254 6222 2254 6222 0 dll_clk
rlabel metal2 22126 2431 22126 2431 0 hkrst_n
rlabel metal1 3726 1326 3726 1326 0 hsxo
rlabel metal2 15042 1734 15042 1734 0 hsxo_en
rlabel metal2 17526 1316 17526 1316 0 hsxo_en_tf
rlabel metal1 18906 2550 18906 2550 0 hsxo_standby
rlabel metal2 23046 1554 23046 1554 0 hsxo_standby_tf
rlabel metal1 9246 2448 9246 2448 0 lsxo
rlabel metal1 18630 2006 18630 2006 0 lsxo_en
rlabel metal2 19366 1316 19366 1316 0 lsxo_en_tf
rlabel via2 20286 1955 20286 1955 0 lsxo_standby
rlabel metal2 21206 1316 21206 1316 0 lsxo_standby_tf
rlabel metal1 14122 1360 14122 1360 0 net1
rlabel metal1 13439 12886 13439 12886 0 net10
rlabel metal1 13800 2618 13800 2618 0 net11
rlabel metal2 13846 2618 13846 2618 0 net12
rlabel metal1 13846 1870 13846 1870 0 net2
rlabel metal1 21712 13294 21712 13294 0 net3
rlabel metal1 13655 8534 13655 8534 0 net4
rlabel metal2 2898 1632 2898 1632 0 net5
rlabel metal2 8326 1632 8326 1632 0 net6
rlabel metal1 10534 2278 10534 2278 0 net7
rlabel metal2 12650 11628 12650 11628 0 net8
rlabel metal1 13984 2958 13984 2958 0 net9
rlabel metal2 17894 13617 17894 13617 0 pclk
rlabel metal1 16054 12240 16054 12240 0 pclk_div
rlabel metal1 16652 13294 16652 13294 0 pclk_div_skewed_delay.dly\[1\]
rlabel metal1 17020 13158 17020 13158 0 pclk_div_skewed_delay.dly\[2\]
rlabel metal1 17388 12410 17388 12410 0 pclk_div_skewed_delay.dly\[3\]
rlabel metal1 18170 13328 18170 13328 0 pclk_div_skewed_delay.dly\[4\]
rlabel metal2 18630 13022 18630 13022 0 pclk_div_skewed_delay.dly\[5\]
rlabel metal2 12006 1384 12006 1384 0 por_n
rlabel metal1 1702 3434 1702 3434 0 rcosc_16m
rlabel metal2 14214 2244 14214 2244 0 rcosc_16m_en
rlabel metal2 15686 1316 15686 1316 0 rcosc_16m_en_tf
rlabel metal1 13938 2006 13938 2006 0 rcosc_500k
rlabel metal2 2491 14348 2491 14348 0 rcosc_500k_en
rlabel metal2 13846 959 13846 959 0 rcosc_500k_en_tf
rlabel metal2 22218 2380 22218 2380 0 rst_n
rlabel metal2 6210 6137 6210 6137 0 sel_clkdiv0[0]
rlabel via2 7038 7395 7038 7395 0 sel_clkdiv0[1]
rlabel metal3 1142 8228 1142 8228 0 sel_clkdiv0[2]
rlabel metal1 15778 9418 15778 9418 0 sel_clkdiv1[0]
rlabel metal2 13938 10234 13938 10234 0 sel_clkdiv1[1]
rlabel metal1 12719 11594 12719 11594 0 sel_clkdiv1[2]
rlabel metal2 1794 12087 1794 12087 0 sel_clkdiv2[0]
rlabel metal1 5704 13430 5704 13430 0 sel_clkdiv2[1]
rlabel metal3 1717 13124 1717 13124 0 sel_clkdiv2[2]
rlabel metal3 1717 1700 1717 1700 0 sel_mux0
rlabel metal2 1794 1394 1794 1394 0 sel_mux1
rlabel metal1 1794 3944 1794 3944 0 sel_mux2
rlabel metal2 2438 3791 2438 3791 0 sel_mux3
rlabel metal3 1717 4964 1717 4964 0 sel_mux4
rlabel metal3 1004 5780 1004 5780 0 sel_mux5
rlabel metal2 18906 13617 18906 13617 0 usb_clk
rlabel metal1 14858 11696 14858 11696 0 usb_clk_delayed.dly\[1\]
rlabel metal1 16146 11152 16146 11152 0 usb_clk_delayed.dly\[2\]
rlabel metal2 16698 11526 16698 11526 0 usb_clk_delayed.dly\[3\]
rlabel metal1 17434 11696 17434 11696 0 usb_clk_delayed.dly\[4\]
rlabel metal1 18170 11696 18170 11696 0 usb_clk_delayed.dly\[5\]
rlabel metal1 18538 11866 18538 11866 0 usb_clk_delayed.dly\[6\]
rlabel metal1 18446 12240 18446 12240 0 usb_clk_delayed.dly\[7\]
rlabel metal2 18906 11900 18906 11900 0 usb_clk_delayed.dly\[8\]
rlabel metal1 19550 11866 19550 11866 0 usb_clk_delayed.dly\[9\]
rlabel metal2 20233 14348 20233 14348 0 user_clk
rlabel metal1 19550 12206 19550 12206 0 user_clk_delay.dly\[1\]
rlabel metal2 1518 1870 1518 1870 0 xclk
rlabel metal2 10166 1248 10166 1248 0 xrst_n
<< properties >>
string FIXED_BBOX 0 0 24000 15000
<< end >>
