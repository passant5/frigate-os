magic
tech sky130A
magscale 1 2
timestamp 1750134269
<< viali >>
rect 3157 18377 3191 18411
rect 13369 18377 13403 18411
rect 22753 18377 22787 18411
rect 2329 18309 2363 18343
rect 2529 18309 2563 18343
rect 8293 18309 8327 18343
rect 8493 18309 8527 18343
rect 10793 18309 10827 18343
rect 16129 18309 16163 18343
rect 16957 18309 16991 18343
rect 21373 18309 21407 18343
rect 1501 18241 1535 18275
rect 1961 18241 1995 18275
rect 2973 18241 3007 18275
rect 3433 18241 3467 18275
rect 3985 18241 4019 18275
rect 4445 18241 4479 18275
rect 5273 18241 5307 18275
rect 6561 18241 6595 18275
rect 7021 18241 7055 18275
rect 9137 18241 9171 18275
rect 9597 18241 9631 18275
rect 11253 18241 11287 18275
rect 12633 18241 12667 18275
rect 13185 18241 13219 18275
rect 13645 18241 13679 18275
rect 14473 18241 14507 18275
rect 15393 18241 15427 18275
rect 16773 18241 16807 18275
rect 17417 18241 17451 18275
rect 18797 18241 18831 18275
rect 19533 18241 19567 18275
rect 19993 18241 20027 18275
rect 20545 18241 20579 18275
rect 21189 18241 21223 18275
rect 23489 18241 23523 18275
rect 24133 18241 24167 18275
rect 5365 18173 5399 18207
rect 5457 18173 5491 18207
rect 11621 18173 11655 18207
rect 12173 18173 12207 18207
rect 14841 18173 14875 18207
rect 15669 18173 15703 18207
rect 16221 18173 16255 18207
rect 17877 18173 17911 18207
rect 18429 18173 18463 18207
rect 20913 18173 20947 18207
rect 21925 18173 21959 18207
rect 22477 18173 22511 18207
rect 4169 18105 4203 18139
rect 6745 18105 6779 18139
rect 12081 18105 12115 18139
rect 12449 18105 12483 18139
rect 14289 18105 14323 18139
rect 15301 18105 15335 18139
rect 17233 18105 17267 18139
rect 17969 18105 18003 18139
rect 21557 18105 21591 18139
rect 22385 18105 22419 18139
rect 1685 18037 1719 18071
rect 2513 18037 2547 18071
rect 2697 18037 2731 18071
rect 4905 18037 4939 18071
rect 8125 18037 8159 18071
rect 8309 18037 8343 18071
rect 9321 18037 9355 18071
rect 11161 18037 11195 18071
rect 13829 18037 13863 18071
rect 18797 18037 18831 18071
rect 19349 18037 19383 18071
rect 19809 18037 19843 18071
rect 20913 18037 20947 18071
rect 23397 18037 23431 18071
rect 23949 18037 23983 18071
rect 13737 17833 13771 17867
rect 15761 17765 15795 17799
rect 17509 17765 17543 17799
rect 20637 17765 20671 17799
rect 23213 17765 23247 17799
rect 1593 17697 1627 17731
rect 4629 17697 4663 17731
rect 6101 17697 6135 17731
rect 8401 17697 8435 17731
rect 10977 17697 11011 17731
rect 21373 17697 21407 17731
rect 4353 17629 4387 17663
rect 8677 17629 8711 17663
rect 9229 17629 9263 17663
rect 11253 17629 11287 17663
rect 12725 17629 12759 17663
rect 13093 17629 13127 17663
rect 14473 17629 14507 17663
rect 15945 17629 15979 17663
rect 16313 17629 16347 17663
rect 16957 17629 16991 17663
rect 17233 17629 17267 17663
rect 18797 17629 18831 17663
rect 21557 17629 21591 17663
rect 21925 17629 21959 17663
rect 23305 17629 23339 17663
rect 23765 17629 23799 17663
rect 1869 17561 1903 17595
rect 12817 17561 12851 17595
rect 13277 17561 13311 17595
rect 18981 17561 19015 17595
rect 19349 17561 19383 17595
rect 3341 17493 3375 17527
rect 6929 17493 6963 17527
rect 13829 17493 13863 17527
rect 23949 17493 23983 17527
rect 2513 17289 2547 17323
rect 2881 17289 2915 17323
rect 8493 17289 8527 17323
rect 20361 17289 20395 17323
rect 24317 17289 24351 17323
rect 1869 17221 1903 17255
rect 2085 17221 2119 17255
rect 2973 17221 3007 17255
rect 10057 17221 10091 17255
rect 11253 17221 11287 17255
rect 12265 17221 12299 17255
rect 12541 17221 12575 17255
rect 14933 17221 14967 17255
rect 15945 17221 15979 17255
rect 18705 17221 18739 17255
rect 19441 17221 19475 17255
rect 19993 17221 20027 17255
rect 21097 17221 21131 17255
rect 22661 17221 22695 17255
rect 8217 17153 8251 17187
rect 8861 17153 8895 17187
rect 9965 17153 9999 17187
rect 10241 17153 10275 17187
rect 11621 17153 11655 17187
rect 12817 17153 12851 17187
rect 14289 17153 14323 17187
rect 14657 17153 14691 17187
rect 15577 17153 15611 17187
rect 16405 17153 16439 17187
rect 17141 17153 17175 17187
rect 18245 17153 18279 17187
rect 21557 17153 21591 17187
rect 23949 17153 23983 17187
rect 3157 17085 3191 17119
rect 3985 17085 4019 17119
rect 4261 17085 4295 17119
rect 7941 17085 7975 17119
rect 8953 17085 8987 17119
rect 9045 17085 9079 17119
rect 10701 17085 10735 17119
rect 11161 17085 11195 17119
rect 15853 17085 15887 17119
rect 18981 17085 19015 17119
rect 19533 17085 19567 17119
rect 20453 17085 20487 17119
rect 21005 17085 21039 17119
rect 22109 17085 22143 17119
rect 23029 17085 23063 17119
rect 2237 17017 2271 17051
rect 5733 17017 5767 17051
rect 14105 17017 14139 17051
rect 19809 17017 19843 17051
rect 22569 17017 22603 17051
rect 2053 16949 2087 16983
rect 6469 16949 6503 16983
rect 10425 16949 10459 16983
rect 4261 16745 4295 16779
rect 4721 16745 4755 16779
rect 5733 16745 5767 16779
rect 5917 16745 5951 16779
rect 6653 16745 6687 16779
rect 6837 16745 6871 16779
rect 7849 16745 7883 16779
rect 8309 16745 8343 16779
rect 15117 16745 15151 16779
rect 16589 16745 16623 16779
rect 18981 16745 19015 16779
rect 20913 16745 20947 16779
rect 4445 16677 4479 16711
rect 10425 16677 10459 16711
rect 13553 16677 13587 16711
rect 20085 16677 20119 16711
rect 21741 16677 21775 16711
rect 23765 16677 23799 16711
rect 1501 16609 1535 16643
rect 5273 16609 5307 16643
rect 7205 16609 7239 16643
rect 7389 16609 7423 16643
rect 10885 16609 10919 16643
rect 13093 16609 13127 16643
rect 19349 16609 19383 16643
rect 5089 16541 5123 16575
rect 7481 16541 7515 16575
rect 9873 16541 9907 16575
rect 11345 16541 11379 16575
rect 12081 16541 12115 16575
rect 12449 16541 12483 16575
rect 14381 16541 14415 16575
rect 14657 16541 14691 16575
rect 15301 16541 15335 16575
rect 15485 16541 15519 16575
rect 15761 16541 15795 16575
rect 16037 16541 16071 16575
rect 16221 16541 16255 16575
rect 16405 16541 16439 16575
rect 17233 16541 17267 16575
rect 17693 16541 17727 16575
rect 18613 16541 18647 16575
rect 20269 16541 20303 16575
rect 20361 16541 20395 16575
rect 20545 16541 20579 16575
rect 20637 16541 20671 16575
rect 21097 16541 21131 16575
rect 21189 16541 21223 16575
rect 21465 16541 21499 16575
rect 21925 16541 21959 16575
rect 22201 16541 22235 16575
rect 22477 16541 22511 16575
rect 23397 16541 23431 16575
rect 1777 16473 1811 16507
rect 4077 16473 4111 16507
rect 6101 16473 6135 16507
rect 6469 16473 6503 16507
rect 8125 16473 8159 16507
rect 10333 16473 10367 16507
rect 11161 16473 11195 16507
rect 12633 16473 12667 16507
rect 13645 16473 13679 16507
rect 14197 16473 14231 16507
rect 15393 16473 15427 16507
rect 15623 16473 15657 16507
rect 16313 16473 16347 16507
rect 18337 16473 18371 16507
rect 19533 16473 19567 16507
rect 21281 16473 21315 16507
rect 3249 16405 3283 16439
rect 4287 16405 4321 16439
rect 5181 16405 5215 16439
rect 5901 16405 5935 16439
rect 6669 16405 6703 16439
rect 8325 16405 8359 16439
rect 8493 16405 8527 16439
rect 10057 16405 10091 16439
rect 14841 16405 14875 16439
rect 17417 16405 17451 16439
rect 22109 16405 22143 16439
rect 2329 16201 2363 16235
rect 2697 16201 2731 16235
rect 2789 16201 2823 16235
rect 8953 16201 8987 16235
rect 10593 16201 10627 16235
rect 11069 16201 11103 16235
rect 14473 16201 14507 16235
rect 15945 16201 15979 16235
rect 17693 16201 17727 16235
rect 20177 16201 20211 16235
rect 24225 16201 24259 16235
rect 10793 16133 10827 16167
rect 17601 16133 17635 16167
rect 18521 16133 18555 16167
rect 18889 16133 18923 16167
rect 22845 16133 22879 16167
rect 23489 16133 23523 16167
rect 1501 16065 1535 16099
rect 1961 16065 1995 16099
rect 3893 16065 3927 16099
rect 7205 16065 7239 16099
rect 11621 16065 11655 16099
rect 12633 16065 12667 16099
rect 13553 16065 13587 16099
rect 13737 16065 13771 16099
rect 13829 16065 13863 16099
rect 13926 16065 13960 16099
rect 15393 16065 15427 16099
rect 15761 16065 15795 16099
rect 17233 16065 17267 16099
rect 18429 16065 18463 16099
rect 19625 16065 19659 16099
rect 20453 16065 20487 16099
rect 20913 16065 20947 16099
rect 21097 16065 21131 16099
rect 21189 16065 21223 16099
rect 21281 16065 21315 16099
rect 22201 16065 22235 16099
rect 23121 16065 23155 16099
rect 23949 16065 23983 16099
rect 24225 16065 24259 16099
rect 24409 16065 24443 16099
rect 2973 15997 3007 16031
rect 4169 15997 4203 16031
rect 7481 15997 7515 16031
rect 16957 15997 16991 16031
rect 17969 15997 18003 16031
rect 18797 15997 18831 16031
rect 19349 15997 19383 16031
rect 19901 15997 19935 16031
rect 23397 15997 23431 16031
rect 5641 15929 5675 15963
rect 12909 15929 12943 15963
rect 14105 15929 14139 15963
rect 20637 15929 20671 15963
rect 1685 15861 1719 15895
rect 10425 15861 10459 15895
rect 10609 15861 10643 15895
rect 11161 15861 11195 15895
rect 15577 15861 15611 15895
rect 19993 15861 20027 15895
rect 21465 15861 21499 15895
rect 4353 15657 4387 15691
rect 5365 15657 5399 15691
rect 5549 15657 5583 15691
rect 7941 15657 7975 15691
rect 14841 15657 14875 15691
rect 15945 15657 15979 15691
rect 19349 15657 19383 15691
rect 20545 15657 20579 15691
rect 15577 15589 15611 15623
rect 15669 15589 15703 15623
rect 16773 15589 16807 15623
rect 18613 15589 18647 15623
rect 2697 15521 2731 15555
rect 2881 15521 2915 15555
rect 4997 15521 5031 15555
rect 6561 15521 6595 15555
rect 8493 15521 8527 15555
rect 11621 15521 11655 15555
rect 12173 15521 12207 15555
rect 21005 15521 21039 15555
rect 21741 15521 21775 15555
rect 24041 15521 24075 15555
rect 4721 15453 4755 15487
rect 6469 15453 6503 15487
rect 8309 15453 8343 15487
rect 10241 15453 10275 15487
rect 10334 15453 10368 15487
rect 10609 15453 10643 15487
rect 10747 15453 10781 15487
rect 12081 15453 12115 15487
rect 12909 15453 12943 15487
rect 14473 15453 14507 15487
rect 15301 15453 15335 15487
rect 15485 15453 15519 15487
rect 15761 15453 15795 15487
rect 16313 15453 16347 15487
rect 16413 15453 16447 15487
rect 16625 15453 16659 15487
rect 16773 15453 16807 15487
rect 17325 15453 17359 15487
rect 18245 15453 18279 15487
rect 19533 15453 19567 15487
rect 19901 15453 19935 15487
rect 20085 15453 20119 15487
rect 20177 15453 20211 15487
rect 20269 15453 20303 15487
rect 21465 15453 21499 15487
rect 21925 15453 21959 15487
rect 22753 15453 22787 15487
rect 23489 15453 23523 15487
rect 23673 15453 23707 15487
rect 5533 15385 5567 15419
rect 5733 15385 5767 15419
rect 10517 15385 10551 15419
rect 13093 15385 13127 15419
rect 16497 15385 16531 15419
rect 21833 15385 21867 15419
rect 1501 15317 1535 15351
rect 2237 15317 2271 15351
rect 2605 15317 2639 15351
rect 4813 15317 4847 15351
rect 6009 15317 6043 15351
rect 6377 15317 6411 15351
rect 8401 15317 8435 15351
rect 10885 15317 10919 15351
rect 14841 15317 14875 15351
rect 15025 15317 15059 15351
rect 23949 15317 23983 15351
rect 2345 15113 2379 15147
rect 4721 15113 4755 15147
rect 8861 15113 8895 15147
rect 10425 15113 10459 15147
rect 11989 15113 12023 15147
rect 13185 15113 13219 15147
rect 14013 15113 14047 15147
rect 14473 15113 14507 15147
rect 15761 15113 15795 15147
rect 16405 15113 16439 15147
rect 17325 15113 17359 15147
rect 19441 15113 19475 15147
rect 20729 15113 20763 15147
rect 21557 15113 21591 15147
rect 22569 15113 22603 15147
rect 2145 15045 2179 15079
rect 5641 15045 5675 15079
rect 5857 15045 5891 15079
rect 12909 15045 12943 15079
rect 15485 15045 15519 15079
rect 18245 15045 18279 15079
rect 18429 15045 18463 15079
rect 23397 15045 23431 15079
rect 23673 15045 23707 15079
rect 1501 14977 1535 15011
rect 2973 14977 3007 15011
rect 7113 14977 7147 15011
rect 9781 14977 9815 15011
rect 9873 14977 9907 15011
rect 10057 14977 10091 15011
rect 10149 14977 10183 15011
rect 10701 14977 10735 15011
rect 11161 14977 11195 15011
rect 11621 14977 11655 15011
rect 11805 14977 11839 15011
rect 12081 14977 12115 15011
rect 12541 14977 12575 15011
rect 12699 14977 12733 15011
rect 12817 14977 12851 15011
rect 13001 14977 13035 15011
rect 13645 14977 13679 15011
rect 13875 14977 13909 15011
rect 14197 14977 14231 15011
rect 14841 14977 14875 15011
rect 15117 14977 15151 15011
rect 16129 14977 16163 15011
rect 16221 14977 16255 15011
rect 16773 14977 16807 15011
rect 16957 14977 16991 15011
rect 17049 14977 17083 15011
rect 17141 14977 17175 15011
rect 17785 14977 17819 15011
rect 19165 14977 19199 15011
rect 19625 14977 19659 15011
rect 20085 14977 20119 15011
rect 20269 14977 20303 15011
rect 20361 14977 20395 15011
rect 20453 14977 20487 15011
rect 21005 14977 21039 15011
rect 21189 14977 21223 15011
rect 21281 14977 21315 15011
rect 21373 14977 21407 15011
rect 21925 14977 21959 15011
rect 22018 14977 22052 15011
rect 22201 14977 22235 15011
rect 22293 14977 22327 15011
rect 22390 14977 22424 15011
rect 23305 14977 23339 15011
rect 23857 14977 23891 15011
rect 24409 14977 24443 15011
rect 3249 14909 3283 14943
rect 7389 14909 7423 14943
rect 14105 14909 14139 14943
rect 14749 14909 14783 14943
rect 15393 14909 15427 14943
rect 15602 14909 15636 14943
rect 22845 14909 22879 14943
rect 1685 14841 1719 14875
rect 9597 14841 9631 14875
rect 10885 14841 10919 14875
rect 17969 14841 18003 14875
rect 2329 14773 2363 14807
rect 2513 14773 2547 14807
rect 5825 14773 5859 14807
rect 6009 14773 6043 14807
rect 10793 14773 10827 14807
rect 10977 14773 11011 14807
rect 13645 14773 13679 14807
rect 14841 14773 14875 14807
rect 24225 14773 24259 14807
rect 3893 14569 3927 14603
rect 7389 14569 7423 14603
rect 7573 14569 7607 14603
rect 7849 14569 7883 14603
rect 9321 14569 9355 14603
rect 9873 14569 9907 14603
rect 11713 14569 11747 14603
rect 12633 14569 12667 14603
rect 16957 14569 16991 14603
rect 17325 14569 17359 14603
rect 21097 14569 21131 14603
rect 21557 14569 21591 14603
rect 11069 14501 11103 14535
rect 11989 14501 12023 14535
rect 16037 14501 16071 14535
rect 23765 14501 23799 14535
rect 1501 14433 1535 14467
rect 4537 14433 4571 14467
rect 4997 14433 5031 14467
rect 8401 14433 8435 14467
rect 15393 14433 15427 14467
rect 19349 14433 19383 14467
rect 19901 14433 19935 14467
rect 4261 14365 4295 14399
rect 8217 14365 8251 14399
rect 10005 14365 10039 14399
rect 10425 14365 10459 14399
rect 10977 14365 11011 14399
rect 11161 14365 11195 14399
rect 11253 14365 11287 14399
rect 11437 14365 11471 14399
rect 11897 14365 11931 14399
rect 12081 14365 12115 14399
rect 12173 14365 12207 14399
rect 12541 14365 12575 14399
rect 12725 14365 12759 14399
rect 13001 14365 13035 14399
rect 13277 14365 13311 14399
rect 14565 14365 14599 14399
rect 14933 14365 14967 14399
rect 15117 14365 15151 14399
rect 15301 14365 15335 14399
rect 16221 14365 16255 14399
rect 16543 14365 16577 14399
rect 16681 14365 16715 14399
rect 16957 14365 16991 14399
rect 17141 14365 17175 14399
rect 17877 14365 17911 14399
rect 20361 14365 20395 14399
rect 20913 14365 20947 14399
rect 21373 14365 21407 14399
rect 21833 14365 21867 14399
rect 22293 14365 22327 14399
rect 23213 14365 23247 14399
rect 1777 14297 1811 14331
rect 5273 14297 5307 14331
rect 7205 14297 7239 14331
rect 8309 14297 8343 14331
rect 9289 14297 9323 14331
rect 9505 14297 9539 14331
rect 10149 14297 10183 14331
rect 10241 14297 10275 14331
rect 10701 14297 10735 14331
rect 16313 14297 16347 14331
rect 16405 14297 16439 14331
rect 18521 14297 18555 14331
rect 18797 14297 18831 14331
rect 19441 14297 19475 14331
rect 3249 14229 3283 14263
rect 4353 14229 4387 14263
rect 6745 14229 6779 14263
rect 7415 14229 7449 14263
rect 9137 14229 9171 14263
rect 13093 14229 13127 14263
rect 13461 14229 13495 14263
rect 20177 14229 20211 14263
rect 22017 14229 22051 14263
rect 3341 14025 3375 14059
rect 3985 14025 4019 14059
rect 6469 14025 6503 14059
rect 6637 14025 6671 14059
rect 8861 14025 8895 14059
rect 9337 14025 9371 14059
rect 13343 14025 13377 14059
rect 14841 14025 14875 14059
rect 15669 14025 15703 14059
rect 16773 14025 16807 14059
rect 20085 14025 20119 14059
rect 21097 14025 21131 14059
rect 3617 13957 3651 13991
rect 3833 13957 3867 13991
rect 6837 13957 6871 13991
rect 9137 13957 9171 13991
rect 11161 13957 11195 13991
rect 19441 13957 19475 13991
rect 20637 13957 20671 13991
rect 22017 13957 22051 13991
rect 22569 13957 22603 13991
rect 22845 13957 22879 13991
rect 23765 13957 23799 13991
rect 23857 13957 23891 13991
rect 1593 13889 1627 13923
rect 6101 13889 6135 13923
rect 7113 13889 7147 13923
rect 10057 13889 10091 13923
rect 10241 13889 10275 13923
rect 10517 13889 10551 13923
rect 10793 13889 10827 13923
rect 11897 13889 11931 13923
rect 11989 13889 12023 13923
rect 12265 13889 12299 13923
rect 13277 13889 13311 13923
rect 13921 13889 13955 13923
rect 14105 13889 14139 13923
rect 14841 13889 14875 13923
rect 15025 13889 15059 13923
rect 15209 13889 15243 13923
rect 16037 13889 16071 13923
rect 16957 13889 16991 13923
rect 17141 13889 17175 13923
rect 17233 13889 17267 13923
rect 17601 13889 17635 13923
rect 17877 13889 17911 13923
rect 19349 13889 19383 13923
rect 19901 13889 19935 13923
rect 21557 13889 21591 13923
rect 22201 13889 22235 13923
rect 23489 13889 23523 13923
rect 1869 13821 1903 13855
rect 7389 13821 7423 13855
rect 10701 13821 10735 13855
rect 10885 13821 10919 13855
rect 10977 13821 11011 13855
rect 15945 13821 15979 13855
rect 19717 13821 19751 13855
rect 24317 13821 24351 13855
rect 11621 13753 11655 13787
rect 3801 13685 3835 13719
rect 4353 13685 4387 13719
rect 5843 13685 5877 13719
rect 6653 13685 6687 13719
rect 9321 13685 9355 13719
rect 9505 13685 9539 13719
rect 10149 13685 10183 13719
rect 11805 13685 11839 13719
rect 12357 13685 12391 13719
rect 15853 13685 15887 13719
rect 20545 13685 20579 13719
rect 21465 13685 21499 13719
rect 2053 13481 2087 13515
rect 2237 13481 2271 13515
rect 6193 13481 6227 13515
rect 7849 13481 7883 13515
rect 9321 13481 9355 13515
rect 11713 13481 11747 13515
rect 12817 13481 12851 13515
rect 16589 13481 16623 13515
rect 16957 13481 16991 13515
rect 2513 13413 2547 13447
rect 18797 13413 18831 13447
rect 21005 13413 21039 13447
rect 22661 13413 22695 13447
rect 3157 13345 3191 13379
rect 5549 13345 5583 13379
rect 5733 13345 5767 13379
rect 8493 13345 8527 13379
rect 10241 13345 10275 13379
rect 12541 13345 12575 13379
rect 16681 13345 16715 13379
rect 18337 13345 18371 13379
rect 20085 13345 20119 13379
rect 21097 13345 21131 13379
rect 23213 13345 23247 13379
rect 2881 13277 2915 13311
rect 8217 13277 8251 13311
rect 9781 13277 9815 13311
rect 9965 13277 9999 13311
rect 11069 13277 11103 13311
rect 12633 13277 12667 13311
rect 13369 13277 13403 13311
rect 13645 13277 13679 13311
rect 13829 13277 13863 13311
rect 15577 13277 15611 13311
rect 16037 13277 16071 13311
rect 16313 13277 16347 13311
rect 16589 13277 16623 13311
rect 17969 13277 18003 13311
rect 19533 13277 19567 13311
rect 20545 13277 20579 13311
rect 21373 13277 21407 13311
rect 22845 13277 22879 13311
rect 23765 13277 23799 13311
rect 1869 13209 1903 13243
rect 5825 13209 5859 13243
rect 8309 13209 8343 13243
rect 9305 13209 9339 13243
rect 9505 13209 9539 13243
rect 10793 13209 10827 13243
rect 11697 13209 11731 13243
rect 11897 13209 11931 13243
rect 18061 13209 18095 13243
rect 18889 13209 18923 13243
rect 19993 13209 20027 13243
rect 23673 13209 23707 13243
rect 1501 13141 1535 13175
rect 2069 13141 2103 13175
rect 2973 13141 3007 13175
rect 9137 13141 9171 13175
rect 11161 13141 11195 13175
rect 11529 13141 11563 13175
rect 12173 13141 12207 13175
rect 15025 13141 15059 13175
rect 24133 13141 24167 13175
rect 1685 12937 1719 12971
rect 10977 12937 11011 12971
rect 12633 12937 12667 12971
rect 18521 12937 18555 12971
rect 2053 12869 2087 12903
rect 2253 12869 2287 12903
rect 3065 12869 3099 12903
rect 3877 12869 3911 12903
rect 4077 12869 4111 12903
rect 5733 12869 5767 12903
rect 5933 12869 5967 12903
rect 10241 12869 10275 12903
rect 15393 12869 15427 12903
rect 24225 12869 24259 12903
rect 1501 12801 1535 12835
rect 7941 12801 7975 12835
rect 11621 12801 11655 12835
rect 11713 12801 11747 12835
rect 11897 12801 11931 12835
rect 12081 12801 12115 12835
rect 12817 12801 12851 12835
rect 12909 12801 12943 12835
rect 13002 12801 13036 12835
rect 14013 12801 14047 12835
rect 14657 12801 14691 12835
rect 14749 12801 14783 12835
rect 14933 12801 14967 12835
rect 15577 12801 15611 12835
rect 15761 12801 15795 12835
rect 16405 12801 16439 12835
rect 16773 12801 16807 12835
rect 18889 12801 18923 12835
rect 20361 12801 20395 12835
rect 21925 12801 21959 12835
rect 22569 12801 22603 12835
rect 22845 12801 22879 12835
rect 23673 12801 23707 12835
rect 23949 12801 23983 12835
rect 3157 12733 3191 12767
rect 3341 12733 3375 12767
rect 8217 12733 8251 12767
rect 8493 12733 8527 12767
rect 10517 12733 10551 12767
rect 13093 12733 13127 12767
rect 14105 12733 14139 12767
rect 16221 12733 16255 12767
rect 17049 12733 17083 12767
rect 20729 12733 20763 12767
rect 21281 12733 21315 12767
rect 23121 12733 23155 12767
rect 2421 12665 2455 12699
rect 16037 12665 16071 12699
rect 16313 12665 16347 12699
rect 20361 12665 20395 12699
rect 21189 12665 21223 12699
rect 23213 12665 23247 12699
rect 2237 12597 2271 12631
rect 2697 12597 2731 12631
rect 3709 12597 3743 12631
rect 3893 12597 3927 12631
rect 5917 12597 5951 12631
rect 6101 12597 6135 12631
rect 7757 12597 7791 12631
rect 14381 12597 14415 12631
rect 15117 12597 15151 12631
rect 16221 12597 16255 12631
rect 9597 12393 9631 12427
rect 15393 12393 15427 12427
rect 15853 12393 15887 12427
rect 16313 12393 16347 12427
rect 17141 12393 17175 12427
rect 17785 12393 17819 12427
rect 21465 12393 21499 12427
rect 17325 12325 17359 12359
rect 23765 12325 23799 12359
rect 1777 12257 1811 12291
rect 4353 12257 4387 12291
rect 4445 12257 4479 12291
rect 4905 12257 4939 12291
rect 7481 12257 7515 12291
rect 8125 12257 8159 12291
rect 10057 12257 10091 12291
rect 11161 12257 11195 12291
rect 13277 12257 13311 12291
rect 13369 12257 13403 12291
rect 15945 12257 15979 12291
rect 18613 12257 18647 12291
rect 21189 12257 21223 12291
rect 21281 12257 21315 12291
rect 22109 12257 22143 12291
rect 1501 12189 1535 12223
rect 4261 12189 4295 12223
rect 7297 12189 7331 12223
rect 8401 12189 8435 12223
rect 9873 12189 9907 12223
rect 10333 12189 10367 12223
rect 11989 12189 12023 12223
rect 12265 12189 12299 12223
rect 12541 12189 12575 12223
rect 12633 12189 12667 12223
rect 13461 12189 13495 12223
rect 13553 12189 13587 12223
rect 14749 12189 14783 12223
rect 14933 12189 14967 12223
rect 15025 12189 15059 12223
rect 15117 12189 15151 12223
rect 15669 12189 15703 12223
rect 15761 12189 15795 12223
rect 16405 12189 16439 12223
rect 18337 12189 18371 12223
rect 19349 12189 19383 12223
rect 19993 12189 20027 12223
rect 20269 12189 20303 12223
rect 21005 12189 21039 12223
rect 21097 12189 21131 12223
rect 21741 12189 21775 12223
rect 21925 12189 21959 12223
rect 22477 12189 22511 12223
rect 23857 12189 23891 12223
rect 5181 12121 5215 12155
rect 7389 12121 7423 12155
rect 9505 12121 9539 12155
rect 10425 12121 10459 12155
rect 10609 12121 10643 12155
rect 12449 12121 12483 12155
rect 16957 12121 16991 12155
rect 17601 12121 17635 12155
rect 3249 12053 3283 12087
rect 3893 12053 3927 12087
rect 6653 12053 6687 12087
rect 6929 12053 6963 12087
rect 10333 12053 10367 12087
rect 12817 12053 12851 12087
rect 13737 12053 13771 12087
rect 17167 12053 17201 12087
rect 17801 12053 17835 12087
rect 17969 12053 18003 12087
rect 4077 11849 4111 11883
rect 4997 11849 5031 11883
rect 5365 11849 5399 11883
rect 5733 11849 5767 11883
rect 6637 11849 6671 11883
rect 10517 11849 10551 11883
rect 15209 11849 15243 11883
rect 19717 11849 19751 11883
rect 20913 11849 20947 11883
rect 22477 11849 22511 11883
rect 2605 11781 2639 11815
rect 6837 11781 6871 11815
rect 7389 11781 7423 11815
rect 9965 11781 9999 11815
rect 10057 11781 10091 11815
rect 14841 11781 14875 11815
rect 20269 11781 20303 11815
rect 20386 11781 20420 11815
rect 22109 11781 22143 11815
rect 23857 11781 23891 11815
rect 24133 11781 24167 11815
rect 1501 11713 1535 11747
rect 1961 11713 1995 11747
rect 4813 11713 4847 11747
rect 9689 11713 9723 11747
rect 10333 11713 10367 11747
rect 11621 11713 11655 11747
rect 11989 11713 12023 11747
rect 12081 11713 12115 11747
rect 13185 11713 13219 11747
rect 13369 11713 13403 11747
rect 13645 11713 13679 11747
rect 14381 11713 14415 11747
rect 14749 11713 14783 11747
rect 15117 11713 15151 11747
rect 15393 11713 15427 11747
rect 15853 11713 15887 11747
rect 16037 11713 16071 11747
rect 20186 11719 20220 11753
rect 20499 11713 20533 11747
rect 20637 11713 20671 11747
rect 21465 11713 21499 11747
rect 21925 11713 21959 11747
rect 22201 11713 22235 11747
rect 22293 11713 22327 11747
rect 22937 11713 22971 11747
rect 23581 11713 23615 11747
rect 24317 11713 24351 11747
rect 2329 11645 2363 11679
rect 5825 11645 5859 11679
rect 5917 11645 5951 11679
rect 7113 11645 7147 11679
rect 9873 11645 9907 11679
rect 10793 11645 10827 11679
rect 10885 11645 10919 11679
rect 13553 11645 13587 11679
rect 14657 11645 14691 11679
rect 17233 11645 17267 11679
rect 17509 11645 17543 11679
rect 18981 11645 19015 11679
rect 19993 11645 20027 11679
rect 21189 11645 21223 11679
rect 1685 11577 1719 11611
rect 6469 11509 6503 11543
rect 6653 11509 6687 11543
rect 8861 11509 8895 11543
rect 14473 11509 14507 11543
rect 15577 11509 15611 11543
rect 16037 11509 16071 11543
rect 19625 11509 19659 11543
rect 21373 11509 21407 11543
rect 2053 11305 2087 11339
rect 4537 11305 4571 11339
rect 4905 11305 4939 11339
rect 7389 11305 7423 11339
rect 9321 11305 9355 11339
rect 13645 11305 13679 11339
rect 19901 11305 19935 11339
rect 22753 11305 22787 11339
rect 2237 11237 2271 11271
rect 8401 11237 8435 11271
rect 11253 11237 11287 11271
rect 22293 11237 22327 11271
rect 3157 11169 3191 11203
rect 6377 11169 6411 11203
rect 7941 11169 7975 11203
rect 11069 11169 11103 11203
rect 13461 11169 13495 11203
rect 15117 11169 15151 11203
rect 16681 11169 16715 11203
rect 19625 11169 19659 11203
rect 21097 11169 21131 11203
rect 23029 11169 23063 11203
rect 23857 11169 23891 11203
rect 2973 11101 3007 11135
rect 4353 11101 4387 11135
rect 6653 11101 6687 11135
rect 7757 11101 7791 11135
rect 9045 11101 9079 11135
rect 9321 11101 9355 11135
rect 9781 11101 9815 11135
rect 9873 11101 9907 11135
rect 10241 11101 10275 11135
rect 10793 11101 10827 11135
rect 11437 11101 11471 11135
rect 11805 11101 11839 11135
rect 12357 11101 12391 11135
rect 13277 11101 13311 11135
rect 13369 11101 13403 11135
rect 13645 11101 13679 11135
rect 15853 11101 15887 11135
rect 16037 11101 16071 11135
rect 16129 11101 16163 11135
rect 19717 11101 19751 11135
rect 20453 11101 20487 11135
rect 20637 11101 20671 11135
rect 20729 11101 20763 11135
rect 20821 11101 20855 11135
rect 21649 11101 21683 11135
rect 21742 11101 21776 11135
rect 21925 11101 21959 11135
rect 22155 11101 22189 11135
rect 22569 11101 22603 11135
rect 24041 11101 24075 11135
rect 1869 11033 1903 11067
rect 2069 11033 2103 11067
rect 8585 11033 8619 11067
rect 9137 11033 9171 11067
rect 9597 11033 9631 11067
rect 12909 11033 12943 11067
rect 15301 11033 15335 11067
rect 16957 11033 16991 11067
rect 18705 11033 18739 11067
rect 22017 11033 22051 11067
rect 23489 11033 23523 11067
rect 23581 11033 23615 11067
rect 2513 10965 2547 10999
rect 2881 10965 2915 10999
rect 7849 10965 7883 10999
rect 10057 10965 10091 10999
rect 10149 10965 10183 10999
rect 15669 10965 15703 10999
rect 3433 10761 3467 10795
rect 7773 10761 7807 10795
rect 10885 10761 10919 10795
rect 16313 10761 16347 10795
rect 18797 10761 18831 10795
rect 20637 10761 20671 10795
rect 21557 10761 21591 10795
rect 24041 10761 24075 10795
rect 1961 10693 1995 10727
rect 7573 10693 7607 10727
rect 8217 10693 8251 10727
rect 10977 10693 11011 10727
rect 11897 10693 11931 10727
rect 15209 10693 15243 10727
rect 20545 10693 20579 10727
rect 22293 10693 22327 10727
rect 23489 10693 23523 10727
rect 6653 10625 6687 10659
rect 8401 10625 8435 10659
rect 8493 10625 8527 10659
rect 9781 10625 9815 10659
rect 11253 10625 11287 10659
rect 12449 10625 12483 10659
rect 13001 10625 13035 10659
rect 13737 10625 13771 10659
rect 14473 10625 14507 10659
rect 15577 10625 15611 10659
rect 16037 10625 16071 10659
rect 16129 10625 16163 10659
rect 16405 10625 16439 10659
rect 21465 10625 21499 10659
rect 23397 10625 23431 10659
rect 24225 10625 24259 10659
rect 1685 10557 1719 10591
rect 4077 10557 4111 10591
rect 5825 10557 5859 10591
rect 6101 10557 6135 10591
rect 6929 10557 6963 10591
rect 9137 10557 9171 10591
rect 10768 10557 10802 10591
rect 12909 10557 12943 10591
rect 16221 10557 16255 10591
rect 17049 10557 17083 10591
rect 17325 10557 17359 10591
rect 22385 10557 22419 10591
rect 22569 10557 22603 10591
rect 23581 10557 23615 10591
rect 8217 10489 8251 10523
rect 10609 10489 10643 10523
rect 6469 10421 6503 10455
rect 6837 10421 6871 10455
rect 7757 10421 7791 10455
rect 7941 10421 7975 10455
rect 13369 10421 13403 10455
rect 21925 10421 21959 10455
rect 23029 10421 23063 10455
rect 4261 10217 4295 10251
rect 4905 10217 4939 10251
rect 5089 10217 5123 10251
rect 5365 10217 5399 10251
rect 12633 10217 12667 10251
rect 13369 10217 13403 10251
rect 15025 10217 15059 10251
rect 17693 10217 17727 10251
rect 17877 10217 17911 10251
rect 18337 10217 18371 10251
rect 18521 10217 18555 10251
rect 23397 10217 23431 10251
rect 24133 10217 24167 10251
rect 13185 10149 13219 10183
rect 14749 10149 14783 10183
rect 1961 10081 1995 10115
rect 5825 10081 5859 10115
rect 8677 10081 8711 10115
rect 15301 10081 15335 10115
rect 20821 10081 20855 10115
rect 21649 10081 21683 10115
rect 1685 10013 1719 10047
rect 4445 10013 4479 10047
rect 5549 10013 5583 10047
rect 5641 10013 5675 10047
rect 5733 10013 5767 10047
rect 6653 10013 6687 10047
rect 9045 10013 9079 10047
rect 11253 10013 11287 10047
rect 11713 10013 11747 10047
rect 12081 10013 12115 10047
rect 12909 10013 12943 10047
rect 14565 10013 14599 10047
rect 14657 10013 14691 10047
rect 14841 10013 14875 10047
rect 15393 10013 15427 10047
rect 16319 10013 16353 10047
rect 16497 10013 16531 10047
rect 20729 10013 20763 10047
rect 23673 10013 23707 10047
rect 23765 10013 23799 10047
rect 23949 10013 23983 10047
rect 4721 9945 4755 9979
rect 6929 9945 6963 9979
rect 9321 9945 9355 9979
rect 13553 9945 13587 9979
rect 16405 9945 16439 9979
rect 17509 9945 17543 9979
rect 18153 9945 18187 9979
rect 21925 9945 21959 9979
rect 3433 9877 3467 9911
rect 4921 9877 4955 9911
rect 10793 9877 10827 9911
rect 13343 9877 13377 9911
rect 17709 9877 17743 9911
rect 18353 9877 18387 9911
rect 20269 9877 20303 9911
rect 20637 9877 20671 9911
rect 21373 9877 21407 9911
rect 2237 9673 2271 9707
rect 2513 9673 2547 9707
rect 2881 9673 2915 9707
rect 6929 9673 6963 9707
rect 12633 9673 12667 9707
rect 15577 9673 15611 9707
rect 18965 9673 18999 9707
rect 1869 9605 1903 9639
rect 2069 9605 2103 9639
rect 8953 9605 8987 9639
rect 9153 9605 9187 9639
rect 9597 9605 9631 9639
rect 17141 9605 17175 9639
rect 18245 9605 18279 9639
rect 19165 9605 19199 9639
rect 22093 9605 22127 9639
rect 22293 9605 22327 9639
rect 22845 9605 22879 9639
rect 6469 9537 6503 9571
rect 6653 9537 6687 9571
rect 7113 9537 7147 9571
rect 9781 9537 9815 9571
rect 10793 9537 10827 9571
rect 10885 9537 10919 9571
rect 10977 9537 11011 9571
rect 11805 9537 11839 9571
rect 11897 9537 11931 9571
rect 13001 9537 13035 9571
rect 14013 9537 14047 9571
rect 14381 9537 14415 9571
rect 14473 9537 14507 9571
rect 14933 9537 14967 9571
rect 15577 9537 15611 9571
rect 16037 9537 16071 9571
rect 16221 9537 16255 9571
rect 18153 9537 18187 9571
rect 19717 9537 19751 9571
rect 22569 9537 22603 9571
rect 2973 9469 3007 9503
rect 3157 9469 3191 9503
rect 4261 9469 4295 9503
rect 4537 9469 4571 9503
rect 6009 9469 6043 9503
rect 7389 9469 7423 9503
rect 11253 9469 11287 9503
rect 12357 9469 12391 9503
rect 15209 9469 15243 9503
rect 15761 9469 15795 9503
rect 17233 9469 17267 9503
rect 17417 9469 17451 9503
rect 18337 9469 18371 9503
rect 19993 9469 20027 9503
rect 21465 9469 21499 9503
rect 24317 9469 24351 9503
rect 9321 9401 9355 9435
rect 11161 9401 11195 9435
rect 13921 9401 13955 9435
rect 14749 9401 14783 9435
rect 16129 9401 16163 9435
rect 21925 9401 21959 9435
rect 2053 9333 2087 9367
rect 6469 9333 6503 9367
rect 7297 9333 7331 9367
rect 9137 9333 9171 9367
rect 10517 9333 10551 9367
rect 12265 9333 12299 9367
rect 13461 9333 13495 9367
rect 14841 9333 14875 9367
rect 16773 9333 16807 9367
rect 17785 9333 17819 9367
rect 18797 9333 18831 9367
rect 18981 9333 19015 9367
rect 22109 9333 22143 9367
rect 4813 9129 4847 9163
rect 4997 9129 5031 9163
rect 5273 9129 5307 9163
rect 8401 9129 8435 9163
rect 9505 9129 9539 9163
rect 9735 9129 9769 9163
rect 18061 9129 18095 9163
rect 18521 9129 18555 9163
rect 22109 9129 22143 9163
rect 22569 9129 22603 9163
rect 22753 9129 22787 9163
rect 23305 9129 23339 9163
rect 23489 9129 23523 9163
rect 23949 9129 23983 9163
rect 9597 9061 9631 9095
rect 7021 8993 7055 9027
rect 10333 8993 10367 9027
rect 12173 8993 12207 9027
rect 16313 8993 16347 9027
rect 19349 8993 19383 9027
rect 1593 8925 1627 8959
rect 5457 8925 5491 8959
rect 5549 8925 5583 8959
rect 5779 8925 5813 8959
rect 5917 8925 5951 8959
rect 6193 8925 6227 8959
rect 6377 8925 6411 8959
rect 6653 8925 6687 8959
rect 7481 8925 7515 8959
rect 9413 8925 9447 8959
rect 9873 8925 9907 8959
rect 10236 8925 10270 8959
rect 10977 8925 11011 8959
rect 11897 8925 11931 8959
rect 13093 8925 13127 8959
rect 14197 8925 14231 8959
rect 21649 8925 21683 8959
rect 21925 8925 21959 8959
rect 24133 8925 24167 8959
rect 1869 8857 1903 8891
rect 4629 8857 4663 8891
rect 4845 8857 4879 8891
rect 5641 8857 5675 8891
rect 7159 8857 7193 8891
rect 7297 8857 7331 8891
rect 7389 8857 7423 8891
rect 8217 8857 8251 8891
rect 8433 8857 8467 8891
rect 10333 8857 10367 8891
rect 10425 8857 10459 8891
rect 10609 8857 10643 8891
rect 11529 8857 11563 8891
rect 13645 8857 13679 8891
rect 14473 8857 14507 8891
rect 16589 8857 16623 8891
rect 18705 8857 18739 8891
rect 19625 8857 19659 8891
rect 22385 8857 22419 8891
rect 23121 8857 23155 8891
rect 23337 8857 23371 8891
rect 3341 8789 3375 8823
rect 6561 8789 6595 8823
rect 7665 8789 7699 8823
rect 8585 8789 8619 8823
rect 15945 8789 15979 8823
rect 18337 8789 18371 8823
rect 18505 8789 18539 8823
rect 21097 8789 21131 8823
rect 21465 8789 21499 8823
rect 22595 8789 22629 8823
rect 2145 8585 2179 8619
rect 2421 8585 2455 8619
rect 2789 8585 2823 8619
rect 9965 8585 9999 8619
rect 14381 8585 14415 8619
rect 15209 8585 15243 8619
rect 18705 8585 18739 8619
rect 19349 8585 19383 8619
rect 19717 8585 19751 8619
rect 20361 8585 20395 8619
rect 20529 8585 20563 8619
rect 21215 8585 21249 8619
rect 24199 8585 24233 8619
rect 1777 8517 1811 8551
rect 1993 8517 2027 8551
rect 5733 8517 5767 8551
rect 5933 8517 5967 8551
rect 7757 8517 7791 8551
rect 15377 8517 15411 8551
rect 15577 8517 15611 8551
rect 17233 8517 17267 8551
rect 19809 8517 19843 8551
rect 20729 8517 20763 8551
rect 21005 8517 21039 8551
rect 24409 8517 24443 8551
rect 2881 8449 2915 8483
rect 3433 8449 3467 8483
rect 3893 8449 3927 8483
rect 6837 8449 6871 8483
rect 6929 8449 6963 8483
rect 7021 8449 7055 8483
rect 7481 8449 7515 8483
rect 9781 8449 9815 8483
rect 9965 8449 9999 8483
rect 10425 8449 10459 8483
rect 10517 8449 10551 8483
rect 10793 8449 10827 8483
rect 10885 8449 10919 8483
rect 11713 8449 11747 8483
rect 11897 8449 11931 8483
rect 12081 8449 12115 8483
rect 12357 8449 12391 8483
rect 12909 8449 12943 8483
rect 14749 8449 14783 8483
rect 15853 8449 15887 8483
rect 22017 8449 22051 8483
rect 3065 8381 3099 8415
rect 6745 8381 6779 8415
rect 7205 8381 7239 8415
rect 9229 8381 9263 8415
rect 13001 8381 13035 8415
rect 14105 8381 14139 8415
rect 14657 8381 14691 8415
rect 16129 8381 16163 8415
rect 16957 8381 16991 8415
rect 19901 8381 19935 8415
rect 22293 8381 22327 8415
rect 3617 8313 3651 8347
rect 11621 8313 11655 8347
rect 15853 8313 15887 8347
rect 15945 8313 15979 8347
rect 18981 8313 19015 8347
rect 21373 8313 21407 8347
rect 23765 8313 23799 8347
rect 24041 8313 24075 8347
rect 1961 8245 1995 8279
rect 5917 8245 5951 8279
rect 6101 8245 6135 8279
rect 13277 8245 13311 8279
rect 13645 8245 13679 8279
rect 15393 8245 15427 8279
rect 20545 8245 20579 8279
rect 21189 8245 21223 8279
rect 24225 8245 24259 8279
rect 1685 8041 1719 8075
rect 6745 8041 6779 8075
rect 10609 8041 10643 8075
rect 13001 8041 13035 8075
rect 13829 8041 13863 8075
rect 17141 8041 17175 8075
rect 18797 8041 18831 8075
rect 22937 8041 22971 8075
rect 12265 7973 12299 8007
rect 2881 7905 2915 7939
rect 3065 7905 3099 7939
rect 3893 7905 3927 7939
rect 5917 7905 5951 7939
rect 7481 7905 7515 7939
rect 10149 7905 10183 7939
rect 10517 7905 10551 7939
rect 14473 7905 14507 7939
rect 18245 7905 18279 7939
rect 19901 7905 19935 7939
rect 21097 7905 21131 7939
rect 22017 7905 22051 7939
rect 23397 7905 23431 7939
rect 23489 7905 23523 7939
rect 1501 7837 1535 7871
rect 2145 7837 2179 7871
rect 6469 7837 6503 7871
rect 6748 7837 6782 7871
rect 7205 7837 7239 7871
rect 7297 7837 7331 7871
rect 7389 7837 7423 7871
rect 8309 7837 8343 7871
rect 8401 7837 8435 7871
rect 8493 7837 8527 7871
rect 9045 7837 9079 7871
rect 9229 7837 9263 7871
rect 9321 7837 9355 7871
rect 9413 7837 9447 7871
rect 10057 7837 10091 7871
rect 10241 7837 10275 7871
rect 10793 7837 10827 7871
rect 11069 7837 11103 7871
rect 11621 7837 11655 7871
rect 11805 7837 11839 7871
rect 11897 7837 11931 7871
rect 11989 7837 12023 7871
rect 13185 7837 13219 7871
rect 13277 7837 13311 7871
rect 13645 7837 13679 7871
rect 13829 7837 13863 7871
rect 14197 7837 14231 7871
rect 16773 7837 16807 7871
rect 17325 7837 17359 7871
rect 17969 7837 18003 7871
rect 22201 7837 22235 7871
rect 23305 7837 23339 7871
rect 24133 7837 24167 7871
rect 3433 7769 3467 7803
rect 5641 7769 5675 7803
rect 8677 7769 8711 7803
rect 11345 7769 11379 7803
rect 18765 7769 18799 7803
rect 18981 7769 19015 7803
rect 19717 7769 19751 7803
rect 21005 7769 21039 7803
rect 22293 7769 22327 7803
rect 2053 7701 2087 7735
rect 2421 7701 2455 7735
rect 2789 7701 2823 7735
rect 6561 7701 6595 7735
rect 7021 7701 7055 7735
rect 9689 7701 9723 7735
rect 15945 7701 15979 7735
rect 16589 7701 16623 7735
rect 17601 7701 17635 7735
rect 18061 7701 18095 7735
rect 18613 7701 18647 7735
rect 19349 7701 19383 7735
rect 19809 7701 19843 7735
rect 20545 7701 20579 7735
rect 20913 7701 20947 7735
rect 21649 7701 21683 7735
rect 22661 7701 22695 7735
rect 23949 7701 23983 7735
rect 3249 7497 3283 7531
rect 4537 7497 4571 7531
rect 7297 7497 7331 7531
rect 7941 7497 7975 7531
rect 12817 7497 12851 7531
rect 12985 7497 13019 7531
rect 14657 7497 14691 7531
rect 15735 7497 15769 7531
rect 16865 7497 16899 7531
rect 18889 7497 18923 7531
rect 20913 7497 20947 7531
rect 21189 7497 21223 7531
rect 1777 7429 1811 7463
rect 4169 7429 4203 7463
rect 4369 7429 4403 7463
rect 6469 7429 6503 7463
rect 7465 7429 7499 7463
rect 7665 7429 7699 7463
rect 9505 7429 9539 7463
rect 13185 7429 13219 7463
rect 14289 7429 14323 7463
rect 14489 7429 14523 7463
rect 14933 7429 14967 7463
rect 15133 7429 15167 7463
rect 15945 7429 15979 7463
rect 17417 7429 17451 7463
rect 19441 7429 19475 7463
rect 21357 7429 21391 7463
rect 21557 7429 21591 7463
rect 22569 7429 22603 7463
rect 3800 7361 3834 7395
rect 3893 7361 3927 7395
rect 5181 7361 5215 7395
rect 5917 7361 5951 7395
rect 6101 7361 6135 7395
rect 6653 7361 6687 7395
rect 6745 7361 6779 7395
rect 8125 7361 8159 7395
rect 8585 7361 8619 7395
rect 13553 7361 13587 7395
rect 13645 7361 13679 7395
rect 13829 7361 13863 7395
rect 16221 7361 16255 7395
rect 16405 7361 16439 7395
rect 22293 7361 22327 7395
rect 1501 7293 1535 7327
rect 5641 7293 5675 7327
rect 8309 7293 8343 7327
rect 9229 7293 9263 7327
rect 11253 7293 11287 7327
rect 11621 7293 11655 7327
rect 11897 7293 11931 7327
rect 17141 7293 17175 7327
rect 19165 7293 19199 7327
rect 24041 7293 24075 7327
rect 3525 7225 3559 7259
rect 4353 7157 4387 7191
rect 4905 7157 4939 7191
rect 5365 7157 5399 7191
rect 5917 7157 5951 7191
rect 6469 7157 6503 7191
rect 7481 7157 7515 7191
rect 8677 7157 8711 7191
rect 13001 7157 13035 7191
rect 14473 7157 14507 7191
rect 15117 7157 15151 7191
rect 15301 7157 15335 7191
rect 15577 7157 15611 7191
rect 15761 7157 15795 7191
rect 16313 7157 16347 7191
rect 21373 7157 21407 7191
rect 21925 7157 21959 7191
rect 24409 7157 24443 7191
rect 1869 6953 1903 6987
rect 6193 6953 6227 6987
rect 7665 6953 7699 6987
rect 17969 6953 18003 6987
rect 18429 6953 18463 6987
rect 19625 6953 19659 6987
rect 20342 6953 20376 6987
rect 21833 6953 21867 6987
rect 2697 6885 2731 6919
rect 3433 6885 3467 6919
rect 6009 6885 6043 6919
rect 6561 6885 6595 6919
rect 12173 6885 12207 6919
rect 2329 6817 2363 6851
rect 4169 6817 4203 6851
rect 5733 6817 5767 6851
rect 6469 6817 6503 6851
rect 10333 6817 10367 6851
rect 13185 6817 13219 6851
rect 16221 6817 16255 6851
rect 22753 6817 22787 6851
rect 23765 6817 23799 6851
rect 3893 6749 3927 6783
rect 5181 6749 5215 6783
rect 5273 6749 5307 6783
rect 5365 6749 5399 6783
rect 7757 6749 7791 6783
rect 8217 6749 8251 6783
rect 8493 6749 8527 6783
rect 9045 6749 9079 6783
rect 9965 6749 9999 6783
rect 10241 6749 10275 6783
rect 10425 6749 10459 6783
rect 10977 6749 11011 6783
rect 11345 6749 11379 6783
rect 11989 6749 12023 6783
rect 12541 6749 12575 6783
rect 12909 6749 12943 6783
rect 14197 6749 14231 6783
rect 20085 6749 20119 6783
rect 23581 6749 23615 6783
rect 1685 6681 1719 6715
rect 1901 6681 1935 6715
rect 3065 6681 3099 6715
rect 6929 6681 6963 6715
rect 9505 6681 9539 6715
rect 14473 6681 14507 6715
rect 16497 6681 16531 6715
rect 18613 6681 18647 6715
rect 19717 6681 19751 6715
rect 22477 6681 22511 6715
rect 2053 6613 2087 6647
rect 2789 6613 2823 6647
rect 3525 6613 3559 6647
rect 4997 6613 5031 6647
rect 8309 6613 8343 6647
rect 8677 6613 8711 6647
rect 15945 6613 15979 6647
rect 18245 6613 18279 6647
rect 18403 6613 18437 6647
rect 18981 6613 19015 6647
rect 22109 6613 22143 6647
rect 22569 6613 22603 6647
rect 23121 6613 23155 6647
rect 23489 6613 23523 6647
rect 6837 6409 6871 6443
rect 7297 6409 7331 6443
rect 8309 6409 8343 6443
rect 8953 6409 8987 6443
rect 9689 6409 9723 6443
rect 14657 6409 14691 6443
rect 16773 6409 16807 6443
rect 17233 6409 17267 6443
rect 17877 6409 17911 6443
rect 19165 6409 19199 6443
rect 24041 6409 24075 6443
rect 7665 6341 7699 6375
rect 7849 6341 7883 6375
rect 15025 6341 15059 6375
rect 21189 6341 21223 6375
rect 21405 6341 21439 6375
rect 22293 6341 22327 6375
rect 24193 6341 24227 6375
rect 24409 6341 24443 6375
rect 1685 6273 1719 6307
rect 1961 6273 1995 6307
rect 2329 6273 2363 6307
rect 2605 6273 2639 6307
rect 2881 6273 2915 6307
rect 3709 6273 3743 6307
rect 3801 6273 3835 6307
rect 4721 6273 4755 6307
rect 4997 6273 5031 6307
rect 5549 6273 5583 6307
rect 6469 6273 6503 6307
rect 6562 6273 6596 6307
rect 7113 6273 7147 6307
rect 7297 6273 7331 6307
rect 7573 6273 7607 6307
rect 8585 6273 8619 6307
rect 9413 6273 9447 6307
rect 10455 6273 10489 6307
rect 10609 6273 10643 6307
rect 10977 6273 11011 6307
rect 11805 6273 11839 6307
rect 15117 6273 15151 6307
rect 15669 6273 15703 6307
rect 15853 6273 15887 6307
rect 16405 6273 16439 6307
rect 17141 6273 17175 6307
rect 17969 6273 18003 6307
rect 18337 6273 18371 6307
rect 18521 6273 18555 6307
rect 20729 6273 20763 6307
rect 1593 6205 1627 6239
rect 2421 6205 2455 6239
rect 8493 6205 8527 6239
rect 9321 6205 9355 6239
rect 9965 6205 9999 6239
rect 10241 6205 10275 6239
rect 12081 6205 12115 6239
rect 13553 6205 13587 6239
rect 13829 6205 13863 6239
rect 15301 6205 15335 6239
rect 17417 6205 17451 6239
rect 18889 6205 18923 6239
rect 19073 6205 19107 6239
rect 20177 6205 20211 6239
rect 22017 6205 22051 6239
rect 5457 6137 5491 6171
rect 15669 6137 15703 6171
rect 18337 6137 18371 6171
rect 3065 6069 3099 6103
rect 6101 6069 6135 6103
rect 7573 6069 7607 6103
rect 11069 6069 11103 6103
rect 14289 6069 14323 6103
rect 16221 6069 16255 6103
rect 19533 6069 19567 6103
rect 21373 6069 21407 6103
rect 21557 6069 21591 6103
rect 23765 6069 23799 6103
rect 24225 6069 24259 6103
rect 4077 5865 4111 5899
rect 8217 5865 8251 5899
rect 12265 5865 12299 5899
rect 16865 5865 16899 5899
rect 17785 5865 17819 5899
rect 19441 5865 19475 5899
rect 19901 5865 19935 5899
rect 21925 5865 21959 5899
rect 14197 5797 14231 5831
rect 2237 5729 2271 5763
rect 4261 5729 4295 5763
rect 6837 5729 6871 5763
rect 7297 5729 7331 5763
rect 7941 5729 7975 5763
rect 15761 5729 15795 5763
rect 21373 5729 21407 5763
rect 21649 5729 21683 5763
rect 22385 5729 22419 5763
rect 24133 5729 24167 5763
rect 1777 5661 1811 5695
rect 2145 5661 2179 5695
rect 2973 5661 3007 5695
rect 3157 5661 3191 5695
rect 3985 5661 4019 5695
rect 4813 5661 4847 5695
rect 4997 5661 5031 5695
rect 5457 5661 5491 5695
rect 5550 5661 5584 5695
rect 5733 5661 5767 5695
rect 5922 5661 5956 5695
rect 6377 5661 6411 5695
rect 6561 5661 6595 5695
rect 7021 5661 7055 5695
rect 7665 5661 7699 5695
rect 8401 5661 8435 5695
rect 8493 5661 8527 5695
rect 8585 5661 8619 5695
rect 9045 5661 9079 5695
rect 9229 5661 9263 5695
rect 9505 5661 9539 5695
rect 10701 5661 10735 5695
rect 10793 5661 10827 5695
rect 10885 5661 10919 5695
rect 11620 5661 11654 5695
rect 11713 5661 11747 5695
rect 12449 5661 12483 5695
rect 12541 5661 12575 5695
rect 12817 5661 12851 5695
rect 13185 5661 13219 5695
rect 13369 5661 13403 5695
rect 13553 5661 13587 5695
rect 15055 5661 15089 5695
rect 15209 5661 15243 5695
rect 15485 5661 15519 5695
rect 16405 5661 16439 5695
rect 18245 5661 18279 5695
rect 18981 5661 19015 5695
rect 19533 5661 19567 5695
rect 22109 5661 22143 5695
rect 5825 5593 5859 5627
rect 6469 5593 6503 5627
rect 7205 5593 7239 5627
rect 12909 5593 12943 5627
rect 14381 5593 14415 5627
rect 16681 5593 16715 5627
rect 16897 5593 16931 5627
rect 17601 5593 17635 5627
rect 22661 5593 22695 5627
rect 4813 5525 4847 5559
rect 6101 5525 6135 5559
rect 9229 5525 9263 5559
rect 10057 5525 10091 5559
rect 11069 5525 11103 5559
rect 11345 5525 11379 5559
rect 14841 5525 14875 5559
rect 17049 5525 17083 5559
rect 17801 5525 17835 5559
rect 17969 5525 18003 5559
rect 18429 5525 18463 5559
rect 18889 5525 18923 5559
rect 4169 5321 4203 5355
rect 7297 5321 7331 5355
rect 7389 5321 7423 5355
rect 8769 5321 8803 5355
rect 12357 5321 12391 5355
rect 15393 5321 15427 5355
rect 18705 5321 18739 5355
rect 20729 5321 20763 5355
rect 21005 5321 21039 5355
rect 21173 5321 21207 5355
rect 22845 5321 22879 5355
rect 23213 5321 23247 5355
rect 23305 5321 23339 5355
rect 24041 5321 24075 5355
rect 1685 5253 1719 5287
rect 14289 5253 14323 5287
rect 14473 5253 14507 5287
rect 14841 5253 14875 5287
rect 19257 5253 19291 5287
rect 21373 5253 21407 5287
rect 22201 5253 22235 5287
rect 22417 5253 22451 5287
rect 24193 5253 24227 5287
rect 24409 5253 24443 5287
rect 2605 5185 2639 5219
rect 3065 5185 3099 5219
rect 3617 5185 3651 5219
rect 4077 5185 4111 5219
rect 4353 5185 4387 5219
rect 5181 5185 5215 5219
rect 5733 5185 5767 5219
rect 7021 5185 7055 5219
rect 7113 5185 7147 5219
rect 7849 5185 7883 5219
rect 8217 5185 8251 5219
rect 8677 5185 8711 5219
rect 10241 5185 10275 5219
rect 10425 5185 10459 5219
rect 10701 5185 10735 5219
rect 10885 5185 10919 5219
rect 11988 5185 12022 5219
rect 12081 5185 12115 5219
rect 12541 5185 12575 5219
rect 13553 5185 13587 5219
rect 13737 5185 13771 5219
rect 13829 5185 13863 5219
rect 14565 5185 14599 5219
rect 15393 5185 15427 5219
rect 15853 5185 15887 5219
rect 15945 5185 15979 5219
rect 4813 5117 4847 5151
rect 5549 5117 5583 5151
rect 7481 5117 7515 5151
rect 9689 5117 9723 5151
rect 10609 5117 10643 5151
rect 12633 5117 12667 5151
rect 12725 5117 12759 5151
rect 12817 5117 12851 5151
rect 15485 5117 15519 5151
rect 16129 5117 16163 5151
rect 16957 5117 16991 5151
rect 17233 5117 17267 5151
rect 18981 5117 19015 5151
rect 23397 5117 23431 5151
rect 2053 5049 2087 5083
rect 6101 5049 6135 5083
rect 11713 5049 11747 5083
rect 13737 5049 13771 5083
rect 14381 5049 14415 5083
rect 2145 4981 2179 5015
rect 3525 4981 3559 5015
rect 4353 4981 4387 5015
rect 6469 4981 6503 5015
rect 6837 4981 6871 5015
rect 9229 4981 9263 5015
rect 16037 4981 16071 5015
rect 21189 4981 21223 5015
rect 22385 4981 22419 5015
rect 22569 4981 22603 5015
rect 24225 4981 24259 5015
rect 1501 4777 1535 4811
rect 2605 4777 2639 4811
rect 5181 4777 5215 4811
rect 9873 4777 9907 4811
rect 13093 4777 13127 4811
rect 15485 4777 15519 4811
rect 17325 4777 17359 4811
rect 19533 4777 19567 4811
rect 19717 4777 19751 4811
rect 22385 4777 22419 4811
rect 24133 4777 24167 4811
rect 1869 4709 1903 4743
rect 12633 4709 12667 4743
rect 15209 4709 15243 4743
rect 18429 4709 18463 4743
rect 2881 4641 2915 4675
rect 2973 4641 3007 4675
rect 3065 4641 3099 4675
rect 5365 4641 5399 4675
rect 6101 4641 6135 4675
rect 6193 4641 6227 4675
rect 6285 4641 6319 4675
rect 6929 4641 6963 4675
rect 7389 4641 7423 4675
rect 8401 4641 8435 4675
rect 14197 4641 14231 4675
rect 16773 4641 16807 4675
rect 17877 4641 17911 4675
rect 23213 4641 23247 4675
rect 2053 4573 2087 4607
rect 2329 4573 2363 4607
rect 2789 4573 2823 4607
rect 3893 4573 3927 4607
rect 4261 4573 4295 4607
rect 4629 4573 4663 4607
rect 5457 4573 5491 4607
rect 6377 4573 6411 4607
rect 7021 4573 7055 4607
rect 7297 4573 7331 4607
rect 8677 4573 8711 4607
rect 9045 4573 9079 4607
rect 9229 4573 9263 4607
rect 9781 4573 9815 4607
rect 9873 4573 9907 4607
rect 10241 4573 10275 4607
rect 10517 4573 10551 4607
rect 10793 4573 10827 4607
rect 10977 4573 11011 4607
rect 11437 4573 11471 4607
rect 11621 4573 11655 4607
rect 11713 4573 11747 4607
rect 12541 4573 12575 4607
rect 12725 4573 12759 4607
rect 13272 4573 13306 4607
rect 13369 4573 13403 4607
rect 13461 4573 13495 4607
rect 13589 4573 13623 4607
rect 13737 4573 13771 4607
rect 14381 4573 14415 4607
rect 14565 4573 14599 4607
rect 14657 4573 14691 4607
rect 14933 4573 14967 4607
rect 15485 4573 15519 4607
rect 15761 4573 15795 4607
rect 17693 4573 17727 4607
rect 18889 4573 18923 4607
rect 19993 4573 20027 4607
rect 9597 4505 9631 4539
rect 10885 4505 10919 4539
rect 15209 4505 15243 4539
rect 17785 4505 17819 4539
rect 19349 4505 19383 4539
rect 19565 4505 19599 4539
rect 20269 4505 20303 4539
rect 22109 4505 22143 4539
rect 2237 4437 2271 4471
rect 3433 4437 3467 4471
rect 5917 4437 5951 4471
rect 6745 4437 6779 4471
rect 9229 4437 9263 4471
rect 11253 4437 11287 4471
rect 11989 4437 12023 4471
rect 15025 4437 15059 4471
rect 15669 4437 15703 4471
rect 16313 4437 16347 4471
rect 21741 4437 21775 4471
rect 23305 4437 23339 4471
rect 23397 4437 23431 4471
rect 23765 4437 23799 4471
rect 4169 4233 4203 4267
rect 12541 4233 12575 4267
rect 16129 4233 16163 4267
rect 19231 4233 19265 4267
rect 19917 4233 19951 4267
rect 20361 4233 20395 4267
rect 20821 4233 20855 4267
rect 21557 4233 21591 4267
rect 1961 4165 1995 4199
rect 5641 4165 5675 4199
rect 6929 4165 6963 4199
rect 18797 4165 18831 4199
rect 19441 4165 19475 4199
rect 19717 4165 19751 4199
rect 20729 4165 20763 4199
rect 3985 4097 4019 4131
rect 4445 4097 4479 4131
rect 4629 4097 4663 4131
rect 5273 4097 5307 4131
rect 5365 4097 5399 4131
rect 9229 4097 9263 4131
rect 9413 4097 9447 4131
rect 9873 4097 9907 4131
rect 9965 4097 9999 4131
rect 10057 4097 10091 4131
rect 10241 4097 10275 4131
rect 10701 4097 10735 4131
rect 10977 4097 11011 4131
rect 11621 4097 11655 4131
rect 11805 4097 11839 4131
rect 13185 4097 13219 4131
rect 13369 4097 13403 4131
rect 13829 4097 13863 4131
rect 14473 4097 14507 4131
rect 14565 4097 14599 4131
rect 15669 4097 15703 4131
rect 16313 4097 16347 4131
rect 16405 4097 16439 4131
rect 21373 4097 21407 4131
rect 24409 4097 24443 4131
rect 1685 4029 1719 4063
rect 3709 4029 3743 4063
rect 4813 4029 4847 4063
rect 5733 4029 5767 4063
rect 6653 4029 6687 4063
rect 10517 4029 10551 4063
rect 10885 4029 10919 4063
rect 12081 4029 12115 4063
rect 15301 4029 15335 4063
rect 15577 4029 15611 4063
rect 16129 4029 16163 4063
rect 16773 4029 16807 4063
rect 17049 4029 17083 4063
rect 21005 4029 21039 4063
rect 22201 4029 22235 4063
rect 22477 4029 22511 4063
rect 23949 4029 23983 4063
rect 3801 3961 3835 3995
rect 9321 3961 9355 3995
rect 12449 3961 12483 3995
rect 24225 3961 24259 3995
rect 3433 3893 3467 3927
rect 5089 3893 5123 3927
rect 6101 3893 6135 3927
rect 8401 3893 8435 3927
rect 9689 3893 9723 3927
rect 11713 3893 11747 3927
rect 12909 3893 12943 3927
rect 13553 3893 13587 3927
rect 13921 3893 13955 3927
rect 19073 3893 19107 3927
rect 19257 3893 19291 3927
rect 19901 3893 19935 3927
rect 20085 3893 20119 3927
rect 2145 3689 2179 3723
rect 2329 3689 2363 3723
rect 7205 3689 7239 3723
rect 7389 3689 7423 3723
rect 10793 3689 10827 3723
rect 15402 3689 15436 3723
rect 16405 3689 16439 3723
rect 19809 3689 19843 3723
rect 20177 3689 20211 3723
rect 22569 3689 22603 3723
rect 23949 3689 23983 3723
rect 1685 3621 1719 3655
rect 2605 3621 2639 3655
rect 11161 3621 11195 3655
rect 23765 3621 23799 3655
rect 2789 3553 2823 3587
rect 2881 3553 2915 3587
rect 3157 3553 3191 3587
rect 4905 3553 4939 3587
rect 7849 3553 7883 3587
rect 9321 3553 9355 3587
rect 13553 3553 13587 3587
rect 13829 3553 13863 3587
rect 18981 3553 19015 3587
rect 21189 3553 21223 3587
rect 23029 3553 23063 3587
rect 23121 3553 23155 3587
rect 1501 3485 1535 3519
rect 2697 3485 2731 3519
rect 2973 3485 3007 3519
rect 3525 3485 3559 3519
rect 4629 3485 4663 3519
rect 7721 3485 7755 3519
rect 7941 3485 7975 3519
rect 8125 3485 8159 3519
rect 8401 3485 8435 3519
rect 9045 3485 9079 3519
rect 11805 3485 11839 3519
rect 12081 3485 12115 3519
rect 14289 3485 14323 3519
rect 14565 3485 14599 3519
rect 14749 3485 14783 3519
rect 15853 3485 15887 3519
rect 16129 3485 16163 3519
rect 16221 3485 16255 3519
rect 16681 3485 16715 3519
rect 19349 3485 19383 3519
rect 20361 3485 20395 3519
rect 22201 3485 22235 3519
rect 22937 3485 22971 3519
rect 1961 3417 1995 3451
rect 4077 3417 4111 3451
rect 5181 3417 5215 3451
rect 7021 3417 7055 3451
rect 7849 3417 7883 3451
rect 11437 3417 11471 3451
rect 15577 3417 15611 3451
rect 16037 3417 16071 3451
rect 18705 3417 18739 3451
rect 21925 3417 21959 3451
rect 24133 3417 24167 3451
rect 2161 3349 2195 3383
rect 3985 3349 4019 3383
rect 4445 3349 4479 3383
rect 6653 3349 6687 3383
rect 7221 3349 7255 3383
rect 8585 3349 8619 3383
rect 15209 3349 15243 3383
rect 15377 3349 15411 3383
rect 16865 3349 16899 3383
rect 17233 3349 17267 3383
rect 20637 3349 20671 3383
rect 21005 3349 21039 3383
rect 21097 3349 21131 3383
rect 23933 3349 23967 3383
rect 3709 3145 3743 3179
rect 5841 3145 5875 3179
rect 6009 3145 6043 3179
rect 8309 3145 8343 3179
rect 12817 3145 12851 3179
rect 16037 3145 16071 3179
rect 17801 3145 17835 3179
rect 17969 3145 18003 3179
rect 18245 3145 18279 3179
rect 19441 3145 19475 3179
rect 21557 3145 21591 3179
rect 21925 3145 21959 3179
rect 22569 3145 22603 3179
rect 4169 3077 4203 3111
rect 5641 3077 5675 3111
rect 11989 3077 12023 3111
rect 14749 3077 14783 3111
rect 17601 3077 17635 3111
rect 18613 3077 18647 3111
rect 22093 3077 22127 3111
rect 22293 3077 22327 3111
rect 1777 3009 1811 3043
rect 2237 3009 2271 3043
rect 2973 3009 3007 3043
rect 3617 3009 3651 3043
rect 3801 3009 3835 3043
rect 4077 3009 4111 3043
rect 4261 3009 4295 3043
rect 4537 3009 4571 3043
rect 4721 3009 4755 3043
rect 4997 3009 5031 3043
rect 5090 3009 5124 3043
rect 6745 3009 6779 3043
rect 7297 3009 7331 3043
rect 7849 3009 7883 3043
rect 8125 3009 8159 3043
rect 9781 3009 9815 3043
rect 10425 3009 10459 3043
rect 10885 3009 10919 3043
rect 11621 3009 11655 3043
rect 11805 3009 11839 3043
rect 12817 3009 12851 3043
rect 13553 3009 13587 3043
rect 14013 3009 14047 3043
rect 14197 3009 14231 3043
rect 14657 3009 14691 3043
rect 15025 3009 15059 3043
rect 15209 3009 15243 3043
rect 15577 3009 15611 3043
rect 15853 3009 15887 3043
rect 18705 3009 18739 3043
rect 19257 3009 19291 3043
rect 19809 3009 19843 3043
rect 24317 3009 24351 3043
rect 2697 2941 2731 2975
rect 2881 2941 2915 2975
rect 6561 2941 6595 2975
rect 9229 2941 9263 2975
rect 10793 2941 10827 2975
rect 12265 2941 12299 2975
rect 12909 2941 12943 2975
rect 13277 2941 13311 2975
rect 16773 2941 16807 2975
rect 18889 2941 18923 2975
rect 20085 2941 20119 2975
rect 24041 2941 24075 2975
rect 2421 2873 2455 2907
rect 5365 2873 5399 2907
rect 7481 2873 7515 2907
rect 8769 2873 8803 2907
rect 11253 2873 11287 2907
rect 15669 2873 15703 2907
rect 16405 2873 16439 2907
rect 1869 2805 1903 2839
rect 2789 2805 2823 2839
rect 4629 2805 4663 2839
rect 5825 2805 5859 2839
rect 9965 2805 9999 2839
rect 17233 2805 17267 2839
rect 17785 2805 17819 2839
rect 22149 2805 22183 2839
rect 1869 2601 1903 2635
rect 11437 2601 11471 2635
rect 17693 2601 17727 2635
rect 18153 2601 18187 2635
rect 18521 2601 18555 2635
rect 3433 2533 3467 2567
rect 9597 2533 9631 2567
rect 13553 2533 13587 2567
rect 18705 2533 18739 2567
rect 22385 2533 22419 2567
rect 2421 2465 2455 2499
rect 2697 2465 2731 2499
rect 6745 2465 6779 2499
rect 7849 2465 7883 2499
rect 8217 2465 8251 2499
rect 11253 2465 11287 2499
rect 14197 2465 14231 2499
rect 14749 2465 14783 2499
rect 15577 2465 15611 2499
rect 15853 2465 15887 2499
rect 16129 2465 16163 2499
rect 16589 2465 16623 2499
rect 16681 2465 16715 2499
rect 16773 2465 16807 2499
rect 16957 2465 16991 2499
rect 17233 2465 17267 2499
rect 19533 2465 19567 2499
rect 19717 2465 19751 2499
rect 23673 2465 23707 2499
rect 1685 2397 1719 2431
rect 2329 2397 2363 2431
rect 2973 2397 3007 2431
rect 3157 2397 3191 2431
rect 3525 2397 3559 2431
rect 3985 2397 4019 2431
rect 4537 2397 4571 2431
rect 4721 2397 4755 2431
rect 5549 2397 5583 2431
rect 5825 2397 5859 2431
rect 6285 2397 6319 2431
rect 6837 2397 6871 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 7941 2397 7975 2431
rect 8389 2391 8423 2425
rect 8493 2407 8527 2441
rect 8585 2397 8619 2431
rect 9045 2397 9079 2431
rect 10057 2397 10091 2431
rect 10609 2397 10643 2431
rect 11161 2397 11195 2431
rect 11989 2397 12023 2431
rect 12357 2397 12391 2431
rect 12449 2397 12483 2431
rect 13185 2397 13219 2431
rect 13369 2397 13403 2431
rect 15025 2397 15059 2431
rect 15761 2397 15795 2431
rect 16037 2397 16071 2431
rect 16497 2397 16531 2431
rect 18061 2397 18095 2431
rect 18245 2397 18279 2431
rect 20637 2397 20671 2431
rect 21649 2397 21683 2431
rect 22293 2397 22327 2431
rect 23489 2397 23523 2431
rect 5089 2329 5123 2363
rect 15945 2329 15979 2363
rect 18981 2329 19015 2363
rect 19809 2329 19843 2363
rect 9229 2261 9263 2295
rect 20177 2261 20211 2295
rect 1501 2057 1535 2091
rect 3985 2057 4019 2091
rect 4261 2057 4295 2091
rect 5197 2057 5231 2091
rect 5365 2057 5399 2091
rect 11161 2057 11195 2091
rect 14841 2057 14875 2091
rect 18889 2057 18923 2091
rect 21389 2057 21423 2091
rect 21557 2057 21591 2091
rect 24041 2057 24075 2091
rect 2973 1989 3007 2023
rect 4997 1989 5031 2023
rect 6561 1989 6595 2023
rect 6745 1989 6779 2023
rect 8033 1989 8067 2023
rect 12173 1989 12207 2023
rect 14993 1989 15027 2023
rect 15209 1989 15243 2023
rect 16037 1989 16071 2023
rect 17049 1989 17083 2023
rect 21189 1989 21223 2023
rect 23489 1989 23523 2023
rect 24204 1989 24238 2023
rect 24409 1989 24443 2023
rect 3249 1921 3283 1955
rect 3801 1921 3835 1955
rect 4721 1921 4755 1955
rect 6469 1921 6503 1955
rect 7389 1921 7423 1955
rect 9781 1921 9815 1955
rect 10057 1921 10091 1955
rect 10211 1921 10245 1955
rect 11989 1921 12023 1955
rect 12357 1921 12391 1955
rect 12725 1921 12759 1955
rect 13553 1921 13587 1955
rect 13645 1921 13679 1955
rect 14197 1921 14231 1955
rect 14565 1921 14599 1955
rect 16313 1921 16347 1955
rect 16773 1921 16807 1955
rect 23765 1921 23799 1955
rect 3525 1853 3559 1887
rect 5641 1853 5675 1887
rect 7757 1853 7791 1887
rect 10701 1853 10735 1887
rect 12817 1853 12851 1887
rect 20361 1853 20395 1887
rect 20637 1853 20671 1887
rect 4353 1785 4387 1819
rect 6009 1785 6043 1819
rect 6745 1785 6779 1819
rect 18521 1785 18555 1819
rect 3617 1717 3651 1751
rect 5181 1717 5215 1751
rect 6101 1717 6135 1751
rect 7297 1717 7331 1751
rect 10241 1717 10275 1751
rect 15025 1717 15059 1751
rect 21373 1717 21407 1751
rect 22017 1717 22051 1751
rect 24225 1717 24259 1751
rect 1961 1513 1995 1547
rect 2145 1513 2179 1547
rect 6101 1513 6135 1547
rect 10793 1513 10827 1547
rect 17049 1513 17083 1547
rect 17233 1513 17267 1547
rect 17509 1513 17543 1547
rect 18153 1513 18187 1547
rect 18797 1513 18831 1547
rect 20072 1513 20106 1547
rect 21557 1513 21591 1547
rect 21925 1513 21959 1547
rect 23869 1513 23903 1547
rect 3065 1445 3099 1479
rect 11805 1445 11839 1479
rect 12173 1445 12207 1479
rect 19441 1445 19475 1479
rect 4997 1377 5031 1411
rect 7113 1377 7147 1411
rect 13185 1377 13219 1411
rect 14473 1377 14507 1411
rect 19809 1377 19843 1411
rect 24133 1377 24167 1411
rect 1501 1309 1535 1343
rect 2789 1309 2823 1343
rect 3279 1309 3313 1343
rect 3433 1309 3467 1343
rect 4123 1309 4157 1343
rect 4261 1309 4295 1343
rect 4537 1309 4571 1343
rect 5181 1309 5215 1343
rect 5365 1309 5399 1343
rect 5641 1309 5675 1343
rect 5733 1309 5767 1343
rect 5917 1309 5951 1343
rect 6469 1309 6503 1343
rect 6929 1309 6963 1343
rect 7849 1309 7883 1343
rect 9413 1309 9447 1343
rect 9965 1309 9999 1343
rect 10425 1309 10459 1343
rect 11069 1309 11103 1343
rect 11621 1309 11655 1343
rect 12081 1309 12115 1343
rect 12541 1309 12575 1343
rect 12909 1309 12943 1343
rect 13553 1309 13587 1343
rect 14197 1309 14231 1343
rect 15761 1309 15795 1343
rect 16037 1309 16071 1343
rect 17509 1309 17543 1343
rect 17705 1309 17739 1343
rect 18827 1309 18861 1343
rect 18981 1309 19015 1343
rect 19349 1309 19383 1343
rect 19533 1309 19567 1343
rect 21925 1309 21959 1343
rect 22109 1309 22143 1343
rect 2129 1241 2163 1275
rect 2329 1241 2363 1275
rect 3893 1241 3927 1275
rect 8585 1241 8619 1275
rect 16865 1241 16899 1275
rect 17065 1241 17099 1275
rect 17969 1241 18003 1275
rect 18185 1241 18219 1275
rect 1685 1173 1719 1207
rect 2697 1173 2731 1207
rect 4721 1173 4755 1207
rect 6653 1173 6687 1207
rect 8493 1173 8527 1207
rect 9137 1173 9171 1207
rect 18337 1173 18371 1207
rect 22385 1173 22419 1207
<< metal1 >>
rect 13814 19252 13820 19304
rect 13872 19292 13878 19304
rect 24394 19292 24400 19304
rect 13872 19264 24400 19292
rect 13872 19252 13878 19264
rect 24394 19252 24400 19264
rect 24452 19252 24458 19304
rect 13354 18640 13360 18692
rect 13412 18680 13418 18692
rect 21450 18680 21456 18692
rect 13412 18652 21456 18680
rect 13412 18640 13418 18652
rect 21450 18640 21456 18652
rect 21508 18640 21514 18692
rect 13170 18572 13176 18624
rect 13228 18612 13234 18624
rect 23474 18612 23480 18624
rect 13228 18584 23480 18612
rect 13228 18572 13234 18584
rect 23474 18572 23480 18584
rect 23532 18572 23538 18624
rect 1104 18522 24840 18544
rect 1104 18470 8214 18522
rect 8266 18470 8278 18522
rect 8330 18470 8342 18522
rect 8394 18470 8406 18522
rect 8458 18470 8470 18522
rect 8522 18470 16214 18522
rect 16266 18470 16278 18522
rect 16330 18470 16342 18522
rect 16394 18470 16406 18522
rect 16458 18470 16470 18522
rect 16522 18470 24214 18522
rect 24266 18470 24278 18522
rect 24330 18470 24342 18522
rect 24394 18470 24406 18522
rect 24458 18470 24470 18522
rect 24522 18470 24840 18522
rect 1104 18448 24840 18470
rect 3145 18411 3203 18417
rect 3145 18377 3157 18411
rect 3191 18408 3203 18411
rect 10870 18408 10876 18420
rect 3191 18380 10876 18408
rect 3191 18377 3203 18380
rect 3145 18371 3203 18377
rect 10870 18368 10876 18380
rect 10928 18368 10934 18420
rect 13354 18368 13360 18420
rect 13412 18368 13418 18420
rect 14182 18368 14188 18420
rect 14240 18408 14246 18420
rect 20622 18408 20628 18420
rect 14240 18380 20628 18408
rect 14240 18368 14246 18380
rect 20622 18368 20628 18380
rect 20680 18368 20686 18420
rect 20898 18368 20904 18420
rect 20956 18408 20962 18420
rect 22741 18411 22799 18417
rect 22741 18408 22753 18411
rect 20956 18380 22753 18408
rect 20956 18368 20962 18380
rect 22741 18377 22753 18380
rect 22787 18377 22799 18411
rect 22741 18371 22799 18377
rect 1854 18300 1860 18352
rect 1912 18340 1918 18352
rect 2317 18343 2375 18349
rect 2317 18340 2329 18343
rect 1912 18312 2329 18340
rect 1912 18300 1918 18312
rect 2317 18309 2329 18312
rect 2363 18309 2375 18343
rect 2317 18303 2375 18309
rect 2406 18300 2412 18352
rect 2464 18340 2470 18352
rect 2517 18343 2575 18349
rect 2517 18340 2529 18343
rect 2464 18312 2529 18340
rect 2464 18300 2470 18312
rect 2517 18309 2529 18312
rect 2563 18309 2575 18343
rect 2517 18303 2575 18309
rect 8281 18343 8339 18349
rect 8281 18309 8293 18343
rect 8327 18340 8339 18343
rect 8481 18343 8539 18349
rect 8327 18309 8340 18340
rect 8281 18303 8340 18309
rect 8481 18309 8493 18343
rect 8527 18340 8539 18343
rect 9674 18340 9680 18352
rect 8527 18312 9680 18340
rect 8527 18309 8539 18312
rect 8481 18303 8539 18309
rect 1302 18232 1308 18284
rect 1360 18272 1366 18284
rect 1489 18275 1547 18281
rect 1489 18272 1501 18275
rect 1360 18244 1501 18272
rect 1360 18232 1366 18244
rect 1489 18241 1501 18244
rect 1535 18272 1547 18275
rect 1949 18275 2007 18281
rect 1949 18272 1961 18275
rect 1535 18244 1961 18272
rect 1535 18241 1547 18244
rect 1489 18235 1547 18241
rect 1949 18241 1961 18244
rect 1995 18241 2007 18275
rect 1949 18235 2007 18241
rect 2958 18232 2964 18284
rect 3016 18272 3022 18284
rect 3421 18275 3479 18281
rect 3421 18272 3433 18275
rect 3016 18244 3433 18272
rect 3016 18232 3022 18244
rect 3421 18241 3433 18244
rect 3467 18241 3479 18275
rect 3421 18235 3479 18241
rect 3878 18232 3884 18284
rect 3936 18272 3942 18284
rect 3973 18275 4031 18281
rect 3973 18272 3985 18275
rect 3936 18244 3985 18272
rect 3936 18232 3942 18244
rect 3973 18241 3985 18244
rect 4019 18272 4031 18275
rect 4433 18275 4491 18281
rect 4433 18272 4445 18275
rect 4019 18244 4445 18272
rect 4019 18241 4031 18244
rect 3973 18235 4031 18241
rect 4433 18241 4445 18244
rect 4479 18241 4491 18275
rect 4433 18235 4491 18241
rect 5258 18232 5264 18284
rect 5316 18232 5322 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 6549 18275 6607 18281
rect 6549 18272 6561 18275
rect 6512 18244 6561 18272
rect 6512 18232 6518 18244
rect 6549 18241 6561 18244
rect 6595 18272 6607 18275
rect 7009 18275 7067 18281
rect 7009 18272 7021 18275
rect 6595 18244 7021 18272
rect 6595 18241 6607 18244
rect 6549 18235 6607 18241
rect 7009 18241 7021 18244
rect 7055 18241 7067 18275
rect 8312 18272 8340 18303
rect 9674 18300 9680 18312
rect 9732 18300 9738 18352
rect 10781 18343 10839 18349
rect 10781 18309 10793 18343
rect 10827 18340 10839 18343
rect 16117 18343 16175 18349
rect 10827 18312 13216 18340
rect 10827 18309 10839 18312
rect 10781 18303 10839 18309
rect 13188 18284 13216 18312
rect 16117 18309 16129 18343
rect 16163 18340 16175 18343
rect 16942 18340 16948 18352
rect 16163 18312 16948 18340
rect 16163 18309 16175 18312
rect 16117 18303 16175 18309
rect 16942 18300 16948 18312
rect 17000 18300 17006 18352
rect 17494 18300 17500 18352
rect 17552 18340 17558 18352
rect 17552 18312 18920 18340
rect 17552 18300 17558 18312
rect 8846 18272 8852 18284
rect 8312 18244 8852 18272
rect 7009 18235 7067 18241
rect 8846 18232 8852 18244
rect 8904 18232 8910 18284
rect 9030 18232 9036 18284
rect 9088 18272 9094 18284
rect 9125 18275 9183 18281
rect 9125 18272 9137 18275
rect 9088 18244 9137 18272
rect 9088 18232 9094 18244
rect 9125 18241 9137 18244
rect 9171 18272 9183 18275
rect 9585 18275 9643 18281
rect 9585 18272 9597 18275
rect 9171 18244 9597 18272
rect 9171 18241 9183 18244
rect 9125 18235 9183 18241
rect 9585 18241 9597 18244
rect 9631 18241 9643 18275
rect 9585 18235 9643 18241
rect 11241 18275 11299 18281
rect 11241 18241 11253 18275
rect 11287 18272 11299 18275
rect 12621 18275 12679 18281
rect 11287 18244 12112 18272
rect 11287 18241 11299 18244
rect 11241 18235 11299 18241
rect 5350 18164 5356 18216
rect 5408 18164 5414 18216
rect 5442 18164 5448 18216
rect 5500 18164 5506 18216
rect 11514 18164 11520 18216
rect 11572 18204 11578 18216
rect 11609 18207 11667 18213
rect 11609 18204 11621 18207
rect 11572 18176 11621 18204
rect 11572 18164 11578 18176
rect 11609 18173 11621 18176
rect 11655 18173 11667 18207
rect 11609 18167 11667 18173
rect 12084 18148 12112 18244
rect 12621 18241 12633 18275
rect 12667 18272 12679 18275
rect 12710 18272 12716 18284
rect 12667 18244 12716 18272
rect 12667 18241 12679 18244
rect 12621 18235 12679 18241
rect 12710 18232 12716 18244
rect 12768 18232 12774 18284
rect 13170 18232 13176 18284
rect 13228 18232 13234 18284
rect 13633 18275 13691 18281
rect 13633 18241 13645 18275
rect 13679 18272 13691 18275
rect 13814 18272 13820 18284
rect 13679 18244 13820 18272
rect 13679 18241 13691 18244
rect 13633 18235 13691 18241
rect 13814 18232 13820 18244
rect 13872 18232 13878 18284
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14461 18235 14519 18241
rect 15381 18275 15439 18281
rect 15381 18241 15393 18275
rect 15427 18272 15439 18275
rect 16761 18275 16819 18281
rect 16761 18272 16773 18275
rect 15427 18244 16773 18272
rect 15427 18241 15439 18244
rect 15381 18235 15439 18241
rect 16761 18241 16773 18244
rect 16807 18241 16819 18275
rect 16761 18235 16819 18241
rect 12161 18207 12219 18213
rect 12161 18173 12173 18207
rect 12207 18173 12219 18207
rect 12161 18167 12219 18173
rect 4157 18139 4215 18145
rect 4157 18105 4169 18139
rect 4203 18136 4215 18139
rect 5166 18136 5172 18148
rect 4203 18108 5172 18136
rect 4203 18105 4215 18108
rect 4157 18099 4215 18105
rect 5166 18096 5172 18108
rect 5224 18096 5230 18148
rect 6733 18139 6791 18145
rect 6733 18105 6745 18139
rect 6779 18136 6791 18139
rect 6779 18108 11284 18136
rect 6779 18105 6791 18108
rect 6733 18099 6791 18105
rect 1670 18028 1676 18080
rect 1728 18028 1734 18080
rect 2498 18028 2504 18080
rect 2556 18028 2562 18080
rect 2590 18028 2596 18080
rect 2648 18068 2654 18080
rect 2685 18071 2743 18077
rect 2685 18068 2697 18071
rect 2648 18040 2697 18068
rect 2648 18028 2654 18040
rect 2685 18037 2697 18040
rect 2731 18037 2743 18071
rect 2685 18031 2743 18037
rect 4614 18028 4620 18080
rect 4672 18068 4678 18080
rect 4893 18071 4951 18077
rect 4893 18068 4905 18071
rect 4672 18040 4905 18068
rect 4672 18028 4678 18040
rect 4893 18037 4905 18040
rect 4939 18037 4951 18071
rect 4893 18031 4951 18037
rect 7926 18028 7932 18080
rect 7984 18068 7990 18080
rect 8113 18071 8171 18077
rect 8113 18068 8125 18071
rect 7984 18040 8125 18068
rect 7984 18028 7990 18040
rect 8113 18037 8125 18040
rect 8159 18037 8171 18071
rect 8113 18031 8171 18037
rect 8297 18071 8355 18077
rect 8297 18037 8309 18071
rect 8343 18068 8355 18071
rect 8570 18068 8576 18080
rect 8343 18040 8576 18068
rect 8343 18037 8355 18040
rect 8297 18031 8355 18037
rect 8570 18028 8576 18040
rect 8628 18028 8634 18080
rect 9306 18028 9312 18080
rect 9364 18028 9370 18080
rect 11146 18028 11152 18080
rect 11204 18028 11210 18080
rect 11256 18068 11284 18108
rect 12066 18096 12072 18148
rect 12124 18096 12130 18148
rect 12176 18136 12204 18167
rect 12437 18139 12495 18145
rect 12437 18136 12449 18139
rect 12176 18108 12449 18136
rect 12437 18105 12449 18108
rect 12483 18105 12495 18139
rect 13906 18136 13912 18148
rect 12437 18099 12495 18105
rect 13188 18108 13912 18136
rect 13188 18068 13216 18108
rect 13906 18096 13912 18108
rect 13964 18096 13970 18148
rect 14274 18096 14280 18148
rect 14332 18096 14338 18148
rect 14476 18136 14504 18235
rect 17402 18232 17408 18284
rect 17460 18232 17466 18284
rect 18690 18232 18696 18284
rect 18748 18272 18754 18284
rect 18785 18275 18843 18281
rect 18785 18272 18797 18275
rect 18748 18244 18797 18272
rect 18748 18232 18754 18244
rect 18785 18241 18797 18244
rect 18831 18241 18843 18275
rect 18892 18272 18920 18312
rect 19334 18300 19340 18352
rect 19392 18340 19398 18352
rect 21361 18343 21419 18349
rect 21361 18340 21373 18343
rect 19392 18312 20024 18340
rect 19392 18300 19398 18312
rect 19996 18281 20024 18312
rect 20548 18312 21373 18340
rect 20548 18281 20576 18312
rect 21361 18309 21373 18312
rect 21407 18340 21419 18343
rect 23658 18340 23664 18352
rect 21407 18312 23664 18340
rect 21407 18309 21419 18312
rect 21361 18303 21419 18309
rect 23658 18300 23664 18312
rect 23716 18300 23722 18352
rect 19521 18275 19579 18281
rect 19521 18272 19533 18275
rect 18892 18244 19533 18272
rect 18785 18235 18843 18241
rect 19521 18241 19533 18244
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19981 18275 20039 18281
rect 19981 18241 19993 18275
rect 20027 18241 20039 18275
rect 19981 18235 20039 18241
rect 20533 18275 20591 18281
rect 20533 18241 20545 18275
rect 20579 18241 20591 18275
rect 20533 18235 20591 18241
rect 20806 18232 20812 18284
rect 20864 18272 20870 18284
rect 21177 18275 21235 18281
rect 21177 18272 21189 18275
rect 20864 18244 21189 18272
rect 20864 18232 20870 18244
rect 21177 18241 21189 18244
rect 21223 18272 21235 18275
rect 21223 18244 21496 18272
rect 21223 18241 21235 18244
rect 21177 18235 21235 18241
rect 14550 18164 14556 18216
rect 14608 18204 14614 18216
rect 14829 18207 14887 18213
rect 14829 18204 14841 18207
rect 14608 18176 14841 18204
rect 14608 18164 14614 18176
rect 14829 18173 14841 18176
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 15657 18207 15715 18213
rect 15657 18173 15669 18207
rect 15703 18204 15715 18207
rect 16114 18204 16120 18216
rect 15703 18176 16120 18204
rect 15703 18173 15715 18176
rect 15657 18167 15715 18173
rect 16114 18164 16120 18176
rect 16172 18164 16178 18216
rect 16209 18207 16267 18213
rect 16209 18173 16221 18207
rect 16255 18173 16267 18207
rect 16209 18167 16267 18173
rect 15286 18136 15292 18148
rect 14476 18108 15292 18136
rect 15286 18096 15292 18108
rect 15344 18096 15350 18148
rect 16224 18136 16252 18167
rect 17862 18164 17868 18216
rect 17920 18164 17926 18216
rect 18414 18164 18420 18216
rect 18472 18164 18478 18216
rect 20898 18164 20904 18216
rect 20956 18164 20962 18216
rect 21468 18204 21496 18244
rect 23474 18232 23480 18284
rect 23532 18232 23538 18284
rect 24118 18232 24124 18284
rect 24176 18232 24182 18284
rect 21913 18207 21971 18213
rect 21913 18204 21925 18207
rect 21468 18176 21925 18204
rect 21913 18173 21925 18176
rect 21959 18173 21971 18207
rect 21913 18167 21971 18173
rect 22462 18164 22468 18216
rect 22520 18164 22526 18216
rect 17221 18139 17279 18145
rect 17221 18136 17233 18139
rect 16224 18108 17233 18136
rect 17221 18105 17233 18108
rect 17267 18105 17279 18139
rect 17221 18099 17279 18105
rect 17957 18139 18015 18145
rect 17957 18105 17969 18139
rect 18003 18136 18015 18139
rect 18322 18136 18328 18148
rect 18003 18108 18328 18136
rect 18003 18105 18015 18108
rect 17957 18099 18015 18105
rect 18322 18096 18328 18108
rect 18380 18096 18386 18148
rect 19978 18136 19984 18148
rect 18708 18108 19984 18136
rect 11256 18040 13216 18068
rect 13817 18071 13875 18077
rect 13817 18037 13829 18071
rect 13863 18068 13875 18071
rect 18708 18068 18736 18108
rect 19978 18096 19984 18108
rect 20036 18096 20042 18148
rect 21545 18139 21603 18145
rect 21545 18105 21557 18139
rect 21591 18136 21603 18139
rect 21818 18136 21824 18148
rect 21591 18108 21824 18136
rect 21591 18105 21603 18108
rect 21545 18099 21603 18105
rect 21818 18096 21824 18108
rect 21876 18096 21882 18148
rect 22373 18139 22431 18145
rect 22373 18105 22385 18139
rect 22419 18105 22431 18139
rect 22373 18099 22431 18105
rect 13863 18040 18736 18068
rect 13863 18037 13875 18040
rect 13817 18031 13875 18037
rect 18782 18028 18788 18080
rect 18840 18028 18846 18080
rect 19337 18071 19395 18077
rect 19337 18037 19349 18071
rect 19383 18068 19395 18071
rect 19426 18068 19432 18080
rect 19383 18040 19432 18068
rect 19383 18037 19395 18040
rect 19337 18031 19395 18037
rect 19426 18028 19432 18040
rect 19484 18028 19490 18080
rect 19794 18028 19800 18080
rect 19852 18028 19858 18080
rect 20901 18071 20959 18077
rect 20901 18037 20913 18071
rect 20947 18068 20959 18071
rect 21634 18068 21640 18080
rect 20947 18040 21640 18068
rect 20947 18037 20959 18040
rect 20901 18031 20959 18037
rect 21634 18028 21640 18040
rect 21692 18068 21698 18080
rect 22388 18068 22416 18099
rect 23198 18068 23204 18080
rect 21692 18040 23204 18068
rect 21692 18028 21698 18040
rect 23198 18028 23204 18040
rect 23256 18028 23262 18080
rect 23382 18028 23388 18080
rect 23440 18028 23446 18080
rect 23750 18028 23756 18080
rect 23808 18068 23814 18080
rect 23937 18071 23995 18077
rect 23937 18068 23949 18071
rect 23808 18040 23949 18068
rect 23808 18028 23814 18040
rect 23937 18037 23949 18040
rect 23983 18037 23995 18071
rect 23937 18031 23995 18037
rect 1104 17978 24840 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 12214 17978
rect 12266 17926 12278 17978
rect 12330 17926 12342 17978
rect 12394 17926 12406 17978
rect 12458 17926 12470 17978
rect 12522 17926 20214 17978
rect 20266 17926 20278 17978
rect 20330 17926 20342 17978
rect 20394 17926 20406 17978
rect 20458 17926 20470 17978
rect 20522 17926 24840 17978
rect 1104 17904 24840 17926
rect 1670 17824 1676 17876
rect 1728 17864 1734 17876
rect 9122 17864 9128 17876
rect 1728 17836 9128 17864
rect 1728 17824 1734 17836
rect 9122 17824 9128 17836
rect 9180 17824 9186 17876
rect 13725 17867 13783 17873
rect 13725 17833 13737 17867
rect 13771 17864 13783 17867
rect 22462 17864 22468 17876
rect 13771 17836 22468 17864
rect 13771 17833 13783 17836
rect 13725 17827 13783 17833
rect 22462 17824 22468 17836
rect 22520 17824 22526 17876
rect 15286 17756 15292 17808
rect 15344 17796 15350 17808
rect 15749 17799 15807 17805
rect 15749 17796 15761 17799
rect 15344 17768 15761 17796
rect 15344 17756 15350 17768
rect 15749 17765 15761 17768
rect 15795 17765 15807 17799
rect 15749 17759 15807 17765
rect 16758 17756 16764 17808
rect 16816 17796 16822 17808
rect 17494 17796 17500 17808
rect 16816 17768 17500 17796
rect 16816 17756 16822 17768
rect 17494 17756 17500 17768
rect 17552 17756 17558 17808
rect 20622 17756 20628 17808
rect 20680 17756 20686 17808
rect 23198 17756 23204 17808
rect 23256 17756 23262 17808
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 1627 17700 4108 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 4080 17672 4108 17700
rect 4614 17688 4620 17740
rect 4672 17688 4678 17740
rect 5258 17688 5264 17740
rect 5316 17728 5322 17740
rect 6089 17731 6147 17737
rect 6089 17728 6101 17731
rect 5316 17700 6101 17728
rect 5316 17688 5322 17700
rect 6089 17697 6101 17700
rect 6135 17697 6147 17731
rect 6089 17691 6147 17697
rect 8389 17731 8447 17737
rect 8389 17697 8401 17731
rect 8435 17728 8447 17731
rect 8754 17728 8760 17740
rect 8435 17700 8760 17728
rect 8435 17697 8447 17700
rect 8389 17691 8447 17697
rect 8754 17688 8760 17700
rect 8812 17688 8818 17740
rect 10965 17731 11023 17737
rect 10965 17697 10977 17731
rect 11011 17728 11023 17731
rect 11606 17728 11612 17740
rect 11011 17700 11612 17728
rect 11011 17697 11023 17700
rect 10965 17691 11023 17697
rect 11606 17688 11612 17700
rect 11664 17688 11670 17740
rect 17402 17728 17408 17740
rect 15948 17700 17408 17728
rect 4062 17620 4068 17672
rect 4120 17660 4126 17672
rect 4341 17663 4399 17669
rect 4341 17660 4353 17663
rect 4120 17632 4353 17660
rect 4120 17620 4126 17632
rect 4341 17629 4353 17632
rect 4387 17629 4399 17663
rect 4341 17623 4399 17629
rect 5718 17620 5724 17672
rect 5776 17620 5782 17672
rect 8665 17663 8723 17669
rect 8665 17629 8677 17663
rect 8711 17660 8723 17663
rect 9217 17663 9275 17669
rect 9217 17660 9229 17663
rect 8711 17632 9229 17660
rect 8711 17629 8723 17632
rect 8665 17623 8723 17629
rect 9217 17629 9229 17632
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 1857 17595 1915 17601
rect 1857 17561 1869 17595
rect 1903 17592 1915 17595
rect 1946 17592 1952 17604
rect 1903 17564 1952 17592
rect 1903 17561 1915 17564
rect 1857 17555 1915 17561
rect 1946 17552 1952 17564
rect 2004 17552 2010 17604
rect 2590 17552 2596 17604
rect 2648 17552 2654 17604
rect 7926 17552 7932 17604
rect 7984 17552 7990 17604
rect 3326 17484 3332 17536
rect 3384 17484 3390 17536
rect 6917 17527 6975 17533
rect 6917 17493 6929 17527
rect 6963 17524 6975 17527
rect 7374 17524 7380 17536
rect 6963 17496 7380 17524
rect 6963 17493 6975 17496
rect 6917 17487 6975 17493
rect 7374 17484 7380 17496
rect 7432 17484 7438 17536
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8680 17524 8708 17623
rect 10686 17620 10692 17672
rect 10744 17660 10750 17672
rect 11241 17663 11299 17669
rect 11241 17660 11253 17663
rect 10744 17632 11253 17660
rect 10744 17620 10750 17632
rect 11241 17629 11253 17632
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 12710 17620 12716 17672
rect 12768 17660 12774 17672
rect 13081 17663 13139 17669
rect 13081 17660 13093 17663
rect 12768 17632 13093 17660
rect 12768 17620 12774 17632
rect 13081 17629 13093 17632
rect 13127 17629 13139 17663
rect 13081 17623 13139 17629
rect 14458 17620 14464 17672
rect 14516 17620 14522 17672
rect 15948 17669 15976 17700
rect 15933 17663 15991 17669
rect 15933 17629 15945 17663
rect 15979 17629 15991 17663
rect 15933 17623 15991 17629
rect 16114 17620 16120 17672
rect 16172 17660 16178 17672
rect 16301 17663 16359 17669
rect 16301 17660 16313 17663
rect 16172 17632 16313 17660
rect 16172 17620 16178 17632
rect 16301 17629 16313 17632
rect 16347 17629 16359 17663
rect 16301 17623 16359 17629
rect 16942 17620 16948 17672
rect 17000 17620 17006 17672
rect 17236 17669 17264 17700
rect 17402 17688 17408 17700
rect 17460 17728 17466 17740
rect 21361 17731 21419 17737
rect 21361 17728 21373 17731
rect 17460 17700 21373 17728
rect 17460 17688 17466 17700
rect 21361 17697 21373 17700
rect 21407 17697 21419 17731
rect 23216 17728 23244 17756
rect 23216 17700 23796 17728
rect 21361 17691 21419 17697
rect 17221 17663 17279 17669
rect 17221 17629 17233 17663
rect 17267 17629 17279 17663
rect 17221 17623 17279 17629
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 21545 17663 21603 17669
rect 21545 17629 21557 17663
rect 21591 17660 21603 17663
rect 21634 17660 21640 17672
rect 21591 17632 21640 17660
rect 21591 17629 21603 17632
rect 21545 17623 21603 17629
rect 21634 17620 21640 17632
rect 21692 17620 21698 17672
rect 21818 17620 21824 17672
rect 21876 17660 21882 17672
rect 21913 17663 21971 17669
rect 21913 17660 21925 17663
rect 21876 17632 21925 17660
rect 21876 17620 21882 17632
rect 21913 17629 21925 17632
rect 21959 17629 21971 17663
rect 21913 17623 21971 17629
rect 23290 17620 23296 17672
rect 23348 17620 23354 17672
rect 23768 17669 23796 17700
rect 23753 17663 23811 17669
rect 23753 17629 23765 17663
rect 23799 17629 23811 17663
rect 23753 17623 23811 17629
rect 12802 17552 12808 17604
rect 12860 17552 12866 17604
rect 13265 17595 13323 17601
rect 13265 17561 13277 17595
rect 13311 17592 13323 17595
rect 13538 17592 13544 17604
rect 13311 17564 13544 17592
rect 13311 17561 13323 17564
rect 13265 17555 13323 17561
rect 13538 17552 13544 17564
rect 13596 17552 13602 17604
rect 18969 17595 19027 17601
rect 18969 17561 18981 17595
rect 19015 17592 19027 17595
rect 19337 17595 19395 17601
rect 19337 17592 19349 17595
rect 19015 17564 19349 17592
rect 19015 17561 19027 17564
rect 18969 17555 19027 17561
rect 19337 17561 19349 17564
rect 19383 17561 19395 17595
rect 19337 17555 19395 17561
rect 8168 17496 8708 17524
rect 13817 17527 13875 17533
rect 8168 17484 8174 17496
rect 13817 17493 13829 17527
rect 13863 17524 13875 17527
rect 20070 17524 20076 17536
rect 13863 17496 20076 17524
rect 13863 17493 13875 17496
rect 13817 17487 13875 17493
rect 20070 17484 20076 17496
rect 20128 17484 20134 17536
rect 23934 17484 23940 17536
rect 23992 17484 23998 17536
rect 1104 17434 24840 17456
rect 1104 17382 8214 17434
rect 8266 17382 8278 17434
rect 8330 17382 8342 17434
rect 8394 17382 8406 17434
rect 8458 17382 8470 17434
rect 8522 17382 16214 17434
rect 16266 17382 16278 17434
rect 16330 17382 16342 17434
rect 16394 17382 16406 17434
rect 16458 17382 16470 17434
rect 16522 17382 24214 17434
rect 24266 17382 24278 17434
rect 24330 17382 24342 17434
rect 24394 17382 24406 17434
rect 24458 17382 24470 17434
rect 24522 17382 24840 17434
rect 1104 17360 24840 17382
rect 1946 17280 1952 17332
rect 2004 17320 2010 17332
rect 2501 17323 2559 17329
rect 2501 17320 2513 17323
rect 2004 17292 2513 17320
rect 2004 17280 2010 17292
rect 2501 17289 2513 17292
rect 2547 17289 2559 17323
rect 2501 17283 2559 17289
rect 2866 17280 2872 17332
rect 2924 17320 2930 17332
rect 3326 17320 3332 17332
rect 2924 17292 3332 17320
rect 2924 17280 2930 17292
rect 3326 17280 3332 17292
rect 3384 17280 3390 17332
rect 5258 17320 5264 17332
rect 4632 17292 5264 17320
rect 1854 17212 1860 17264
rect 1912 17212 1918 17264
rect 2073 17255 2131 17261
rect 2073 17221 2085 17255
rect 2119 17252 2131 17255
rect 2406 17252 2412 17264
rect 2119 17224 2412 17252
rect 2119 17221 2131 17224
rect 2073 17215 2131 17221
rect 2406 17212 2412 17224
rect 2464 17212 2470 17264
rect 2961 17255 3019 17261
rect 2961 17221 2973 17255
rect 3007 17252 3019 17255
rect 4632 17252 4660 17292
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 8110 17280 8116 17332
rect 8168 17280 8174 17332
rect 8481 17323 8539 17329
rect 8481 17289 8493 17323
rect 8527 17320 8539 17323
rect 8754 17320 8760 17332
rect 8527 17292 8760 17320
rect 8527 17289 8539 17292
rect 8481 17283 8539 17289
rect 8754 17280 8760 17292
rect 8812 17280 8818 17332
rect 9950 17280 9956 17332
rect 10008 17320 10014 17332
rect 10008 17292 16528 17320
rect 10008 17280 10014 17292
rect 3007 17224 4660 17252
rect 3007 17221 3019 17224
rect 2961 17215 3019 17221
rect 4798 17212 4804 17264
rect 4856 17212 4862 17264
rect 8128 17252 8156 17280
rect 10045 17255 10103 17261
rect 8128 17224 8248 17252
rect 6822 17144 6828 17196
rect 6880 17144 6886 17196
rect 8220 17193 8248 17224
rect 10045 17221 10057 17255
rect 10091 17252 10103 17255
rect 10594 17252 10600 17264
rect 10091 17224 10600 17252
rect 10091 17221 10103 17224
rect 10045 17215 10103 17221
rect 10594 17212 10600 17224
rect 10652 17212 10658 17264
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 11241 17255 11299 17261
rect 11241 17252 11253 17255
rect 11204 17224 11253 17252
rect 11204 17212 11210 17224
rect 11241 17221 11253 17224
rect 11287 17221 11299 17255
rect 11241 17215 11299 17221
rect 12066 17212 12072 17264
rect 12124 17252 12130 17264
rect 12253 17255 12311 17261
rect 12253 17252 12265 17255
rect 12124 17224 12265 17252
rect 12124 17212 12130 17224
rect 12253 17221 12265 17224
rect 12299 17221 12311 17255
rect 12253 17215 12311 17221
rect 12529 17255 12587 17261
rect 12529 17221 12541 17255
rect 12575 17252 12587 17255
rect 12710 17252 12716 17264
rect 12575 17224 12716 17252
rect 12575 17221 12587 17224
rect 12529 17215 12587 17221
rect 12710 17212 12716 17224
rect 12768 17212 12774 17264
rect 14366 17212 14372 17264
rect 14424 17252 14430 17264
rect 14921 17255 14979 17261
rect 14921 17252 14933 17255
rect 14424 17224 14933 17252
rect 14424 17212 14430 17224
rect 14921 17221 14933 17224
rect 14967 17252 14979 17255
rect 15933 17255 15991 17261
rect 15933 17252 15945 17255
rect 14967 17224 15945 17252
rect 14967 17221 14979 17224
rect 14921 17215 14979 17221
rect 15933 17221 15945 17224
rect 15979 17221 15991 17255
rect 15933 17215 15991 17221
rect 8205 17187 8263 17193
rect 8205 17153 8217 17187
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 8849 17187 8907 17193
rect 8849 17153 8861 17187
rect 8895 17153 8907 17187
rect 8849 17147 8907 17153
rect 3145 17119 3203 17125
rect 3145 17085 3157 17119
rect 3191 17085 3203 17119
rect 3145 17079 3203 17085
rect 2225 17051 2283 17057
rect 2225 17017 2237 17051
rect 2271 17048 2283 17051
rect 2774 17048 2780 17060
rect 2271 17020 2780 17048
rect 2271 17017 2283 17020
rect 2225 17011 2283 17017
rect 2774 17008 2780 17020
rect 2832 17008 2838 17060
rect 1946 16940 1952 16992
rect 2004 16980 2010 16992
rect 2041 16983 2099 16989
rect 2041 16980 2053 16983
rect 2004 16952 2053 16980
rect 2004 16940 2010 16952
rect 2041 16949 2053 16952
rect 2087 16980 2099 16983
rect 2498 16980 2504 16992
rect 2087 16952 2504 16980
rect 2087 16949 2099 16952
rect 2041 16943 2099 16949
rect 2498 16940 2504 16952
rect 2556 16940 2562 16992
rect 3160 16980 3188 17079
rect 3970 17076 3976 17128
rect 4028 17076 4034 17128
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17116 4307 17119
rect 4706 17116 4712 17128
rect 4295 17088 4712 17116
rect 4295 17085 4307 17088
rect 4249 17079 4307 17085
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 7926 17076 7932 17128
rect 7984 17076 7990 17128
rect 5350 17008 5356 17060
rect 5408 17048 5414 17060
rect 5721 17051 5779 17057
rect 5721 17048 5733 17051
rect 5408 17020 5733 17048
rect 5408 17008 5414 17020
rect 5721 17017 5733 17020
rect 5767 17017 5779 17051
rect 5721 17011 5779 17017
rect 4982 16980 4988 16992
rect 3160 16952 4988 16980
rect 4982 16940 4988 16952
rect 5040 16940 5046 16992
rect 6457 16983 6515 16989
rect 6457 16949 6469 16983
rect 6503 16980 6515 16983
rect 6730 16980 6736 16992
rect 6503 16952 6736 16980
rect 6503 16949 6515 16952
rect 6457 16943 6515 16949
rect 6730 16940 6736 16952
rect 6788 16940 6794 16992
rect 7374 16940 7380 16992
rect 7432 16980 7438 16992
rect 8864 16980 8892 17147
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9953 17187 10011 17193
rect 9953 17184 9965 17187
rect 9364 17156 9965 17184
rect 9364 17144 9370 17156
rect 9953 17153 9965 17156
rect 9999 17153 10011 17187
rect 9953 17147 10011 17153
rect 10226 17144 10232 17196
rect 10284 17144 10290 17196
rect 11606 17144 11612 17196
rect 11664 17144 11670 17196
rect 12805 17187 12863 17193
rect 12805 17153 12817 17187
rect 12851 17184 12863 17187
rect 13078 17184 13084 17196
rect 12851 17156 13084 17184
rect 12851 17153 12863 17156
rect 12805 17147 12863 17153
rect 13078 17144 13084 17156
rect 13136 17144 13142 17196
rect 14274 17144 14280 17196
rect 14332 17184 14338 17196
rect 14642 17184 14648 17196
rect 14332 17156 14648 17184
rect 14332 17144 14338 17156
rect 14642 17144 14648 17156
rect 14700 17144 14706 17196
rect 15562 17144 15568 17196
rect 15620 17184 15626 17196
rect 16393 17187 16451 17193
rect 16393 17184 16405 17187
rect 15620 17156 16405 17184
rect 15620 17144 15626 17156
rect 16393 17153 16405 17156
rect 16439 17153 16451 17187
rect 16500 17184 16528 17292
rect 18322 17280 18328 17332
rect 18380 17320 18386 17332
rect 20349 17323 20407 17329
rect 20349 17320 20361 17323
rect 18380 17292 20361 17320
rect 18380 17280 18386 17292
rect 20349 17289 20361 17292
rect 20395 17289 20407 17323
rect 20349 17283 20407 17289
rect 24118 17280 24124 17332
rect 24176 17320 24182 17332
rect 24305 17323 24363 17329
rect 24305 17320 24317 17323
rect 24176 17292 24317 17320
rect 24176 17280 24182 17292
rect 24305 17289 24317 17292
rect 24351 17320 24363 17323
rect 24578 17320 24584 17332
rect 24351 17292 24584 17320
rect 24351 17289 24363 17292
rect 24305 17283 24363 17289
rect 24578 17280 24584 17292
rect 24636 17280 24642 17332
rect 18690 17212 18696 17264
rect 18748 17252 18754 17264
rect 19429 17255 19487 17261
rect 19429 17252 19441 17255
rect 18748 17224 19441 17252
rect 18748 17212 18754 17224
rect 19429 17221 19441 17224
rect 19475 17252 19487 17255
rect 19981 17255 20039 17261
rect 19981 17252 19993 17255
rect 19475 17224 19993 17252
rect 19475 17221 19487 17224
rect 19429 17215 19487 17221
rect 19981 17221 19993 17224
rect 20027 17221 20039 17255
rect 19981 17215 20039 17221
rect 20070 17212 20076 17264
rect 20128 17252 20134 17264
rect 21085 17255 21143 17261
rect 21085 17252 21097 17255
rect 20128 17224 21097 17252
rect 20128 17212 20134 17224
rect 21085 17221 21097 17224
rect 21131 17252 21143 17255
rect 22649 17255 22707 17261
rect 21131 17224 21496 17252
rect 21131 17221 21143 17224
rect 21085 17215 21143 17221
rect 17129 17187 17187 17193
rect 17129 17184 17141 17187
rect 16500 17156 17141 17184
rect 16393 17147 16451 17153
rect 17129 17153 17141 17156
rect 17175 17153 17187 17187
rect 17129 17147 17187 17153
rect 8938 17076 8944 17128
rect 8996 17076 9002 17128
rect 9030 17076 9036 17128
rect 9088 17076 9094 17128
rect 10686 17076 10692 17128
rect 10744 17076 10750 17128
rect 11149 17119 11207 17125
rect 11149 17085 11161 17119
rect 11195 17116 11207 17119
rect 12710 17116 12716 17128
rect 11195 17088 12716 17116
rect 11195 17085 11207 17088
rect 11149 17079 11207 17085
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 13354 17076 13360 17128
rect 13412 17116 13418 17128
rect 13412 17088 15148 17116
rect 13412 17076 13418 17088
rect 11606 17008 11612 17060
rect 11664 17048 11670 17060
rect 11664 17020 13492 17048
rect 11664 17008 11670 17020
rect 7432 16952 8892 16980
rect 10413 16983 10471 16989
rect 7432 16940 7438 16952
rect 10413 16949 10425 16983
rect 10459 16980 10471 16983
rect 13354 16980 13360 16992
rect 10459 16952 13360 16980
rect 10459 16949 10471 16952
rect 10413 16943 10471 16949
rect 13354 16940 13360 16952
rect 13412 16940 13418 16992
rect 13464 16980 13492 17020
rect 13538 17008 13544 17060
rect 13596 17048 13602 17060
rect 14093 17051 14151 17057
rect 14093 17048 14105 17051
rect 13596 17020 14105 17048
rect 13596 17008 13602 17020
rect 14093 17017 14105 17020
rect 14139 17017 14151 17051
rect 15120 17048 15148 17088
rect 15194 17076 15200 17128
rect 15252 17116 15258 17128
rect 15841 17119 15899 17125
rect 15841 17116 15853 17119
rect 15252 17088 15853 17116
rect 15252 17076 15258 17088
rect 15841 17085 15853 17088
rect 15887 17085 15899 17119
rect 17144 17116 17172 17147
rect 18230 17144 18236 17196
rect 18288 17144 18294 17196
rect 20806 17184 20812 17196
rect 19306 17156 20812 17184
rect 18969 17119 19027 17125
rect 18969 17116 18981 17119
rect 17144 17088 18981 17116
rect 15841 17079 15899 17085
rect 18969 17085 18981 17088
rect 19015 17085 19027 17119
rect 18969 17079 19027 17085
rect 19306 17048 19334 17156
rect 20806 17144 20812 17156
rect 20864 17144 20870 17196
rect 19521 17119 19579 17125
rect 19521 17085 19533 17119
rect 19567 17116 19579 17119
rect 20441 17119 20499 17125
rect 20441 17116 20453 17119
rect 19567 17088 20453 17116
rect 19567 17085 19579 17088
rect 19521 17079 19579 17085
rect 20441 17085 20453 17088
rect 20487 17085 20499 17119
rect 20441 17079 20499 17085
rect 20993 17119 21051 17125
rect 20993 17085 21005 17119
rect 21039 17116 21051 17119
rect 21358 17116 21364 17128
rect 21039 17088 21364 17116
rect 21039 17085 21051 17088
rect 20993 17079 21051 17085
rect 21358 17076 21364 17088
rect 21416 17076 21422 17128
rect 15120 17020 19334 17048
rect 14093 17011 14151 17017
rect 19610 17008 19616 17060
rect 19668 17048 19674 17060
rect 19797 17051 19855 17057
rect 19797 17048 19809 17051
rect 19668 17020 19809 17048
rect 19668 17008 19674 17020
rect 19797 17017 19809 17020
rect 19843 17017 19855 17051
rect 21468 17048 21496 17224
rect 22649 17221 22661 17255
rect 22695 17252 22707 17255
rect 23382 17252 23388 17264
rect 22695 17224 23388 17252
rect 22695 17221 22707 17224
rect 22649 17215 22707 17221
rect 23382 17212 23388 17224
rect 23440 17212 23446 17264
rect 21545 17187 21603 17193
rect 21545 17153 21557 17187
rect 21591 17184 21603 17187
rect 22186 17184 22192 17196
rect 21591 17156 22192 17184
rect 21591 17153 21603 17156
rect 21545 17147 21603 17153
rect 22186 17144 22192 17156
rect 22244 17144 22250 17196
rect 23934 17144 23940 17196
rect 23992 17144 23998 17196
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17116 22155 17119
rect 22462 17116 22468 17128
rect 22143 17088 22468 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 22462 17076 22468 17088
rect 22520 17076 22526 17128
rect 22922 17076 22928 17128
rect 22980 17116 22986 17128
rect 23017 17119 23075 17125
rect 23017 17116 23029 17119
rect 22980 17088 23029 17116
rect 22980 17076 22986 17088
rect 23017 17085 23029 17088
rect 23063 17085 23075 17119
rect 23017 17079 23075 17085
rect 22278 17048 22284 17060
rect 21468 17020 22284 17048
rect 19797 17011 19855 17017
rect 22278 17008 22284 17020
rect 22336 17008 22342 17060
rect 22557 17051 22615 17057
rect 22557 17017 22569 17051
rect 22603 17048 22615 17051
rect 23290 17048 23296 17060
rect 22603 17020 23296 17048
rect 22603 17017 22615 17020
rect 22557 17011 22615 17017
rect 23290 17008 23296 17020
rect 23348 17008 23354 17060
rect 20898 16980 20904 16992
rect 13464 16952 20904 16980
rect 20898 16940 20904 16952
rect 20956 16940 20962 16992
rect 1104 16890 24840 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 12214 16890
rect 12266 16838 12278 16890
rect 12330 16838 12342 16890
rect 12394 16838 12406 16890
rect 12458 16838 12470 16890
rect 12522 16838 20214 16890
rect 20266 16838 20278 16890
rect 20330 16838 20342 16890
rect 20394 16838 20406 16890
rect 20458 16838 20470 16890
rect 20522 16838 24840 16890
rect 1104 16816 24840 16838
rect 4249 16779 4307 16785
rect 4249 16745 4261 16779
rect 4295 16745 4307 16779
rect 4249 16739 4307 16745
rect 1489 16643 1547 16649
rect 1489 16609 1501 16643
rect 1535 16640 1547 16643
rect 4062 16640 4068 16652
rect 1535 16612 4068 16640
rect 1535 16609 1547 16612
rect 1489 16603 1547 16609
rect 4062 16600 4068 16612
rect 4120 16600 4126 16652
rect 4264 16640 4292 16739
rect 4706 16736 4712 16788
rect 4764 16736 4770 16788
rect 5718 16736 5724 16788
rect 5776 16736 5782 16788
rect 5902 16736 5908 16788
rect 5960 16776 5966 16788
rect 6641 16779 6699 16785
rect 6641 16776 6653 16779
rect 5960 16748 6653 16776
rect 5960 16736 5966 16748
rect 6641 16745 6653 16748
rect 6687 16745 6699 16779
rect 6641 16739 6699 16745
rect 6822 16736 6828 16788
rect 6880 16736 6886 16788
rect 7837 16779 7895 16785
rect 7837 16745 7849 16779
rect 7883 16776 7895 16779
rect 7926 16776 7932 16788
rect 7883 16748 7932 16776
rect 7883 16745 7895 16748
rect 7837 16739 7895 16745
rect 7926 16736 7932 16748
rect 7984 16736 7990 16788
rect 8297 16779 8355 16785
rect 8297 16745 8309 16779
rect 8343 16776 8355 16779
rect 8570 16776 8576 16788
rect 8343 16748 8576 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 4433 16711 4491 16717
rect 4433 16677 4445 16711
rect 4479 16708 4491 16711
rect 4798 16708 4804 16720
rect 4479 16680 4804 16708
rect 4479 16677 4491 16680
rect 4433 16671 4491 16677
rect 4798 16668 4804 16680
rect 4856 16668 4862 16720
rect 8312 16708 8340 16739
rect 8570 16736 8576 16748
rect 8628 16736 8634 16788
rect 15105 16779 15163 16785
rect 12406 16748 15056 16776
rect 4908 16680 8340 16708
rect 10413 16711 10471 16717
rect 4908 16640 4936 16680
rect 10413 16677 10425 16711
rect 10459 16708 10471 16711
rect 11054 16708 11060 16720
rect 10459 16680 11060 16708
rect 10459 16677 10471 16680
rect 10413 16671 10471 16677
rect 11054 16668 11060 16680
rect 11112 16668 11118 16720
rect 4264 16612 4936 16640
rect 4982 16600 4988 16652
rect 5040 16640 5046 16652
rect 5261 16643 5319 16649
rect 5261 16640 5273 16643
rect 5040 16612 5273 16640
rect 5040 16600 5046 16612
rect 5261 16609 5273 16612
rect 5307 16640 5319 16643
rect 5442 16640 5448 16652
rect 5307 16612 5448 16640
rect 5307 16609 5319 16612
rect 5261 16603 5319 16609
rect 5442 16600 5448 16612
rect 5500 16600 5506 16652
rect 7190 16600 7196 16652
rect 7248 16600 7254 16652
rect 7374 16600 7380 16652
rect 7432 16600 7438 16652
rect 10873 16643 10931 16649
rect 10873 16609 10885 16643
rect 10919 16640 10931 16643
rect 12406 16640 12434 16748
rect 13538 16668 13544 16720
rect 13596 16668 13602 16720
rect 15028 16708 15056 16748
rect 15105 16745 15117 16779
rect 15151 16776 15163 16779
rect 15562 16776 15568 16788
rect 15151 16748 15568 16776
rect 15151 16745 15163 16748
rect 15105 16739 15163 16745
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 16114 16736 16120 16788
rect 16172 16776 16178 16788
rect 16577 16779 16635 16785
rect 16577 16776 16589 16779
rect 16172 16748 16589 16776
rect 16172 16736 16178 16748
rect 16577 16745 16589 16748
rect 16623 16745 16635 16779
rect 16577 16739 16635 16745
rect 17678 16736 17684 16788
rect 17736 16776 17742 16788
rect 18414 16776 18420 16788
rect 17736 16748 18420 16776
rect 17736 16736 17742 16748
rect 18414 16736 18420 16748
rect 18472 16776 18478 16788
rect 18690 16776 18696 16788
rect 18472 16748 18696 16776
rect 18472 16736 18478 16748
rect 18690 16736 18696 16748
rect 18748 16736 18754 16788
rect 18969 16779 19027 16785
rect 18969 16745 18981 16779
rect 19015 16776 19027 16779
rect 19334 16776 19340 16788
rect 19015 16748 19340 16776
rect 19015 16745 19027 16748
rect 18969 16739 19027 16745
rect 19334 16736 19340 16748
rect 19392 16736 19398 16788
rect 20898 16736 20904 16788
rect 20956 16736 20962 16788
rect 20073 16711 20131 16717
rect 20073 16708 20085 16711
rect 15028 16680 20085 16708
rect 20073 16677 20085 16680
rect 20119 16677 20131 16711
rect 21729 16711 21787 16717
rect 21729 16708 21741 16711
rect 20073 16671 20131 16677
rect 20180 16680 21741 16708
rect 10919 16612 12434 16640
rect 10919 16609 10931 16612
rect 10873 16603 10931 16609
rect 5077 16575 5135 16581
rect 5077 16541 5089 16575
rect 5123 16572 5135 16575
rect 5350 16572 5356 16584
rect 5123 16544 5356 16572
rect 5123 16541 5135 16544
rect 5077 16535 5135 16541
rect 5350 16532 5356 16544
rect 5408 16532 5414 16584
rect 6730 16532 6736 16584
rect 6788 16572 6794 16584
rect 7469 16575 7527 16581
rect 7469 16572 7481 16575
rect 6788 16544 7481 16572
rect 6788 16532 6794 16544
rect 7469 16541 7481 16544
rect 7515 16541 7527 16575
rect 7469 16535 7527 16541
rect 9861 16575 9919 16581
rect 9861 16541 9873 16575
rect 9907 16572 9919 16575
rect 9907 16544 11008 16572
rect 9907 16541 9919 16544
rect 9861 16535 9919 16541
rect 1762 16464 1768 16516
rect 1820 16464 1826 16516
rect 2774 16464 2780 16516
rect 2832 16464 2838 16516
rect 3050 16464 3056 16516
rect 3108 16504 3114 16516
rect 4065 16507 4123 16513
rect 4065 16504 4077 16507
rect 3108 16476 4077 16504
rect 3108 16464 3114 16476
rect 4065 16473 4077 16476
rect 4111 16504 4123 16507
rect 5718 16504 5724 16516
rect 4111 16476 5724 16504
rect 4111 16473 4123 16476
rect 4065 16467 4123 16473
rect 5718 16464 5724 16476
rect 5776 16504 5782 16516
rect 6089 16507 6147 16513
rect 6089 16504 6101 16507
rect 5776 16476 6101 16504
rect 5776 16464 5782 16476
rect 6089 16473 6101 16476
rect 6135 16473 6147 16507
rect 6089 16467 6147 16473
rect 6457 16507 6515 16513
rect 6457 16473 6469 16507
rect 6503 16504 6515 16507
rect 8018 16504 8024 16516
rect 6503 16476 8024 16504
rect 6503 16473 6515 16476
rect 6457 16467 6515 16473
rect 8018 16464 8024 16476
rect 8076 16504 8082 16516
rect 8113 16507 8171 16513
rect 8113 16504 8125 16507
rect 8076 16476 8125 16504
rect 8076 16464 8082 16476
rect 8113 16473 8125 16476
rect 8159 16473 8171 16507
rect 8846 16504 8852 16516
rect 8113 16467 8171 16473
rect 8404 16476 8852 16504
rect 2682 16396 2688 16448
rect 2740 16436 2746 16448
rect 3237 16439 3295 16445
rect 3237 16436 3249 16439
rect 2740 16408 3249 16436
rect 2740 16396 2746 16408
rect 3237 16405 3249 16408
rect 3283 16405 3295 16439
rect 3237 16399 3295 16405
rect 4275 16439 4333 16445
rect 4275 16405 4287 16439
rect 4321 16436 4333 16439
rect 5074 16436 5080 16448
rect 4321 16408 5080 16436
rect 4321 16405 4333 16408
rect 4275 16399 4333 16405
rect 5074 16396 5080 16408
rect 5132 16396 5138 16448
rect 5169 16439 5227 16445
rect 5169 16405 5181 16439
rect 5215 16436 5227 16439
rect 5350 16436 5356 16448
rect 5215 16408 5356 16436
rect 5215 16405 5227 16408
rect 5169 16399 5227 16405
rect 5350 16396 5356 16408
rect 5408 16396 5414 16448
rect 5889 16439 5947 16445
rect 5889 16405 5901 16439
rect 5935 16436 5947 16439
rect 5994 16436 6000 16448
rect 5935 16408 6000 16436
rect 5935 16405 5947 16408
rect 5889 16399 5947 16405
rect 5994 16396 6000 16408
rect 6052 16436 6058 16448
rect 6657 16439 6715 16445
rect 6657 16436 6669 16439
rect 6052 16408 6669 16436
rect 6052 16396 6058 16408
rect 6657 16405 6669 16408
rect 6703 16405 6715 16439
rect 6657 16399 6715 16405
rect 7098 16396 7104 16448
rect 7156 16436 7162 16448
rect 8313 16439 8371 16445
rect 8313 16436 8325 16439
rect 7156 16408 8325 16436
rect 7156 16396 7162 16408
rect 8313 16405 8325 16408
rect 8359 16436 8371 16439
rect 8404 16436 8432 16476
rect 8846 16464 8852 16476
rect 8904 16464 8910 16516
rect 10321 16507 10379 16513
rect 10321 16473 10333 16507
rect 10367 16473 10379 16507
rect 10980 16504 11008 16544
rect 11054 16532 11060 16584
rect 11112 16572 11118 16584
rect 12084 16581 12112 16612
rect 13078 16600 13084 16652
rect 13136 16600 13142 16652
rect 17954 16640 17960 16652
rect 15672 16612 16160 16640
rect 11333 16575 11391 16581
rect 11333 16572 11345 16575
rect 11112 16544 11345 16572
rect 11112 16532 11118 16544
rect 11333 16541 11345 16544
rect 11379 16541 11391 16575
rect 11333 16535 11391 16541
rect 12069 16575 12127 16581
rect 12069 16541 12081 16575
rect 12115 16541 12127 16575
rect 12069 16535 12127 16541
rect 12437 16575 12495 16581
rect 12437 16541 12449 16575
rect 12483 16572 12495 16575
rect 12802 16572 12808 16584
rect 12483 16544 12808 16572
rect 12483 16541 12495 16544
rect 12437 16535 12495 16541
rect 12802 16532 12808 16544
rect 12860 16532 12866 16584
rect 14366 16532 14372 16584
rect 14424 16532 14430 16584
rect 14642 16532 14648 16584
rect 14700 16532 14706 16584
rect 15286 16532 15292 16584
rect 15344 16532 15350 16584
rect 15473 16575 15531 16581
rect 15473 16541 15485 16575
rect 15519 16572 15531 16575
rect 15672 16572 15700 16612
rect 16132 16584 16160 16612
rect 16408 16612 17960 16640
rect 15519 16544 15700 16572
rect 15749 16575 15807 16581
rect 15519 16541 15531 16544
rect 15473 16535 15531 16541
rect 15749 16541 15761 16575
rect 15795 16572 15807 16575
rect 15838 16572 15844 16584
rect 15795 16544 15844 16572
rect 15795 16541 15807 16544
rect 15749 16535 15807 16541
rect 15838 16532 15844 16544
rect 15896 16532 15902 16584
rect 16022 16532 16028 16584
rect 16080 16532 16086 16584
rect 16114 16532 16120 16584
rect 16172 16572 16178 16584
rect 16408 16581 16436 16612
rect 17954 16600 17960 16612
rect 18012 16600 18018 16652
rect 19337 16643 19395 16649
rect 19337 16640 19349 16643
rect 18616 16612 19349 16640
rect 16209 16575 16267 16581
rect 16209 16572 16221 16575
rect 16172 16544 16221 16572
rect 16172 16532 16178 16544
rect 16209 16541 16221 16544
rect 16255 16541 16267 16575
rect 16209 16535 16267 16541
rect 16393 16575 16451 16581
rect 16393 16541 16405 16575
rect 16439 16541 16451 16575
rect 16393 16535 16451 16541
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16541 17279 16575
rect 17221 16535 17279 16541
rect 11149 16507 11207 16513
rect 11149 16504 11161 16507
rect 10980 16476 11161 16504
rect 10321 16467 10379 16473
rect 11149 16473 11161 16476
rect 11195 16504 11207 16507
rect 11195 16476 12434 16504
rect 11195 16473 11207 16476
rect 11149 16467 11207 16473
rect 8359 16408 8432 16436
rect 8481 16439 8539 16445
rect 8359 16405 8371 16408
rect 8313 16399 8371 16405
rect 8481 16405 8493 16439
rect 8527 16436 8539 16439
rect 8570 16436 8576 16448
rect 8527 16408 8576 16436
rect 8527 16405 8539 16408
rect 8481 16399 8539 16405
rect 8570 16396 8576 16408
rect 8628 16396 8634 16448
rect 10045 16439 10103 16445
rect 10045 16405 10057 16439
rect 10091 16436 10103 16439
rect 10336 16436 10364 16467
rect 10091 16408 10364 16436
rect 12406 16436 12434 16476
rect 12618 16464 12624 16516
rect 12676 16464 12682 16516
rect 13633 16507 13691 16513
rect 13633 16473 13645 16507
rect 13679 16504 13691 16507
rect 14185 16507 14243 16513
rect 14185 16504 14197 16507
rect 13679 16476 14197 16504
rect 13679 16473 13691 16476
rect 13633 16467 13691 16473
rect 14185 16473 14197 16476
rect 14231 16473 14243 16507
rect 15194 16504 15200 16516
rect 14185 16467 14243 16473
rect 14844 16476 15200 16504
rect 12636 16436 12664 16464
rect 14844 16445 14872 16476
rect 15194 16464 15200 16476
rect 15252 16464 15258 16516
rect 15654 16513 15660 16516
rect 15381 16507 15439 16513
rect 15381 16473 15393 16507
rect 15427 16473 15439 16507
rect 15381 16467 15439 16473
rect 15611 16507 15660 16513
rect 15611 16473 15623 16507
rect 15657 16473 15660 16507
rect 15611 16467 15660 16473
rect 12406 16408 12664 16436
rect 14829 16439 14887 16445
rect 10091 16405 10103 16408
rect 10045 16399 10103 16405
rect 14829 16405 14841 16439
rect 14875 16405 14887 16439
rect 15396 16436 15424 16467
rect 15654 16464 15660 16467
rect 15712 16464 15718 16516
rect 15856 16504 15884 16532
rect 16301 16507 16359 16513
rect 16301 16504 16313 16507
rect 15856 16476 16313 16504
rect 16301 16473 16313 16476
rect 16347 16473 16359 16507
rect 17236 16504 17264 16535
rect 17678 16532 17684 16584
rect 17736 16532 17742 16584
rect 18230 16572 18236 16584
rect 17804 16544 18236 16572
rect 17804 16504 17832 16544
rect 18230 16532 18236 16544
rect 18288 16572 18294 16584
rect 18616 16581 18644 16612
rect 19337 16609 19349 16612
rect 19383 16609 19395 16643
rect 20180 16640 20208 16680
rect 21729 16677 21741 16680
rect 21775 16677 21787 16711
rect 21729 16671 21787 16677
rect 23290 16668 23296 16720
rect 23348 16708 23354 16720
rect 23753 16711 23811 16717
rect 23753 16708 23765 16711
rect 23348 16680 23765 16708
rect 23348 16668 23354 16680
rect 23753 16677 23765 16680
rect 23799 16677 23811 16711
rect 23753 16671 23811 16677
rect 19337 16603 19395 16609
rect 19444 16612 20208 16640
rect 20548 16612 21496 16640
rect 18601 16575 18659 16581
rect 18601 16572 18613 16575
rect 18288 16544 18613 16572
rect 18288 16532 18294 16544
rect 18601 16541 18613 16544
rect 18647 16541 18659 16575
rect 18601 16535 18659 16541
rect 18690 16532 18696 16584
rect 18748 16572 18754 16584
rect 19444 16572 19472 16612
rect 18748 16544 19472 16572
rect 18748 16532 18754 16544
rect 19978 16532 19984 16584
rect 20036 16572 20042 16584
rect 20548 16581 20576 16612
rect 20257 16575 20315 16581
rect 20257 16572 20269 16575
rect 20036 16544 20269 16572
rect 20036 16532 20042 16544
rect 20257 16541 20269 16544
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20349 16575 20407 16581
rect 20349 16541 20361 16575
rect 20395 16541 20407 16575
rect 20349 16535 20407 16541
rect 20533 16575 20591 16581
rect 20533 16541 20545 16575
rect 20579 16541 20591 16575
rect 20533 16535 20591 16541
rect 17236 16476 17832 16504
rect 16301 16467 16359 16473
rect 18322 16464 18328 16516
rect 18380 16464 18386 16516
rect 19518 16464 19524 16516
rect 19576 16464 19582 16516
rect 16022 16436 16028 16448
rect 15396 16408 16028 16436
rect 14829 16399 14887 16405
rect 16022 16396 16028 16408
rect 16080 16396 16086 16448
rect 17405 16439 17463 16445
rect 17405 16405 17417 16439
rect 17451 16436 17463 16439
rect 17862 16436 17868 16448
rect 17451 16408 17868 16436
rect 17451 16405 17463 16408
rect 17405 16399 17463 16405
rect 17862 16396 17868 16408
rect 17920 16396 17926 16448
rect 17954 16396 17960 16448
rect 18012 16436 18018 16448
rect 19426 16436 19432 16448
rect 18012 16408 19432 16436
rect 18012 16396 18018 16408
rect 19426 16396 19432 16408
rect 19484 16396 19490 16448
rect 20364 16436 20392 16535
rect 20622 16532 20628 16584
rect 20680 16532 20686 16584
rect 21082 16532 21088 16584
rect 21140 16532 21146 16584
rect 21174 16532 21180 16584
rect 21232 16532 21238 16584
rect 21468 16581 21496 16612
rect 21453 16575 21511 16581
rect 21453 16541 21465 16575
rect 21499 16572 21511 16575
rect 21542 16572 21548 16584
rect 21499 16544 21548 16572
rect 21499 16541 21511 16544
rect 21453 16535 21511 16541
rect 21542 16532 21548 16544
rect 21600 16572 21606 16584
rect 21913 16575 21971 16581
rect 21913 16572 21925 16575
rect 21600 16544 21925 16572
rect 21600 16532 21606 16544
rect 21913 16541 21925 16544
rect 21959 16541 21971 16575
rect 21913 16535 21971 16541
rect 22189 16575 22247 16581
rect 22189 16541 22201 16575
rect 22235 16572 22247 16575
rect 22370 16572 22376 16584
rect 22235 16544 22376 16572
rect 22235 16541 22247 16544
rect 22189 16535 22247 16541
rect 22370 16532 22376 16544
rect 22428 16532 22434 16584
rect 22462 16532 22468 16584
rect 22520 16532 22526 16584
rect 23385 16575 23443 16581
rect 23385 16541 23397 16575
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 21266 16464 21272 16516
rect 21324 16464 21330 16516
rect 21726 16464 21732 16516
rect 21784 16504 21790 16516
rect 23400 16504 23428 16535
rect 23566 16504 23572 16516
rect 21784 16476 23572 16504
rect 21784 16464 21790 16476
rect 23566 16464 23572 16476
rect 23624 16464 23630 16516
rect 21174 16436 21180 16448
rect 20364 16408 21180 16436
rect 21174 16396 21180 16408
rect 21232 16436 21238 16448
rect 22097 16439 22155 16445
rect 22097 16436 22109 16439
rect 21232 16408 22109 16436
rect 21232 16396 21238 16408
rect 22097 16405 22109 16408
rect 22143 16405 22155 16439
rect 22097 16399 22155 16405
rect 1104 16346 24840 16368
rect 1104 16294 8214 16346
rect 8266 16294 8278 16346
rect 8330 16294 8342 16346
rect 8394 16294 8406 16346
rect 8458 16294 8470 16346
rect 8522 16294 16214 16346
rect 16266 16294 16278 16346
rect 16330 16294 16342 16346
rect 16394 16294 16406 16346
rect 16458 16294 16470 16346
rect 16522 16294 24214 16346
rect 24266 16294 24278 16346
rect 24330 16294 24342 16346
rect 24394 16294 24406 16346
rect 24458 16294 24470 16346
rect 24522 16294 24840 16346
rect 1104 16272 24840 16294
rect 1762 16192 1768 16244
rect 1820 16232 1826 16244
rect 2317 16235 2375 16241
rect 2317 16232 2329 16235
rect 1820 16204 2329 16232
rect 1820 16192 1826 16204
rect 2317 16201 2329 16204
rect 2363 16201 2375 16235
rect 2317 16195 2375 16201
rect 2682 16192 2688 16244
rect 2740 16192 2746 16244
rect 2777 16235 2835 16241
rect 2777 16201 2789 16235
rect 2823 16232 2835 16235
rect 2866 16232 2872 16244
rect 2823 16204 2872 16232
rect 2823 16201 2835 16204
rect 2777 16195 2835 16201
rect 2866 16192 2872 16204
rect 2924 16192 2930 16244
rect 4982 16232 4988 16244
rect 2976 16204 4988 16232
rect 2130 16124 2136 16176
rect 2188 16164 2194 16176
rect 2188 16136 2912 16164
rect 2188 16124 2194 16136
rect 2884 16108 2912 16136
rect 1486 16056 1492 16108
rect 1544 16096 1550 16108
rect 1949 16099 2007 16105
rect 1949 16096 1961 16099
rect 1544 16068 1961 16096
rect 1544 16056 1550 16068
rect 1949 16065 1961 16068
rect 1995 16065 2007 16099
rect 1949 16059 2007 16065
rect 2866 16056 2872 16108
rect 2924 16056 2930 16108
rect 2976 16037 3004 16204
rect 4982 16192 4988 16204
rect 5040 16192 5046 16244
rect 5074 16192 5080 16244
rect 5132 16232 5138 16244
rect 7098 16232 7104 16244
rect 5132 16204 7104 16232
rect 5132 16192 5138 16204
rect 7098 16192 7104 16204
rect 7156 16192 7162 16244
rect 8110 16232 8116 16244
rect 7208 16204 8116 16232
rect 4062 16164 4068 16176
rect 3896 16136 4068 16164
rect 3896 16105 3924 16136
rect 4062 16124 4068 16136
rect 4120 16124 4126 16176
rect 3881 16099 3939 16105
rect 3881 16065 3893 16099
rect 3927 16065 3939 16099
rect 3881 16059 3939 16065
rect 5258 16056 5264 16108
rect 5316 16056 5322 16108
rect 7098 16056 7104 16108
rect 7156 16096 7162 16108
rect 7208 16105 7236 16204
rect 8110 16192 8116 16204
rect 8168 16192 8174 16244
rect 8938 16192 8944 16244
rect 8996 16192 9002 16244
rect 10581 16235 10639 16241
rect 10581 16201 10593 16235
rect 10627 16232 10639 16235
rect 10627 16204 11008 16232
rect 10627 16201 10639 16204
rect 10581 16195 10639 16201
rect 9674 16124 9680 16176
rect 9732 16164 9738 16176
rect 10781 16167 10839 16173
rect 10781 16164 10793 16167
rect 9732 16136 10793 16164
rect 9732 16124 9738 16136
rect 10781 16133 10793 16136
rect 10827 16133 10839 16167
rect 10980 16164 11008 16204
rect 11054 16192 11060 16244
rect 11112 16192 11118 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14461 16235 14519 16241
rect 14461 16232 14473 16235
rect 13872 16204 14473 16232
rect 13872 16192 13878 16204
rect 14461 16201 14473 16204
rect 14507 16201 14519 16235
rect 14461 16195 14519 16201
rect 15933 16235 15991 16241
rect 15933 16201 15945 16235
rect 15979 16232 15991 16235
rect 16022 16232 16028 16244
rect 15979 16204 16028 16232
rect 15979 16201 15991 16204
rect 15933 16195 15991 16201
rect 16022 16192 16028 16204
rect 16080 16192 16086 16244
rect 17681 16235 17739 16241
rect 17681 16201 17693 16235
rect 17727 16232 17739 16235
rect 18414 16232 18420 16244
rect 17727 16204 18420 16232
rect 17727 16201 17739 16204
rect 17681 16195 17739 16201
rect 18414 16192 18420 16204
rect 18472 16232 18478 16244
rect 20165 16235 20223 16241
rect 18472 16204 18920 16232
rect 18472 16192 18478 16204
rect 11146 16164 11152 16176
rect 10980 16136 11152 16164
rect 10781 16127 10839 16133
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 18892 16173 18920 16204
rect 20165 16201 20177 16235
rect 20211 16232 20223 16235
rect 21266 16232 21272 16244
rect 20211 16204 21272 16232
rect 20211 16201 20223 16204
rect 20165 16195 20223 16201
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 23658 16192 23664 16244
rect 23716 16232 23722 16244
rect 24213 16235 24271 16241
rect 24213 16232 24225 16235
rect 23716 16204 24225 16232
rect 23716 16192 23722 16204
rect 24213 16201 24225 16204
rect 24259 16201 24271 16235
rect 24213 16195 24271 16201
rect 17589 16167 17647 16173
rect 17589 16133 17601 16167
rect 17635 16164 17647 16167
rect 18509 16167 18567 16173
rect 18509 16164 18521 16167
rect 17635 16136 18521 16164
rect 17635 16133 17647 16136
rect 17589 16127 17647 16133
rect 18509 16133 18521 16136
rect 18555 16133 18567 16167
rect 18509 16127 18567 16133
rect 18877 16167 18935 16173
rect 18877 16133 18889 16167
rect 18923 16133 18935 16167
rect 18877 16127 18935 16133
rect 18966 16124 18972 16176
rect 19024 16164 19030 16176
rect 21726 16164 21732 16176
rect 19024 16136 19656 16164
rect 19024 16124 19030 16136
rect 7193 16099 7251 16105
rect 7193 16096 7205 16099
rect 7156 16068 7205 16096
rect 7156 16056 7162 16068
rect 7193 16065 7205 16068
rect 7239 16065 7251 16099
rect 7193 16059 7251 16065
rect 8570 16056 8576 16108
rect 8628 16056 8634 16108
rect 11606 16056 11612 16108
rect 11664 16056 11670 16108
rect 12618 16056 12624 16108
rect 12676 16056 12682 16108
rect 13262 16056 13268 16108
rect 13320 16096 13326 16108
rect 13541 16099 13599 16105
rect 13541 16096 13553 16099
rect 13320 16068 13553 16096
rect 13320 16056 13326 16068
rect 13541 16065 13553 16068
rect 13587 16065 13599 16099
rect 13541 16059 13599 16065
rect 13722 16056 13728 16108
rect 13780 16056 13786 16108
rect 13817 16099 13875 16105
rect 13817 16065 13829 16099
rect 13863 16065 13875 16099
rect 13817 16059 13875 16065
rect 2961 16031 3019 16037
rect 2961 15997 2973 16031
rect 3007 15997 3019 16031
rect 2961 15991 3019 15997
rect 4157 16031 4215 16037
rect 4157 15997 4169 16031
rect 4203 16028 4215 16031
rect 4614 16028 4620 16040
rect 4203 16000 4620 16028
rect 4203 15997 4215 16000
rect 4157 15991 4215 15997
rect 4614 15988 4620 16000
rect 4672 15988 4678 16040
rect 7469 16031 7527 16037
rect 7469 15997 7481 16031
rect 7515 16028 7527 16031
rect 7926 16028 7932 16040
rect 7515 16000 7932 16028
rect 7515 15997 7527 16000
rect 7469 15991 7527 15997
rect 7926 15988 7932 16000
rect 7984 15988 7990 16040
rect 8018 15988 8024 16040
rect 8076 16028 8082 16040
rect 9674 16028 9680 16040
rect 8076 16000 9680 16028
rect 8076 15988 8082 16000
rect 9674 15988 9680 16000
rect 9732 15988 9738 16040
rect 13354 15988 13360 16040
rect 13412 16028 13418 16040
rect 13832 16028 13860 16059
rect 13906 16056 13912 16108
rect 13964 16105 13970 16108
rect 13964 16059 13972 16105
rect 13964 16056 13970 16059
rect 15102 16056 15108 16108
rect 15160 16096 15166 16108
rect 15381 16099 15439 16105
rect 15381 16096 15393 16099
rect 15160 16068 15393 16096
rect 15160 16056 15166 16068
rect 15381 16065 15393 16068
rect 15427 16065 15439 16099
rect 15381 16059 15439 16065
rect 15470 16056 15476 16108
rect 15528 16096 15534 16108
rect 15749 16099 15807 16105
rect 15749 16096 15761 16099
rect 15528 16068 15761 16096
rect 15528 16056 15534 16068
rect 15749 16065 15761 16068
rect 15795 16096 15807 16099
rect 16574 16096 16580 16108
rect 15795 16068 16580 16096
rect 15795 16065 15807 16068
rect 15749 16059 15807 16065
rect 16574 16056 16580 16068
rect 16632 16056 16638 16108
rect 17221 16099 17279 16105
rect 17221 16065 17233 16099
rect 17267 16096 17279 16099
rect 18230 16096 18236 16108
rect 17267 16068 18236 16096
rect 17267 16065 17279 16068
rect 17221 16059 17279 16065
rect 18230 16056 18236 16068
rect 18288 16056 18294 16108
rect 18417 16099 18475 16105
rect 18417 16065 18429 16099
rect 18463 16096 18475 16099
rect 18598 16096 18604 16108
rect 18463 16068 18604 16096
rect 18463 16065 18475 16068
rect 18417 16059 18475 16065
rect 18598 16056 18604 16068
rect 18656 16096 18662 16108
rect 19518 16096 19524 16108
rect 18656 16068 19524 16096
rect 18656 16056 18662 16068
rect 19518 16056 19524 16068
rect 19576 16056 19582 16108
rect 19628 16105 19656 16136
rect 20456 16136 21732 16164
rect 20456 16105 20484 16136
rect 21726 16124 21732 16136
rect 21784 16124 21790 16176
rect 22278 16124 22284 16176
rect 22336 16164 22342 16176
rect 22833 16167 22891 16173
rect 22833 16164 22845 16167
rect 22336 16136 22845 16164
rect 22336 16124 22342 16136
rect 22833 16133 22845 16136
rect 22879 16133 22891 16167
rect 22833 16127 22891 16133
rect 23474 16124 23480 16176
rect 23532 16124 23538 16176
rect 19613 16099 19671 16105
rect 19613 16065 19625 16099
rect 19659 16065 19671 16099
rect 19613 16059 19671 16065
rect 20441 16099 20499 16105
rect 20441 16065 20453 16099
rect 20487 16065 20499 16099
rect 20441 16059 20499 16065
rect 20714 16056 20720 16108
rect 20772 16096 20778 16108
rect 20901 16099 20959 16105
rect 20901 16096 20913 16099
rect 20772 16068 20913 16096
rect 20772 16056 20778 16068
rect 20901 16065 20913 16068
rect 20947 16065 20959 16099
rect 20901 16059 20959 16065
rect 20990 16056 20996 16108
rect 21048 16096 21054 16108
rect 21085 16099 21143 16105
rect 21085 16096 21097 16099
rect 21048 16068 21097 16096
rect 21048 16056 21054 16068
rect 21085 16065 21097 16068
rect 21131 16065 21143 16099
rect 21085 16059 21143 16065
rect 21174 16056 21180 16108
rect 21232 16056 21238 16108
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16096 21327 16099
rect 21450 16096 21456 16108
rect 21315 16068 21456 16096
rect 21315 16065 21327 16068
rect 21269 16059 21327 16065
rect 21450 16056 21456 16068
rect 21508 16056 21514 16108
rect 22186 16056 22192 16108
rect 22244 16056 22250 16108
rect 23106 16056 23112 16108
rect 23164 16056 23170 16108
rect 23198 16056 23204 16108
rect 23256 16096 23262 16108
rect 23937 16099 23995 16105
rect 23937 16096 23949 16099
rect 23256 16068 23949 16096
rect 23256 16056 23262 16068
rect 23937 16065 23949 16068
rect 23983 16065 23995 16099
rect 23937 16059 23995 16065
rect 24213 16099 24271 16105
rect 24213 16065 24225 16099
rect 24259 16065 24271 16099
rect 24213 16059 24271 16065
rect 24397 16099 24455 16105
rect 24397 16065 24409 16099
rect 24443 16096 24455 16099
rect 24670 16096 24676 16108
rect 24443 16068 24676 16096
rect 24443 16065 24455 16068
rect 24397 16059 24455 16065
rect 15838 16028 15844 16040
rect 13412 16000 15844 16028
rect 13412 15988 13418 16000
rect 15838 15988 15844 16000
rect 15896 16028 15902 16040
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 15896 16000 16957 16028
rect 15896 15988 15902 16000
rect 16945 15997 16957 16000
rect 16991 16028 17003 16031
rect 17034 16028 17040 16040
rect 16991 16000 17040 16028
rect 16991 15997 17003 16000
rect 16945 15991 17003 15997
rect 17034 15988 17040 16000
rect 17092 15988 17098 16040
rect 17310 15988 17316 16040
rect 17368 16028 17374 16040
rect 17957 16031 18015 16037
rect 17957 16028 17969 16031
rect 17368 16000 17969 16028
rect 17368 15988 17374 16000
rect 17957 15997 17969 16000
rect 18003 15997 18015 16031
rect 17957 15991 18015 15997
rect 18782 15988 18788 16040
rect 18840 15988 18846 16040
rect 19334 15988 19340 16040
rect 19392 15988 19398 16040
rect 19886 15988 19892 16040
rect 19944 15988 19950 16040
rect 23385 16031 23443 16037
rect 23385 15997 23397 16031
rect 23431 15997 23443 16031
rect 23385 15991 23443 15997
rect 5350 15920 5356 15972
rect 5408 15960 5414 15972
rect 5629 15963 5687 15969
rect 5629 15960 5641 15963
rect 5408 15932 5641 15960
rect 5408 15920 5414 15932
rect 5629 15929 5641 15932
rect 5675 15929 5687 15963
rect 5629 15923 5687 15929
rect 10318 15920 10324 15972
rect 10376 15960 10382 15972
rect 10376 15932 10640 15960
rect 10376 15920 10382 15932
rect 1673 15895 1731 15901
rect 1673 15861 1685 15895
rect 1719 15892 1731 15895
rect 5442 15892 5448 15904
rect 1719 15864 5448 15892
rect 1719 15861 1731 15864
rect 1673 15855 1731 15861
rect 5442 15852 5448 15864
rect 5500 15852 5506 15904
rect 10134 15852 10140 15904
rect 10192 15892 10198 15904
rect 10612 15901 10640 15932
rect 12894 15920 12900 15972
rect 12952 15920 12958 15972
rect 14093 15963 14151 15969
rect 14093 15929 14105 15963
rect 14139 15960 14151 15963
rect 18690 15960 18696 15972
rect 14139 15932 18696 15960
rect 14139 15929 14151 15932
rect 14093 15923 14151 15929
rect 18690 15920 18696 15932
rect 18748 15920 18754 15972
rect 19794 15960 19800 15972
rect 18800 15932 19800 15960
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 10192 15864 10425 15892
rect 10192 15852 10198 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 10597 15895 10655 15901
rect 10597 15861 10609 15895
rect 10643 15861 10655 15895
rect 10597 15855 10655 15861
rect 11149 15895 11207 15901
rect 11149 15861 11161 15895
rect 11195 15892 11207 15895
rect 11974 15892 11980 15904
rect 11195 15864 11980 15892
rect 11195 15861 11207 15864
rect 11149 15855 11207 15861
rect 11974 15852 11980 15864
rect 12032 15852 12038 15904
rect 15562 15852 15568 15904
rect 15620 15852 15626 15904
rect 15654 15852 15660 15904
rect 15712 15892 15718 15904
rect 18800 15892 18828 15932
rect 19794 15920 19800 15932
rect 19852 15920 19858 15972
rect 20625 15963 20683 15969
rect 20625 15929 20637 15963
rect 20671 15960 20683 15963
rect 23400 15960 23428 15991
rect 20671 15932 23428 15960
rect 20671 15929 20683 15932
rect 20625 15923 20683 15929
rect 15712 15864 18828 15892
rect 15712 15852 15718 15864
rect 19978 15852 19984 15904
rect 20036 15852 20042 15904
rect 20990 15852 20996 15904
rect 21048 15892 21054 15904
rect 21174 15892 21180 15904
rect 21048 15864 21180 15892
rect 21048 15852 21054 15864
rect 21174 15852 21180 15864
rect 21232 15852 21238 15904
rect 21450 15852 21456 15904
rect 21508 15852 21514 15904
rect 23290 15852 23296 15904
rect 23348 15892 23354 15904
rect 24228 15892 24256 16059
rect 24670 16056 24676 16068
rect 24728 16056 24734 16108
rect 23348 15864 24256 15892
rect 23348 15852 23354 15864
rect 1104 15802 24840 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 12214 15802
rect 12266 15750 12278 15802
rect 12330 15750 12342 15802
rect 12394 15750 12406 15802
rect 12458 15750 12470 15802
rect 12522 15750 20214 15802
rect 20266 15750 20278 15802
rect 20330 15750 20342 15802
rect 20394 15750 20406 15802
rect 20458 15750 20470 15802
rect 20522 15750 24840 15802
rect 1104 15728 24840 15750
rect 4341 15691 4399 15697
rect 4341 15657 4353 15691
rect 4387 15688 4399 15691
rect 4614 15688 4620 15700
rect 4387 15660 4620 15688
rect 4387 15657 4399 15660
rect 4341 15651 4399 15657
rect 4614 15648 4620 15660
rect 4672 15648 4678 15700
rect 5258 15648 5264 15700
rect 5316 15688 5322 15700
rect 5353 15691 5411 15697
rect 5353 15688 5365 15691
rect 5316 15660 5365 15688
rect 5316 15648 5322 15660
rect 5353 15657 5365 15660
rect 5399 15657 5411 15691
rect 5353 15651 5411 15657
rect 5537 15691 5595 15697
rect 5537 15657 5549 15691
rect 5583 15688 5595 15691
rect 5902 15688 5908 15700
rect 5583 15660 5908 15688
rect 5583 15657 5595 15660
rect 5537 15651 5595 15657
rect 5902 15648 5908 15660
rect 5960 15648 5966 15700
rect 7926 15648 7932 15700
rect 7984 15648 7990 15700
rect 14826 15648 14832 15700
rect 14884 15648 14890 15700
rect 15194 15648 15200 15700
rect 15252 15688 15258 15700
rect 15933 15691 15991 15697
rect 15252 15660 15700 15688
rect 15252 15648 15258 15660
rect 2884 15592 5396 15620
rect 2682 15512 2688 15564
rect 2740 15512 2746 15564
rect 2884 15561 2912 15592
rect 2869 15555 2927 15561
rect 2869 15521 2881 15555
rect 2915 15521 2927 15555
rect 2869 15515 2927 15521
rect 4982 15512 4988 15564
rect 5040 15512 5046 15564
rect 5368 15552 5396 15592
rect 5442 15580 5448 15632
rect 5500 15620 5506 15632
rect 13814 15620 13820 15632
rect 5500 15592 13820 15620
rect 5500 15580 5506 15592
rect 13814 15580 13820 15592
rect 13872 15580 13878 15632
rect 15010 15580 15016 15632
rect 15068 15620 15074 15632
rect 15672 15629 15700 15660
rect 15933 15657 15945 15691
rect 15979 15688 15991 15691
rect 16114 15688 16120 15700
rect 15979 15660 16120 15688
rect 15979 15657 15991 15660
rect 15933 15651 15991 15657
rect 16114 15648 16120 15660
rect 16172 15648 16178 15700
rect 16574 15688 16580 15700
rect 16500 15660 16580 15688
rect 15565 15623 15623 15629
rect 15565 15620 15577 15623
rect 15068 15592 15577 15620
rect 15068 15580 15074 15592
rect 15565 15589 15577 15592
rect 15611 15589 15623 15623
rect 15565 15583 15623 15589
rect 15657 15623 15715 15629
rect 15657 15589 15669 15623
rect 15703 15589 15715 15623
rect 15657 15583 15715 15589
rect 6549 15555 6607 15561
rect 6549 15552 6561 15555
rect 5368 15524 6561 15552
rect 6549 15521 6561 15524
rect 6595 15552 6607 15555
rect 7190 15552 7196 15564
rect 6595 15524 7196 15552
rect 6595 15521 6607 15524
rect 6549 15515 6607 15521
rect 7190 15512 7196 15524
rect 7248 15552 7254 15564
rect 8481 15555 8539 15561
rect 8481 15552 8493 15555
rect 7248 15524 8493 15552
rect 7248 15512 7254 15524
rect 8481 15521 8493 15524
rect 8527 15552 8539 15555
rect 8570 15552 8576 15564
rect 8527 15524 8576 15552
rect 8527 15521 8539 15524
rect 8481 15515 8539 15521
rect 8570 15512 8576 15524
rect 8628 15552 8634 15564
rect 9030 15552 9036 15564
rect 8628 15524 9036 15552
rect 8628 15512 8634 15524
rect 9030 15512 9036 15524
rect 9088 15512 9094 15564
rect 11606 15512 11612 15564
rect 11664 15512 11670 15564
rect 11974 15512 11980 15564
rect 12032 15552 12038 15564
rect 12161 15555 12219 15561
rect 12161 15552 12173 15555
rect 12032 15524 12173 15552
rect 12032 15512 12038 15524
rect 12161 15521 12173 15524
rect 12207 15521 12219 15555
rect 12161 15515 12219 15521
rect 15102 15512 15108 15564
rect 15160 15552 15166 15564
rect 15160 15524 16252 15552
rect 15160 15512 15166 15524
rect 4709 15487 4767 15493
rect 4709 15453 4721 15487
rect 4755 15484 4767 15487
rect 5350 15484 5356 15496
rect 4755 15456 5356 15484
rect 4755 15453 4767 15456
rect 4709 15447 4767 15453
rect 5350 15444 5356 15456
rect 5408 15444 5414 15496
rect 5994 15484 6000 15496
rect 5552 15456 6000 15484
rect 5552 15425 5580 15456
rect 5994 15444 6000 15456
rect 6052 15444 6058 15496
rect 6457 15487 6515 15493
rect 6457 15453 6469 15487
rect 6503 15484 6515 15487
rect 6730 15484 6736 15496
rect 6503 15456 6736 15484
rect 6503 15453 6515 15456
rect 6457 15447 6515 15453
rect 6730 15444 6736 15456
rect 6788 15444 6794 15496
rect 8297 15487 8355 15493
rect 8297 15453 8309 15487
rect 8343 15484 8355 15487
rect 8938 15484 8944 15496
rect 8343 15456 8944 15484
rect 8343 15453 8355 15456
rect 8297 15447 8355 15453
rect 8938 15444 8944 15456
rect 8996 15444 9002 15496
rect 10226 15444 10232 15496
rect 10284 15444 10290 15496
rect 10318 15444 10324 15496
rect 10376 15484 10382 15496
rect 10376 15456 10421 15484
rect 10376 15444 10382 15456
rect 10594 15444 10600 15496
rect 10652 15444 10658 15496
rect 10735 15487 10793 15493
rect 10735 15453 10747 15487
rect 10781 15484 10793 15487
rect 10870 15484 10876 15496
rect 10781 15456 10876 15484
rect 10781 15453 10793 15456
rect 10735 15447 10793 15453
rect 10870 15444 10876 15456
rect 10928 15444 10934 15496
rect 12069 15487 12127 15493
rect 12069 15453 12081 15487
rect 12115 15484 12127 15487
rect 12894 15484 12900 15496
rect 12115 15456 12900 15484
rect 12115 15453 12127 15456
rect 12069 15447 12127 15453
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 14461 15487 14519 15493
rect 14461 15453 14473 15487
rect 14507 15484 14519 15487
rect 14918 15484 14924 15496
rect 14507 15456 14924 15484
rect 14507 15453 14519 15456
rect 14461 15447 14519 15453
rect 14918 15444 14924 15456
rect 14976 15444 14982 15496
rect 15289 15487 15347 15493
rect 15289 15484 15301 15487
rect 15028 15456 15301 15484
rect 5521 15419 5580 15425
rect 5521 15385 5533 15419
rect 5567 15388 5580 15419
rect 5567 15385 5579 15388
rect 5521 15379 5579 15385
rect 5718 15376 5724 15428
rect 5776 15416 5782 15428
rect 6822 15416 6828 15428
rect 5776 15388 6828 15416
rect 5776 15376 5782 15388
rect 6822 15376 6828 15388
rect 6880 15376 6886 15428
rect 10505 15419 10563 15425
rect 10505 15385 10517 15419
rect 10551 15385 10563 15419
rect 10505 15379 10563 15385
rect 13081 15419 13139 15425
rect 13081 15385 13093 15419
rect 13127 15416 13139 15419
rect 14642 15416 14648 15428
rect 13127 15388 14648 15416
rect 13127 15385 13139 15388
rect 13081 15379 13139 15385
rect 1394 15308 1400 15360
rect 1452 15348 1458 15360
rect 1489 15351 1547 15357
rect 1489 15348 1501 15351
rect 1452 15320 1501 15348
rect 1452 15308 1458 15320
rect 1489 15317 1501 15320
rect 1535 15317 1547 15351
rect 1489 15311 1547 15317
rect 1762 15308 1768 15360
rect 1820 15348 1826 15360
rect 2225 15351 2283 15357
rect 2225 15348 2237 15351
rect 1820 15320 2237 15348
rect 1820 15308 1826 15320
rect 2225 15317 2237 15320
rect 2271 15317 2283 15351
rect 2225 15311 2283 15317
rect 2593 15351 2651 15357
rect 2593 15317 2605 15351
rect 2639 15348 2651 15351
rect 2682 15348 2688 15360
rect 2639 15320 2688 15348
rect 2639 15317 2651 15320
rect 2593 15311 2651 15317
rect 2682 15308 2688 15320
rect 2740 15308 2746 15360
rect 4798 15308 4804 15360
rect 4856 15308 4862 15360
rect 5626 15308 5632 15360
rect 5684 15348 5690 15360
rect 5997 15351 6055 15357
rect 5997 15348 6009 15351
rect 5684 15320 6009 15348
rect 5684 15308 5690 15320
rect 5997 15317 6009 15320
rect 6043 15317 6055 15351
rect 5997 15311 6055 15317
rect 6365 15351 6423 15357
rect 6365 15317 6377 15351
rect 6411 15348 6423 15351
rect 6730 15348 6736 15360
rect 6411 15320 6736 15348
rect 6411 15317 6423 15320
rect 6365 15311 6423 15317
rect 6730 15308 6736 15320
rect 6788 15308 6794 15360
rect 7926 15308 7932 15360
rect 7984 15348 7990 15360
rect 8389 15351 8447 15357
rect 8389 15348 8401 15351
rect 7984 15320 8401 15348
rect 7984 15308 7990 15320
rect 8389 15317 8401 15320
rect 8435 15348 8447 15351
rect 8846 15348 8852 15360
rect 8435 15320 8852 15348
rect 8435 15317 8447 15320
rect 8389 15311 8447 15317
rect 8846 15308 8852 15320
rect 8904 15308 8910 15360
rect 10410 15308 10416 15360
rect 10468 15348 10474 15360
rect 10520 15348 10548 15379
rect 14642 15376 14648 15388
rect 14700 15376 14706 15428
rect 14734 15376 14740 15428
rect 14792 15416 14798 15428
rect 15028 15416 15056 15456
rect 15289 15453 15301 15456
rect 15335 15484 15347 15487
rect 15378 15484 15384 15496
rect 15335 15456 15384 15484
rect 15335 15453 15347 15456
rect 15289 15447 15347 15453
rect 15378 15444 15384 15456
rect 15436 15444 15442 15496
rect 15470 15444 15476 15496
rect 15528 15444 15534 15496
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 16224 15481 16252 15524
rect 16301 15487 16359 15493
rect 16301 15481 16313 15487
rect 16224 15453 16313 15481
rect 16347 15453 16359 15487
rect 16301 15447 16359 15453
rect 16401 15487 16459 15493
rect 16401 15453 16413 15487
rect 16447 15484 16459 15487
rect 16500 15484 16528 15660
rect 16574 15648 16580 15660
rect 16632 15688 16638 15700
rect 17126 15688 17132 15700
rect 16632 15660 17132 15688
rect 16632 15648 16638 15660
rect 17126 15648 17132 15660
rect 17184 15648 17190 15700
rect 18782 15648 18788 15700
rect 18840 15688 18846 15700
rect 19337 15691 19395 15697
rect 19337 15688 19349 15691
rect 18840 15660 19349 15688
rect 18840 15648 18846 15660
rect 19337 15657 19349 15660
rect 19383 15657 19395 15691
rect 19337 15651 19395 15657
rect 20533 15691 20591 15697
rect 20533 15657 20545 15691
rect 20579 15688 20591 15691
rect 20622 15688 20628 15700
rect 20579 15660 20628 15688
rect 20579 15657 20591 15660
rect 20533 15651 20591 15657
rect 20622 15648 20628 15660
rect 20680 15648 20686 15700
rect 16758 15580 16764 15632
rect 16816 15580 16822 15632
rect 18598 15580 18604 15632
rect 18656 15580 18662 15632
rect 18690 15580 18696 15632
rect 18748 15620 18754 15632
rect 22462 15620 22468 15632
rect 18748 15592 22468 15620
rect 18748 15580 18754 15592
rect 22462 15580 22468 15592
rect 22520 15580 22526 15632
rect 19334 15512 19340 15564
rect 19392 15552 19398 15564
rect 20993 15555 21051 15561
rect 20993 15552 21005 15555
rect 19392 15524 21005 15552
rect 19392 15512 19398 15524
rect 20993 15521 21005 15524
rect 21039 15521 21051 15555
rect 20993 15515 21051 15521
rect 21174 15512 21180 15564
rect 21232 15552 21238 15564
rect 21726 15552 21732 15564
rect 21232 15524 21732 15552
rect 21232 15512 21238 15524
rect 21726 15512 21732 15524
rect 21784 15512 21790 15564
rect 23382 15512 23388 15564
rect 23440 15552 23446 15564
rect 24029 15555 24087 15561
rect 24029 15552 24041 15555
rect 23440 15524 24041 15552
rect 23440 15512 23446 15524
rect 24029 15521 24041 15524
rect 24075 15521 24087 15555
rect 24029 15515 24087 15521
rect 16447 15456 16528 15484
rect 16447 15453 16459 15456
rect 16401 15447 16459 15453
rect 16574 15444 16580 15496
rect 16632 15493 16638 15496
rect 16632 15487 16671 15493
rect 16659 15453 16671 15487
rect 16632 15447 16671 15453
rect 16761 15487 16819 15493
rect 16761 15453 16773 15487
rect 16807 15481 16819 15487
rect 16807 15453 16896 15481
rect 16761 15447 16819 15453
rect 16632 15444 16638 15447
rect 14792 15388 15056 15416
rect 16485 15419 16543 15425
rect 14792 15376 14798 15388
rect 16485 15385 16497 15419
rect 16531 15385 16543 15419
rect 16485 15379 16543 15385
rect 10468 15320 10548 15348
rect 10468 15308 10474 15320
rect 10870 15308 10876 15360
rect 10928 15308 10934 15360
rect 14826 15308 14832 15360
rect 14884 15308 14890 15360
rect 15013 15351 15071 15357
rect 15013 15317 15025 15351
rect 15059 15348 15071 15351
rect 15102 15348 15108 15360
rect 15059 15320 15108 15348
rect 15059 15317 15071 15320
rect 15013 15311 15071 15317
rect 15102 15308 15108 15320
rect 15160 15308 15166 15360
rect 16022 15308 16028 15360
rect 16080 15348 16086 15360
rect 16500 15348 16528 15379
rect 16080 15320 16528 15348
rect 16592 15348 16620 15444
rect 16868 15416 16896 15453
rect 17310 15444 17316 15496
rect 17368 15444 17374 15496
rect 18138 15444 18144 15496
rect 18196 15484 18202 15496
rect 18233 15487 18291 15493
rect 18233 15484 18245 15487
rect 18196 15456 18245 15484
rect 18196 15444 18202 15456
rect 18233 15453 18245 15456
rect 18279 15484 18291 15487
rect 19521 15487 19579 15493
rect 19521 15484 19533 15487
rect 18279 15456 19533 15484
rect 18279 15453 18291 15456
rect 18233 15447 18291 15453
rect 19521 15453 19533 15456
rect 19567 15453 19579 15487
rect 19521 15447 19579 15453
rect 19886 15444 19892 15496
rect 19944 15444 19950 15496
rect 20073 15487 20131 15493
rect 20073 15453 20085 15487
rect 20119 15453 20131 15487
rect 20073 15447 20131 15453
rect 20165 15487 20223 15493
rect 20165 15453 20177 15487
rect 20211 15453 20223 15487
rect 20165 15447 20223 15453
rect 20257 15487 20315 15493
rect 20257 15453 20269 15487
rect 20303 15484 20315 15487
rect 20898 15484 20904 15496
rect 20303 15456 20904 15484
rect 20303 15453 20315 15456
rect 20257 15447 20315 15453
rect 16942 15416 16948 15428
rect 16868 15388 16948 15416
rect 16942 15376 16948 15388
rect 17000 15416 17006 15428
rect 18966 15416 18972 15428
rect 17000 15388 18972 15416
rect 17000 15376 17006 15388
rect 18966 15376 18972 15388
rect 19024 15376 19030 15428
rect 19242 15376 19248 15428
rect 19300 15416 19306 15428
rect 20088 15416 20116 15447
rect 19300 15388 20116 15416
rect 19300 15376 19306 15388
rect 19518 15348 19524 15360
rect 16592 15320 19524 15348
rect 16080 15308 16086 15320
rect 19518 15308 19524 15320
rect 19576 15308 19582 15360
rect 19978 15308 19984 15360
rect 20036 15348 20042 15360
rect 20180 15348 20208 15447
rect 20898 15444 20904 15456
rect 20956 15444 20962 15496
rect 21450 15444 21456 15496
rect 21508 15444 21514 15496
rect 21634 15484 21640 15496
rect 21560 15456 21640 15484
rect 20622 15376 20628 15428
rect 20680 15416 20686 15428
rect 21560 15416 21588 15456
rect 21634 15444 21640 15456
rect 21692 15484 21698 15496
rect 21913 15487 21971 15493
rect 21913 15484 21925 15487
rect 21692 15456 21925 15484
rect 21692 15444 21698 15456
rect 21913 15453 21925 15456
rect 21959 15453 21971 15487
rect 21913 15447 21971 15453
rect 22094 15444 22100 15496
rect 22152 15484 22158 15496
rect 22741 15487 22799 15493
rect 22741 15484 22753 15487
rect 22152 15456 22753 15484
rect 22152 15444 22158 15456
rect 22741 15453 22753 15456
rect 22787 15484 22799 15487
rect 23198 15484 23204 15496
rect 22787 15456 23204 15484
rect 22787 15453 22799 15456
rect 22741 15447 22799 15453
rect 23198 15444 23204 15456
rect 23256 15444 23262 15496
rect 23474 15444 23480 15496
rect 23532 15444 23538 15496
rect 23566 15444 23572 15496
rect 23624 15484 23630 15496
rect 23661 15487 23719 15493
rect 23661 15484 23673 15487
rect 23624 15456 23673 15484
rect 23624 15444 23630 15456
rect 23661 15453 23673 15456
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 20680 15388 21588 15416
rect 21821 15419 21879 15425
rect 20680 15376 20686 15388
rect 21821 15385 21833 15419
rect 21867 15385 21879 15419
rect 21821 15379 21879 15385
rect 20036 15320 20208 15348
rect 20036 15308 20042 15320
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 21836 15348 21864 15379
rect 22002 15348 22008 15360
rect 20864 15320 22008 15348
rect 20864 15308 20870 15320
rect 22002 15308 22008 15320
rect 22060 15308 22066 15360
rect 23934 15308 23940 15360
rect 23992 15308 23998 15360
rect 1104 15258 24840 15280
rect 1104 15206 8214 15258
rect 8266 15206 8278 15258
rect 8330 15206 8342 15258
rect 8394 15206 8406 15258
rect 8458 15206 8470 15258
rect 8522 15206 16214 15258
rect 16266 15206 16278 15258
rect 16330 15206 16342 15258
rect 16394 15206 16406 15258
rect 16458 15206 16470 15258
rect 16522 15206 24214 15258
rect 24266 15206 24278 15258
rect 24330 15206 24342 15258
rect 24394 15206 24406 15258
rect 24458 15206 24470 15258
rect 24522 15206 24840 15258
rect 1104 15184 24840 15206
rect 2038 15104 2044 15156
rect 2096 15144 2102 15156
rect 2314 15144 2320 15156
rect 2372 15153 2378 15156
rect 2372 15147 2391 15153
rect 2096 15116 2320 15144
rect 2096 15104 2102 15116
rect 2314 15104 2320 15116
rect 2379 15113 2391 15147
rect 4062 15144 4068 15156
rect 2372 15107 2391 15113
rect 2976 15116 4068 15144
rect 2372 15104 2378 15107
rect 2130 15036 2136 15088
rect 2188 15036 2194 15088
rect 2976 15020 3004 15116
rect 4062 15104 4068 15116
rect 4120 15104 4126 15156
rect 4709 15147 4767 15153
rect 4709 15113 4721 15147
rect 4755 15144 4767 15147
rect 4798 15144 4804 15156
rect 4755 15116 4804 15144
rect 4755 15113 4767 15116
rect 4709 15107 4767 15113
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 5166 15104 5172 15156
rect 5224 15144 5230 15156
rect 5224 15116 8708 15144
rect 5224 15104 5230 15116
rect 3970 15036 3976 15088
rect 4028 15036 4034 15088
rect 5629 15079 5687 15085
rect 5629 15045 5641 15079
rect 5675 15045 5687 15079
rect 5629 15039 5687 15045
rect 5845 15079 5903 15085
rect 5845 15045 5857 15079
rect 5891 15076 5903 15079
rect 5994 15076 6000 15088
rect 5891 15048 6000 15076
rect 5891 15045 5903 15048
rect 5845 15039 5903 15045
rect 1394 14968 1400 15020
rect 1452 15008 1458 15020
rect 1489 15011 1547 15017
rect 1489 15008 1501 15011
rect 1452 14980 1501 15008
rect 1452 14968 1458 14980
rect 1489 14977 1501 14980
rect 1535 14977 1547 15011
rect 1489 14971 1547 14977
rect 2958 14968 2964 15020
rect 3016 14968 3022 15020
rect 5644 15008 5672 15039
rect 5994 15036 6000 15048
rect 6052 15036 6058 15088
rect 7650 15036 7656 15088
rect 7708 15076 7714 15088
rect 7708 15048 7866 15076
rect 7708 15036 7714 15048
rect 7006 15008 7012 15020
rect 5644 14980 7012 15008
rect 7006 14968 7012 14980
rect 7064 14968 7070 15020
rect 7098 14968 7104 15020
rect 7156 14968 7162 15020
rect 8680 15008 8708 15116
rect 8846 15104 8852 15156
rect 8904 15104 8910 15156
rect 10226 15104 10232 15156
rect 10284 15144 10290 15156
rect 10413 15147 10471 15153
rect 10413 15144 10425 15147
rect 10284 15116 10425 15144
rect 10284 15104 10290 15116
rect 10413 15113 10425 15116
rect 10459 15113 10471 15147
rect 10413 15107 10471 15113
rect 11977 15147 12035 15153
rect 11977 15113 11989 15147
rect 12023 15113 12035 15147
rect 11977 15107 12035 15113
rect 10594 15076 10600 15088
rect 9876 15048 10600 15076
rect 9876 15020 9904 15048
rect 10594 15036 10600 15048
rect 10652 15076 10658 15088
rect 11698 15076 11704 15088
rect 10652 15048 11704 15076
rect 10652 15036 10658 15048
rect 11698 15036 11704 15048
rect 11756 15076 11762 15088
rect 11992 15076 12020 15107
rect 13078 15104 13084 15156
rect 13136 15144 13142 15156
rect 13173 15147 13231 15153
rect 13173 15144 13185 15147
rect 13136 15116 13185 15144
rect 13136 15104 13142 15116
rect 13173 15113 13185 15116
rect 13219 15113 13231 15147
rect 13173 15107 13231 15113
rect 14001 15147 14059 15153
rect 14001 15113 14013 15147
rect 14047 15144 14059 15147
rect 14461 15147 14519 15153
rect 14461 15144 14473 15147
rect 14047 15116 14473 15144
rect 14047 15113 14059 15116
rect 14001 15107 14059 15113
rect 14461 15113 14473 15116
rect 14507 15113 14519 15147
rect 15010 15144 15016 15156
rect 14461 15107 14519 15113
rect 14936 15116 15016 15144
rect 12897 15079 12955 15085
rect 11756 15048 12572 15076
rect 11756 15036 11762 15048
rect 9769 15011 9827 15017
rect 9769 15008 9781 15011
rect 8680 14980 9781 15008
rect 9769 14977 9781 14980
rect 9815 14977 9827 15011
rect 9769 14971 9827 14977
rect 9858 14968 9864 15020
rect 9916 14968 9922 15020
rect 10045 15011 10103 15017
rect 10045 14977 10057 15011
rect 10091 14977 10103 15011
rect 10045 14971 10103 14977
rect 3237 14943 3295 14949
rect 3237 14909 3249 14943
rect 3283 14940 3295 14943
rect 3878 14940 3884 14952
rect 3283 14912 3884 14940
rect 3283 14909 3295 14912
rect 3237 14903 3295 14909
rect 3878 14900 3884 14912
rect 3936 14900 3942 14952
rect 7377 14943 7435 14949
rect 7377 14909 7389 14943
rect 7423 14940 7435 14943
rect 7834 14940 7840 14952
rect 7423 14912 7840 14940
rect 7423 14909 7435 14912
rect 7377 14903 7435 14909
rect 7834 14900 7840 14912
rect 7892 14900 7898 14952
rect 10060 14940 10088 14971
rect 10134 14968 10140 15020
rect 10192 14968 10198 15020
rect 10689 15011 10747 15017
rect 10689 14977 10701 15011
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 11149 15011 11207 15017
rect 11149 14977 11161 15011
rect 11195 15008 11207 15011
rect 11330 15008 11336 15020
rect 11195 14980 11336 15008
rect 11195 14977 11207 14980
rect 11149 14971 11207 14977
rect 10410 14940 10416 14952
rect 10060 14912 10416 14940
rect 10410 14900 10416 14912
rect 10468 14940 10474 14952
rect 10704 14940 10732 14971
rect 11330 14968 11336 14980
rect 11388 14968 11394 15020
rect 11606 14968 11612 15020
rect 11664 14968 11670 15020
rect 11790 14968 11796 15020
rect 11848 14968 11854 15020
rect 11974 14968 11980 15020
rect 12032 15008 12038 15020
rect 12544 15017 12572 15048
rect 12897 15045 12909 15079
rect 12943 15076 12955 15079
rect 13722 15076 13728 15088
rect 12943 15048 13728 15076
rect 12943 15045 12955 15048
rect 12897 15039 12955 15045
rect 13722 15036 13728 15048
rect 13780 15076 13786 15088
rect 14016 15076 14044 15107
rect 14734 15076 14740 15088
rect 13780 15048 14044 15076
rect 14200 15048 14740 15076
rect 13780 15036 13786 15048
rect 12710 15017 12716 15020
rect 12069 15011 12127 15017
rect 12069 15008 12081 15011
rect 12032 14980 12081 15008
rect 12032 14968 12038 14980
rect 12069 14977 12081 14980
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 12529 15011 12587 15017
rect 12529 14977 12541 15011
rect 12575 14977 12587 15011
rect 12529 14971 12587 14977
rect 12687 15011 12716 15017
rect 12687 14977 12699 15011
rect 12687 14971 12716 14977
rect 12710 14968 12716 14971
rect 12768 14968 12774 15020
rect 12802 14968 12808 15020
rect 12860 14968 12866 15020
rect 12989 15011 13047 15017
rect 12989 14977 13001 15011
rect 13035 15008 13047 15011
rect 13262 15008 13268 15020
rect 13035 14980 13268 15008
rect 13035 14977 13047 14980
rect 12989 14971 13047 14977
rect 13262 14968 13268 14980
rect 13320 14968 13326 15020
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13633 15011 13691 15017
rect 13633 15008 13645 15011
rect 13412 14980 13645 15008
rect 13412 14968 13418 14980
rect 13633 14977 13645 14980
rect 13679 14977 13691 15011
rect 13633 14971 13691 14977
rect 13814 14968 13820 15020
rect 13872 15017 13878 15020
rect 14200 15017 14228 15048
rect 14734 15036 14740 15048
rect 14792 15036 14798 15088
rect 13872 15011 13921 15017
rect 13872 14977 13875 15011
rect 13909 14977 13921 15011
rect 13872 14971 13921 14977
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14829 15011 14887 15017
rect 14829 14977 14841 15011
rect 14875 15008 14887 15011
rect 14936 15008 14964 15116
rect 15010 15104 15016 15116
rect 15068 15144 15074 15156
rect 15654 15144 15660 15156
rect 15068 15116 15660 15144
rect 15068 15104 15074 15116
rect 15654 15104 15660 15116
rect 15712 15104 15718 15156
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 16022 15144 16028 15156
rect 15795 15116 16028 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16022 15104 16028 15116
rect 16080 15104 16086 15156
rect 16393 15147 16451 15153
rect 16393 15113 16405 15147
rect 16439 15144 16451 15147
rect 16942 15144 16948 15156
rect 16439 15116 16948 15144
rect 16439 15113 16451 15116
rect 16393 15107 16451 15113
rect 16942 15104 16948 15116
rect 17000 15104 17006 15156
rect 17310 15104 17316 15156
rect 17368 15104 17374 15156
rect 18782 15144 18788 15156
rect 17420 15116 18788 15144
rect 15473 15079 15531 15085
rect 15473 15045 15485 15079
rect 15519 15076 15531 15079
rect 15562 15076 15568 15088
rect 15519 15048 15568 15076
rect 15519 15045 15531 15048
rect 15473 15039 15531 15045
rect 15562 15036 15568 15048
rect 15620 15036 15626 15088
rect 17420 15076 17448 15116
rect 18782 15104 18788 15116
rect 18840 15144 18846 15156
rect 19242 15144 19248 15156
rect 18840 15116 19248 15144
rect 18840 15104 18846 15116
rect 19242 15104 19248 15116
rect 19300 15104 19306 15156
rect 19426 15104 19432 15156
rect 19484 15104 19490 15156
rect 19702 15104 19708 15156
rect 19760 15144 19766 15156
rect 19760 15116 20300 15144
rect 19760 15104 19766 15116
rect 16224 15048 17448 15076
rect 14875 14980 14964 15008
rect 15105 15011 15163 15017
rect 14875 14977 14887 14980
rect 14829 14971 14887 14977
rect 15105 14977 15117 15011
rect 15151 15008 15163 15011
rect 15286 15008 15292 15020
rect 15151 14980 15292 15008
rect 15151 14977 15163 14980
rect 15105 14971 15163 14977
rect 13872 14968 13878 14971
rect 15286 14968 15292 14980
rect 15344 14968 15350 15020
rect 15488 14980 16068 15008
rect 11808 14940 11836 14968
rect 10468 14912 11836 14940
rect 13280 14940 13308 14968
rect 15488 14952 15516 14980
rect 14093 14943 14151 14949
rect 14093 14940 14105 14943
rect 13280 14912 14105 14940
rect 10468 14900 10474 14912
rect 14093 14909 14105 14912
rect 14139 14909 14151 14943
rect 14093 14903 14151 14909
rect 14642 14900 14648 14952
rect 14700 14940 14706 14952
rect 14737 14943 14795 14949
rect 14737 14940 14749 14943
rect 14700 14912 14749 14940
rect 14700 14900 14706 14912
rect 14737 14909 14749 14912
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 14918 14900 14924 14952
rect 14976 14940 14982 14952
rect 15381 14943 15439 14949
rect 15381 14940 15393 14943
rect 14976 14912 15393 14940
rect 14976 14900 14982 14912
rect 15381 14909 15393 14912
rect 15427 14909 15439 14943
rect 15381 14903 15439 14909
rect 15470 14900 15476 14952
rect 15528 14900 15534 14952
rect 15590 14943 15648 14949
rect 15590 14909 15602 14943
rect 15636 14940 15648 14943
rect 15838 14940 15844 14952
rect 15636 14912 15844 14940
rect 15636 14909 15648 14912
rect 15590 14903 15648 14909
rect 15838 14900 15844 14912
rect 15896 14900 15902 14952
rect 16040 14940 16068 14980
rect 16114 14968 16120 15020
rect 16172 14968 16178 15020
rect 16224 15017 16252 15048
rect 18138 15036 18144 15088
rect 18196 15076 18202 15088
rect 18233 15079 18291 15085
rect 18233 15076 18245 15079
rect 18196 15048 18245 15076
rect 18196 15036 18202 15048
rect 18233 15045 18245 15048
rect 18279 15045 18291 15079
rect 18233 15039 18291 15045
rect 18414 15036 18420 15088
rect 18472 15036 18478 15088
rect 16209 15011 16267 15017
rect 16209 14977 16221 15011
rect 16255 14977 16267 15011
rect 16209 14971 16267 14977
rect 16761 15011 16819 15017
rect 16761 14977 16773 15011
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 16945 15011 17003 15017
rect 16945 14977 16957 15011
rect 16991 14977 17003 15011
rect 16945 14971 17003 14977
rect 16776 14940 16804 14971
rect 16040 14912 16804 14940
rect 16960 14940 16988 14971
rect 17034 14968 17040 15020
rect 17092 14968 17098 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 15008 17187 15011
rect 17218 15008 17224 15020
rect 17175 14980 17224 15008
rect 17175 14977 17187 14980
rect 17129 14971 17187 14977
rect 17218 14968 17224 14980
rect 17276 14968 17282 15020
rect 17773 15011 17831 15017
rect 17773 14977 17785 15011
rect 17819 15008 17831 15011
rect 19153 15011 19211 15017
rect 17819 14980 17908 15008
rect 17819 14977 17831 14980
rect 17773 14971 17831 14977
rect 17310 14940 17316 14952
rect 16960 14912 17316 14940
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 1673 14875 1731 14881
rect 1673 14841 1685 14875
rect 1719 14872 1731 14875
rect 9585 14875 9643 14881
rect 1719 14844 2774 14872
rect 1719 14841 1731 14844
rect 1673 14835 1731 14841
rect 1946 14764 1952 14816
rect 2004 14804 2010 14816
rect 2317 14807 2375 14813
rect 2317 14804 2329 14807
rect 2004 14776 2329 14804
rect 2004 14764 2010 14776
rect 2317 14773 2329 14776
rect 2363 14773 2375 14807
rect 2317 14767 2375 14773
rect 2498 14764 2504 14816
rect 2556 14764 2562 14816
rect 2746 14804 2774 14844
rect 4264 14844 6684 14872
rect 4264 14804 4292 14844
rect 2746 14776 4292 14804
rect 5810 14764 5816 14816
rect 5868 14764 5874 14816
rect 5994 14764 6000 14816
rect 6052 14764 6058 14816
rect 6656 14804 6684 14844
rect 9585 14841 9597 14875
rect 9631 14872 9643 14875
rect 10594 14872 10600 14884
rect 9631 14844 10600 14872
rect 9631 14841 9643 14844
rect 9585 14835 9643 14841
rect 10594 14832 10600 14844
rect 10652 14832 10658 14884
rect 10873 14875 10931 14881
rect 10873 14841 10885 14875
rect 10919 14872 10931 14875
rect 11146 14872 11152 14884
rect 10919 14844 11152 14872
rect 10919 14841 10931 14844
rect 10873 14835 10931 14841
rect 11146 14832 11152 14844
rect 11204 14832 11210 14884
rect 17770 14872 17776 14884
rect 14660 14844 17776 14872
rect 10502 14804 10508 14816
rect 6656 14776 10508 14804
rect 10502 14764 10508 14776
rect 10560 14764 10566 14816
rect 10778 14764 10784 14816
rect 10836 14764 10842 14816
rect 10962 14764 10968 14816
rect 11020 14764 11026 14816
rect 13633 14807 13691 14813
rect 13633 14773 13645 14807
rect 13679 14804 13691 14807
rect 14660 14804 14688 14844
rect 17770 14832 17776 14844
rect 17828 14832 17834 14884
rect 13679 14776 14688 14804
rect 14829 14807 14887 14813
rect 13679 14773 13691 14776
rect 13633 14767 13691 14773
rect 14829 14773 14841 14807
rect 14875 14804 14887 14807
rect 15010 14804 15016 14816
rect 14875 14776 15016 14804
rect 14875 14773 14887 14776
rect 14829 14767 14887 14773
rect 15010 14764 15016 14776
rect 15068 14804 15074 14816
rect 15194 14804 15200 14816
rect 15068 14776 15200 14804
rect 15068 14764 15074 14776
rect 15194 14764 15200 14776
rect 15252 14804 15258 14816
rect 17034 14804 17040 14816
rect 15252 14776 17040 14804
rect 15252 14764 15258 14776
rect 17034 14764 17040 14776
rect 17092 14764 17098 14816
rect 17586 14764 17592 14816
rect 17644 14804 17650 14816
rect 17880 14804 17908 14980
rect 19153 14977 19165 15011
rect 19199 15008 19211 15011
rect 19334 15008 19340 15020
rect 19199 14980 19340 15008
rect 19199 14977 19211 14980
rect 19153 14971 19211 14977
rect 19334 14968 19340 14980
rect 19392 14968 19398 15020
rect 19610 14968 19616 15020
rect 19668 14968 19674 15020
rect 19886 14968 19892 15020
rect 19944 15008 19950 15020
rect 20272 15017 20300 15116
rect 20622 15104 20628 15156
rect 20680 15104 20686 15156
rect 20717 15147 20775 15153
rect 20717 15113 20729 15147
rect 20763 15144 20775 15147
rect 21545 15147 21603 15153
rect 20763 15116 21496 15144
rect 20763 15113 20775 15116
rect 20717 15107 20775 15113
rect 20640 15076 20668 15104
rect 20364 15048 20668 15076
rect 20364 15017 20392 15048
rect 20898 15036 20904 15088
rect 20956 15076 20962 15088
rect 20956 15048 21404 15076
rect 20956 15036 20962 15048
rect 20073 15011 20131 15017
rect 20073 15008 20085 15011
rect 19944 14980 20085 15008
rect 19944 14968 19950 14980
rect 20073 14977 20085 14980
rect 20119 14977 20131 15011
rect 20073 14971 20131 14977
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20257 14971 20315 14977
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 14977 20407 15011
rect 20349 14971 20407 14977
rect 20441 15011 20499 15017
rect 20441 14977 20453 15011
rect 20487 15008 20499 15011
rect 20622 15008 20628 15020
rect 20487 14980 20628 15008
rect 20487 14977 20499 14980
rect 20441 14971 20499 14977
rect 20622 14968 20628 14980
rect 20680 14968 20686 15020
rect 20990 14968 20996 15020
rect 21048 14968 21054 15020
rect 21174 14968 21180 15020
rect 21232 14968 21238 15020
rect 21266 14968 21272 15020
rect 21324 14968 21330 15020
rect 21376 15017 21404 15048
rect 21361 15011 21419 15017
rect 21361 14977 21373 15011
rect 21407 14977 21419 15011
rect 21468 15008 21496 15116
rect 21545 15113 21557 15147
rect 21591 15144 21603 15147
rect 22094 15144 22100 15156
rect 21591 15116 22100 15144
rect 21591 15113 21603 15116
rect 21545 15107 21603 15113
rect 22094 15104 22100 15116
rect 22152 15104 22158 15156
rect 22186 15104 22192 15156
rect 22244 15144 22250 15156
rect 22557 15147 22615 15153
rect 22557 15144 22569 15147
rect 22244 15116 22569 15144
rect 22244 15104 22250 15116
rect 22557 15113 22569 15116
rect 22603 15113 22615 15147
rect 22557 15107 22615 15113
rect 21726 15036 21732 15088
rect 21784 15076 21790 15088
rect 21784 15048 22048 15076
rect 21784 15036 21790 15048
rect 21542 15008 21548 15020
rect 21468 14980 21548 15008
rect 21361 14971 21419 14977
rect 21542 14968 21548 14980
rect 21600 15008 21606 15020
rect 22020 15017 22048 15048
rect 23382 15036 23388 15088
rect 23440 15036 23446 15088
rect 23566 15036 23572 15088
rect 23624 15076 23630 15088
rect 23661 15079 23719 15085
rect 23661 15076 23673 15079
rect 23624 15048 23673 15076
rect 23624 15036 23630 15048
rect 23661 15045 23673 15048
rect 23707 15045 23719 15079
rect 23661 15039 23719 15045
rect 21913 15011 21971 15017
rect 21913 15008 21925 15011
rect 21600 14980 21925 15008
rect 21600 14968 21606 14980
rect 21913 14977 21925 14980
rect 21959 14977 21971 15011
rect 21913 14971 21971 14977
rect 22006 15011 22064 15017
rect 22006 14977 22018 15011
rect 22052 14977 22064 15011
rect 22006 14971 22064 14977
rect 22094 14968 22100 15020
rect 22152 15008 22158 15020
rect 22189 15011 22247 15017
rect 22189 15008 22201 15011
rect 22152 14980 22201 15008
rect 22152 14968 22158 14980
rect 22189 14977 22201 14980
rect 22235 14977 22247 15011
rect 22189 14971 22247 14977
rect 22278 14968 22284 15020
rect 22336 14968 22342 15020
rect 22370 14968 22376 15020
rect 22428 15017 22434 15020
rect 22428 15008 22436 15017
rect 23293 15011 23351 15017
rect 22428 14980 22473 15008
rect 22428 14971 22436 14980
rect 23293 14977 23305 15011
rect 23339 15008 23351 15011
rect 23750 15008 23756 15020
rect 23339 14980 23756 15008
rect 23339 14977 23351 14980
rect 23293 14971 23351 14977
rect 22428 14968 22434 14971
rect 23750 14968 23756 14980
rect 23808 15008 23814 15020
rect 23845 15011 23903 15017
rect 23845 15008 23857 15011
rect 23808 14980 23857 15008
rect 23808 14968 23814 14980
rect 23845 14977 23857 14980
rect 23891 14977 23903 15011
rect 23845 14971 23903 14977
rect 24118 14968 24124 15020
rect 24176 15008 24182 15020
rect 24397 15011 24455 15017
rect 24397 15008 24409 15011
rect 24176 14980 24409 15008
rect 24176 14968 24182 14980
rect 24397 14977 24409 14980
rect 24443 14977 24455 15011
rect 24397 14971 24455 14977
rect 22462 14940 22468 14952
rect 17972 14912 22468 14940
rect 17972 14881 18000 14912
rect 22462 14900 22468 14912
rect 22520 14900 22526 14952
rect 22833 14943 22891 14949
rect 22833 14909 22845 14943
rect 22879 14909 22891 14943
rect 22833 14903 22891 14909
rect 17957 14875 18015 14881
rect 17957 14841 17969 14875
rect 18003 14841 18015 14875
rect 17957 14835 18015 14841
rect 18046 14832 18052 14884
rect 18104 14872 18110 14884
rect 22278 14872 22284 14884
rect 18104 14844 22284 14872
rect 18104 14832 18110 14844
rect 22278 14832 22284 14844
rect 22336 14872 22342 14884
rect 22848 14872 22876 14903
rect 25038 14872 25044 14884
rect 22336 14844 22876 14872
rect 22940 14844 25044 14872
rect 22336 14832 22342 14844
rect 22940 14804 22968 14844
rect 25038 14832 25044 14844
rect 25096 14832 25102 14884
rect 17644 14776 22968 14804
rect 17644 14764 17650 14776
rect 23014 14764 23020 14816
rect 23072 14804 23078 14816
rect 24213 14807 24271 14813
rect 24213 14804 24225 14807
rect 23072 14776 24225 14804
rect 23072 14764 23078 14776
rect 24213 14773 24225 14776
rect 24259 14773 24271 14807
rect 24213 14767 24271 14773
rect 1104 14714 24840 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 12214 14714
rect 12266 14662 12278 14714
rect 12330 14662 12342 14714
rect 12394 14662 12406 14714
rect 12458 14662 12470 14714
rect 12522 14662 20214 14714
rect 20266 14662 20278 14714
rect 20330 14662 20342 14714
rect 20394 14662 20406 14714
rect 20458 14662 20470 14714
rect 20522 14662 24840 14714
rect 1104 14640 24840 14662
rect 3878 14560 3884 14612
rect 3936 14560 3942 14612
rect 7377 14603 7435 14609
rect 7377 14569 7389 14603
rect 7423 14600 7435 14603
rect 7561 14603 7619 14609
rect 7423 14572 7512 14600
rect 7423 14569 7435 14572
rect 7377 14563 7435 14569
rect 4062 14492 4068 14544
rect 4120 14532 4126 14544
rect 7484 14532 7512 14572
rect 7561 14569 7573 14603
rect 7607 14600 7619 14603
rect 7650 14600 7656 14612
rect 7607 14572 7656 14600
rect 7607 14569 7619 14572
rect 7561 14563 7619 14569
rect 7650 14560 7656 14572
rect 7708 14560 7714 14612
rect 7834 14560 7840 14612
rect 7892 14560 7898 14612
rect 8662 14600 8668 14612
rect 7944 14572 8668 14600
rect 7944 14532 7972 14572
rect 8662 14560 8668 14572
rect 8720 14600 8726 14612
rect 9306 14600 9312 14612
rect 8720 14572 9312 14600
rect 8720 14560 8726 14572
rect 9306 14560 9312 14572
rect 9364 14560 9370 14612
rect 9861 14603 9919 14609
rect 9861 14569 9873 14603
rect 9907 14600 9919 14603
rect 9950 14600 9956 14612
rect 9907 14572 9956 14600
rect 9907 14569 9919 14572
rect 9861 14563 9919 14569
rect 9950 14560 9956 14572
rect 10008 14560 10014 14612
rect 11701 14603 11759 14609
rect 11701 14569 11713 14603
rect 11747 14600 11759 14603
rect 11790 14600 11796 14612
rect 11747 14572 11796 14600
rect 11747 14569 11759 14572
rect 11701 14563 11759 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 12621 14603 12679 14609
rect 12621 14569 12633 14603
rect 12667 14600 12679 14603
rect 12802 14600 12808 14612
rect 12667 14572 12808 14600
rect 12667 14569 12679 14572
rect 12621 14563 12679 14569
rect 12802 14560 12808 14572
rect 12860 14560 12866 14612
rect 13262 14560 13268 14612
rect 13320 14600 13326 14612
rect 15470 14600 15476 14612
rect 13320 14572 15476 14600
rect 13320 14560 13326 14572
rect 15470 14560 15476 14572
rect 15528 14560 15534 14612
rect 16942 14560 16948 14612
rect 17000 14560 17006 14612
rect 17310 14560 17316 14612
rect 17368 14560 17374 14612
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19610 14600 19616 14612
rect 19392 14572 19616 14600
rect 19392 14560 19398 14572
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 21082 14560 21088 14612
rect 21140 14560 21146 14612
rect 21358 14560 21364 14612
rect 21416 14600 21422 14612
rect 21545 14603 21603 14609
rect 21545 14600 21557 14603
rect 21416 14572 21557 14600
rect 21416 14560 21422 14572
rect 21545 14569 21557 14572
rect 21591 14569 21603 14603
rect 21545 14563 21603 14569
rect 4120 14504 5028 14532
rect 7484 14504 7972 14532
rect 4120 14492 4126 14504
rect 1486 14424 1492 14476
rect 1544 14464 1550 14476
rect 2958 14464 2964 14476
rect 1544 14436 2964 14464
rect 1544 14424 1550 14436
rect 2958 14424 2964 14436
rect 3016 14424 3022 14476
rect 4525 14467 4583 14473
rect 4525 14433 4537 14467
rect 4571 14464 4583 14467
rect 4890 14464 4896 14476
rect 4571 14436 4896 14464
rect 4571 14433 4583 14436
rect 4525 14427 4583 14433
rect 4890 14424 4896 14436
rect 4948 14424 4954 14476
rect 5000 14473 5028 14504
rect 10962 14492 10968 14544
rect 11020 14532 11026 14544
rect 11057 14535 11115 14541
rect 11057 14532 11069 14535
rect 11020 14504 11069 14532
rect 11020 14492 11026 14504
rect 11057 14501 11069 14504
rect 11103 14532 11115 14535
rect 11882 14532 11888 14544
rect 11103 14504 11888 14532
rect 11103 14501 11115 14504
rect 11057 14495 11115 14501
rect 11882 14492 11888 14504
rect 11940 14532 11946 14544
rect 11977 14535 12035 14541
rect 11977 14532 11989 14535
rect 11940 14504 11989 14532
rect 11940 14492 11946 14504
rect 11977 14501 11989 14504
rect 12023 14501 12035 14535
rect 11977 14495 12035 14501
rect 12066 14492 12072 14544
rect 12124 14492 12130 14544
rect 12894 14492 12900 14544
rect 12952 14532 12958 14544
rect 13538 14532 13544 14544
rect 12952 14504 13544 14532
rect 12952 14492 12958 14504
rect 13538 14492 13544 14504
rect 13596 14532 13602 14544
rect 16025 14535 16083 14541
rect 13596 14504 14964 14532
rect 13596 14492 13602 14504
rect 4985 14467 5043 14473
rect 4985 14433 4997 14467
rect 5031 14464 5043 14467
rect 7098 14464 7104 14476
rect 5031 14436 7104 14464
rect 5031 14433 5043 14436
rect 4985 14427 5043 14433
rect 7098 14424 7104 14436
rect 7156 14424 7162 14476
rect 7926 14424 7932 14476
rect 7984 14464 7990 14476
rect 8389 14467 8447 14473
rect 7984 14436 8248 14464
rect 7984 14424 7990 14436
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4798 14396 4804 14408
rect 4295 14368 4804 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 4798 14356 4804 14368
rect 4856 14356 4862 14408
rect 8220 14405 8248 14436
rect 8389 14433 8401 14467
rect 8435 14464 8447 14467
rect 8435 14436 8524 14464
rect 8435 14433 8447 14436
rect 8389 14427 8447 14433
rect 8205 14399 8263 14405
rect 8205 14365 8217 14399
rect 8251 14365 8263 14399
rect 8496 14396 8524 14436
rect 9122 14424 9128 14476
rect 9180 14464 9186 14476
rect 12084 14464 12112 14492
rect 9180 14436 12020 14464
rect 12084 14436 12204 14464
rect 9180 14424 9186 14436
rect 8570 14396 8576 14408
rect 8496 14368 8576 14396
rect 8205 14359 8263 14365
rect 8570 14356 8576 14368
rect 8628 14356 8634 14408
rect 9766 14356 9772 14408
rect 9824 14396 9830 14408
rect 9993 14399 10051 14405
rect 9993 14396 10005 14399
rect 9824 14368 10005 14396
rect 9824 14356 9830 14368
rect 9993 14365 10005 14368
rect 10039 14365 10051 14399
rect 9993 14359 10051 14365
rect 10410 14356 10416 14408
rect 10468 14356 10474 14408
rect 10778 14356 10784 14408
rect 10836 14396 10842 14408
rect 10965 14399 11023 14405
rect 10965 14396 10977 14399
rect 10836 14368 10977 14396
rect 10836 14356 10842 14368
rect 10965 14365 10977 14368
rect 11011 14365 11023 14399
rect 10965 14359 11023 14365
rect 11149 14399 11207 14405
rect 11149 14365 11161 14399
rect 11195 14365 11207 14399
rect 11149 14359 11207 14365
rect 1762 14288 1768 14340
rect 1820 14288 1826 14340
rect 2498 14288 2504 14340
rect 2556 14288 2562 14340
rect 5261 14331 5319 14337
rect 5261 14297 5273 14331
rect 5307 14328 5319 14331
rect 5534 14328 5540 14340
rect 5307 14300 5540 14328
rect 5307 14297 5319 14300
rect 5261 14291 5319 14297
rect 5534 14288 5540 14300
rect 5592 14288 5598 14340
rect 5994 14288 6000 14340
rect 6052 14288 6058 14340
rect 7006 14288 7012 14340
rect 7064 14328 7070 14340
rect 7193 14331 7251 14337
rect 7193 14328 7205 14331
rect 7064 14300 7205 14328
rect 7064 14288 7070 14300
rect 7193 14297 7205 14300
rect 7239 14328 7251 14331
rect 8018 14328 8024 14340
rect 7239 14300 8024 14328
rect 7239 14297 7251 14300
rect 7193 14291 7251 14297
rect 8018 14288 8024 14300
rect 8076 14288 8082 14340
rect 8110 14288 8116 14340
rect 8168 14328 8174 14340
rect 8297 14331 8355 14337
rect 8297 14328 8309 14331
rect 8168 14300 8309 14328
rect 8168 14288 8174 14300
rect 8297 14297 8309 14300
rect 8343 14297 8355 14331
rect 9214 14328 9220 14340
rect 8297 14291 8355 14297
rect 8772 14300 9220 14328
rect 8772 14272 8800 14300
rect 9214 14288 9220 14300
rect 9272 14337 9278 14340
rect 9272 14331 9335 14337
rect 9272 14297 9289 14331
rect 9323 14297 9335 14331
rect 9272 14291 9335 14297
rect 9493 14331 9551 14337
rect 9493 14297 9505 14331
rect 9539 14297 9551 14331
rect 9493 14291 9551 14297
rect 9272 14288 9278 14291
rect 2682 14220 2688 14272
rect 2740 14260 2746 14272
rect 3237 14263 3295 14269
rect 3237 14260 3249 14263
rect 2740 14232 3249 14260
rect 2740 14220 2746 14232
rect 3237 14229 3249 14232
rect 3283 14229 3295 14263
rect 3237 14223 3295 14229
rect 3326 14220 3332 14272
rect 3384 14260 3390 14272
rect 4341 14263 4399 14269
rect 4341 14260 4353 14263
rect 3384 14232 4353 14260
rect 3384 14220 3390 14232
rect 4341 14229 4353 14232
rect 4387 14229 4399 14263
rect 4341 14223 4399 14229
rect 6730 14220 6736 14272
rect 6788 14220 6794 14272
rect 6914 14220 6920 14272
rect 6972 14260 6978 14272
rect 7403 14263 7461 14269
rect 7403 14260 7415 14263
rect 6972 14232 7415 14260
rect 6972 14220 6978 14232
rect 7403 14229 7415 14232
rect 7449 14260 7461 14263
rect 8754 14260 8760 14272
rect 7449 14232 8760 14260
rect 7449 14229 7461 14232
rect 7403 14223 7461 14229
rect 8754 14220 8760 14232
rect 8812 14220 8818 14272
rect 9030 14220 9036 14272
rect 9088 14260 9094 14272
rect 9125 14263 9183 14269
rect 9125 14260 9137 14263
rect 9088 14232 9137 14260
rect 9088 14220 9094 14232
rect 9125 14229 9137 14232
rect 9171 14229 9183 14263
rect 9508 14260 9536 14291
rect 9858 14288 9864 14340
rect 9916 14328 9922 14340
rect 10137 14331 10195 14337
rect 10137 14328 10149 14331
rect 9916 14300 10149 14328
rect 9916 14288 9922 14300
rect 10137 14297 10149 14300
rect 10183 14297 10195 14331
rect 10137 14291 10195 14297
rect 10229 14331 10287 14337
rect 10229 14297 10241 14331
rect 10275 14328 10287 14331
rect 10689 14331 10747 14337
rect 10689 14328 10701 14331
rect 10275 14300 10701 14328
rect 10275 14297 10287 14300
rect 10229 14291 10287 14297
rect 10689 14297 10701 14300
rect 10735 14297 10747 14331
rect 11164 14328 11192 14359
rect 11238 14356 11244 14408
rect 11296 14356 11302 14408
rect 11422 14356 11428 14408
rect 11480 14356 11486 14408
rect 11790 14356 11796 14408
rect 11848 14398 11854 14408
rect 11885 14399 11943 14405
rect 11885 14398 11897 14399
rect 11848 14370 11897 14398
rect 11848 14356 11854 14370
rect 11885 14365 11897 14370
rect 11931 14365 11943 14399
rect 11885 14359 11943 14365
rect 11330 14328 11336 14340
rect 11164 14300 11336 14328
rect 10689 14291 10747 14297
rect 11330 14288 11336 14300
rect 11388 14328 11394 14340
rect 11808 14328 11836 14356
rect 11388 14300 11836 14328
rect 11992 14328 12020 14436
rect 12066 14356 12072 14408
rect 12124 14356 12130 14408
rect 12176 14405 12204 14436
rect 12268 14436 13032 14464
rect 12161 14399 12219 14405
rect 12161 14365 12173 14399
rect 12207 14365 12219 14399
rect 12161 14359 12219 14365
rect 12268 14328 12296 14436
rect 12529 14399 12587 14405
rect 12529 14365 12541 14399
rect 12575 14365 12587 14399
rect 12529 14359 12587 14365
rect 12713 14399 12771 14405
rect 12713 14365 12725 14399
rect 12759 14396 12771 14399
rect 12894 14396 12900 14408
rect 12759 14368 12900 14396
rect 12759 14365 12771 14368
rect 12713 14359 12771 14365
rect 11992 14300 12296 14328
rect 12544 14328 12572 14359
rect 12894 14356 12900 14368
rect 12952 14356 12958 14408
rect 13004 14405 13032 14436
rect 12989 14399 13047 14405
rect 12989 14365 13001 14399
rect 13035 14365 13047 14399
rect 12989 14359 13047 14365
rect 13262 14356 13268 14408
rect 13320 14356 13326 14408
rect 14936 14405 14964 14504
rect 16025 14501 16037 14535
rect 16071 14532 16083 14535
rect 23106 14532 23112 14544
rect 16071 14504 19932 14532
rect 16071 14501 16083 14504
rect 16025 14495 16083 14501
rect 15378 14424 15384 14476
rect 15436 14424 15442 14476
rect 16546 14436 17832 14464
rect 14553 14399 14611 14405
rect 14553 14365 14565 14399
rect 14599 14365 14611 14399
rect 14553 14359 14611 14365
rect 14921 14399 14979 14405
rect 14921 14365 14933 14399
rect 14967 14396 14979 14399
rect 15010 14396 15016 14408
rect 14967 14368 15016 14396
rect 14967 14365 14979 14368
rect 14921 14359 14979 14365
rect 14090 14328 14096 14340
rect 12544 14300 14096 14328
rect 11388 14288 11394 14300
rect 14090 14288 14096 14300
rect 14148 14328 14154 14340
rect 14568 14328 14596 14359
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15102 14356 15108 14408
rect 15160 14356 15166 14408
rect 15289 14399 15347 14405
rect 15289 14365 15301 14399
rect 15335 14365 15347 14399
rect 15396 14396 15424 14424
rect 16546 14405 16574 14436
rect 16209 14399 16267 14405
rect 16209 14396 16221 14399
rect 15396 14368 16221 14396
rect 15289 14359 15347 14365
rect 16209 14365 16221 14368
rect 16255 14365 16267 14399
rect 16209 14359 16267 14365
rect 16531 14399 16589 14405
rect 16531 14365 16543 14399
rect 16577 14365 16589 14399
rect 16531 14359 16589 14365
rect 16669 14399 16727 14405
rect 16669 14365 16681 14399
rect 16715 14365 16727 14399
rect 16669 14359 16727 14365
rect 14148 14300 14596 14328
rect 14148 14288 14154 14300
rect 14642 14288 14648 14340
rect 14700 14328 14706 14340
rect 15304 14328 15332 14359
rect 14700 14300 15332 14328
rect 14700 14288 14706 14300
rect 9674 14260 9680 14272
rect 9508 14232 9680 14260
rect 9125 14223 9183 14229
rect 9674 14220 9680 14232
rect 9732 14220 9738 14272
rect 11238 14220 11244 14272
rect 11296 14260 11302 14272
rect 11974 14260 11980 14272
rect 11296 14232 11980 14260
rect 11296 14220 11302 14232
rect 11974 14220 11980 14232
rect 12032 14220 12038 14272
rect 12986 14220 12992 14272
rect 13044 14260 13050 14272
rect 13081 14263 13139 14269
rect 13081 14260 13093 14263
rect 13044 14232 13093 14260
rect 13044 14220 13050 14232
rect 13081 14229 13093 14232
rect 13127 14260 13139 14263
rect 13354 14260 13360 14272
rect 13127 14232 13360 14260
rect 13127 14229 13139 14232
rect 13081 14223 13139 14229
rect 13354 14220 13360 14232
rect 13412 14220 13418 14272
rect 13446 14220 13452 14272
rect 13504 14220 13510 14272
rect 13906 14220 13912 14272
rect 13964 14260 13970 14272
rect 14660 14260 14688 14288
rect 13964 14232 14688 14260
rect 15304 14260 15332 14300
rect 15470 14288 15476 14340
rect 15528 14328 15534 14340
rect 16301 14331 16359 14337
rect 16301 14328 16313 14331
rect 15528 14300 16313 14328
rect 15528 14288 15534 14300
rect 16301 14297 16313 14300
rect 16347 14297 16359 14331
rect 16301 14291 16359 14297
rect 16393 14331 16451 14337
rect 16393 14297 16405 14331
rect 16439 14297 16451 14331
rect 16684 14328 16712 14359
rect 16942 14356 16948 14408
rect 17000 14356 17006 14408
rect 17126 14356 17132 14408
rect 17184 14356 17190 14408
rect 17678 14328 17684 14340
rect 16684 14300 17684 14328
rect 16393 14291 16451 14297
rect 15746 14260 15752 14272
rect 15304 14232 15752 14260
rect 13964 14220 13970 14232
rect 15746 14220 15752 14232
rect 15804 14220 15810 14272
rect 16408 14260 16436 14291
rect 17678 14288 17684 14300
rect 17736 14288 17742 14340
rect 17804 14328 17832 14436
rect 17880 14405 17908 14504
rect 19337 14467 19395 14473
rect 19337 14433 19349 14467
rect 19383 14464 19395 14467
rect 19426 14464 19432 14476
rect 19383 14436 19432 14464
rect 19383 14433 19395 14436
rect 19337 14427 19395 14433
rect 19426 14424 19432 14436
rect 19484 14424 19490 14476
rect 19904 14473 19932 14504
rect 21376 14504 23112 14532
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14433 19947 14467
rect 19889 14427 19947 14433
rect 17865 14399 17923 14405
rect 17865 14365 17877 14399
rect 17911 14365 17923 14399
rect 20349 14399 20407 14405
rect 17865 14359 17923 14365
rect 17972 14368 19564 14396
rect 17972 14328 18000 14368
rect 17804 14300 18000 14328
rect 18506 14288 18512 14340
rect 18564 14288 18570 14340
rect 18785 14331 18843 14337
rect 18785 14297 18797 14331
rect 18831 14328 18843 14331
rect 19334 14328 19340 14340
rect 18831 14300 19340 14328
rect 18831 14297 18843 14300
rect 18785 14291 18843 14297
rect 19334 14288 19340 14300
rect 19392 14288 19398 14340
rect 19429 14331 19487 14337
rect 19429 14297 19441 14331
rect 19475 14297 19487 14331
rect 19536 14328 19564 14368
rect 20349 14365 20361 14399
rect 20395 14396 20407 14399
rect 20622 14396 20628 14408
rect 20395 14368 20628 14396
rect 20395 14365 20407 14368
rect 20349 14359 20407 14365
rect 20622 14356 20628 14368
rect 20680 14356 20686 14408
rect 20901 14399 20959 14405
rect 20901 14365 20913 14399
rect 20947 14396 20959 14399
rect 21082 14396 21088 14408
rect 20947 14368 21088 14396
rect 20947 14365 20959 14368
rect 20901 14359 20959 14365
rect 21082 14356 21088 14368
rect 21140 14356 21146 14408
rect 21376 14405 21404 14504
rect 23106 14492 23112 14504
rect 23164 14492 23170 14544
rect 23750 14492 23756 14544
rect 23808 14492 23814 14544
rect 22066 14436 22600 14464
rect 21361 14399 21419 14405
rect 21361 14365 21373 14399
rect 21407 14365 21419 14399
rect 21361 14359 21419 14365
rect 21821 14399 21879 14405
rect 21821 14365 21833 14399
rect 21867 14396 21879 14399
rect 22066 14396 22094 14436
rect 22572 14408 22600 14436
rect 21867 14368 22094 14396
rect 21867 14365 21879 14368
rect 21821 14359 21879 14365
rect 22278 14356 22284 14408
rect 22336 14356 22342 14408
rect 22554 14356 22560 14408
rect 22612 14396 22618 14408
rect 23201 14399 23259 14405
rect 23201 14396 23213 14399
rect 22612 14368 23213 14396
rect 22612 14356 22618 14368
rect 23201 14365 23213 14368
rect 23247 14365 23259 14399
rect 23201 14359 23259 14365
rect 23658 14328 23664 14340
rect 19536 14300 23664 14328
rect 19429 14291 19487 14297
rect 16758 14260 16764 14272
rect 16408 14232 16764 14260
rect 16758 14220 16764 14232
rect 16816 14220 16822 14272
rect 18524 14260 18552 14288
rect 19444 14260 19472 14291
rect 23658 14288 23664 14300
rect 23716 14288 23722 14340
rect 18524 14232 19472 14260
rect 20070 14220 20076 14272
rect 20128 14260 20134 14272
rect 20165 14263 20223 14269
rect 20165 14260 20177 14263
rect 20128 14232 20177 14260
rect 20128 14220 20134 14232
rect 20165 14229 20177 14232
rect 20211 14229 20223 14263
rect 20165 14223 20223 14229
rect 22005 14263 22063 14269
rect 22005 14229 22017 14263
rect 22051 14260 22063 14263
rect 23750 14260 23756 14272
rect 22051 14232 23756 14260
rect 22051 14229 22063 14232
rect 22005 14223 22063 14229
rect 23750 14220 23756 14232
rect 23808 14220 23814 14272
rect 1104 14170 24840 14192
rect 1104 14118 8214 14170
rect 8266 14118 8278 14170
rect 8330 14118 8342 14170
rect 8394 14118 8406 14170
rect 8458 14118 8470 14170
rect 8522 14118 16214 14170
rect 16266 14118 16278 14170
rect 16330 14118 16342 14170
rect 16394 14118 16406 14170
rect 16458 14118 16470 14170
rect 16522 14118 24214 14170
rect 24266 14118 24278 14170
rect 24330 14118 24342 14170
rect 24394 14118 24406 14170
rect 24458 14118 24470 14170
rect 24522 14118 24840 14170
rect 1104 14096 24840 14118
rect 2130 14016 2136 14068
rect 2188 14056 2194 14068
rect 2188 14028 3280 14056
rect 2188 14016 2194 14028
rect 2866 13948 2872 14000
rect 2924 13948 2930 14000
rect 3252 13988 3280 14028
rect 3326 14016 3332 14068
rect 3384 14016 3390 14068
rect 3970 14016 3976 14068
rect 4028 14016 4034 14068
rect 5902 14056 5908 14068
rect 4540 14028 5908 14056
rect 3605 13991 3663 13997
rect 3605 13988 3617 13991
rect 3252 13960 3617 13988
rect 3605 13957 3617 13960
rect 3651 13957 3663 13991
rect 3605 13951 3663 13957
rect 3821 13991 3879 13997
rect 3821 13957 3833 13991
rect 3867 13988 3879 13991
rect 4540 13988 4568 14028
rect 5902 14016 5908 14028
rect 5960 14016 5966 14068
rect 6457 14059 6515 14065
rect 6457 14025 6469 14059
rect 6503 14025 6515 14059
rect 6457 14019 6515 14025
rect 6625 14059 6683 14065
rect 6625 14025 6637 14059
rect 6671 14056 6683 14059
rect 6914 14056 6920 14068
rect 6671 14028 6920 14056
rect 6671 14025 6683 14028
rect 6625 14019 6683 14025
rect 6472 13988 6500 14019
rect 6914 14016 6920 14028
rect 6972 14016 6978 14068
rect 8110 14016 8116 14068
rect 8168 14056 8174 14068
rect 8849 14059 8907 14065
rect 8849 14056 8861 14059
rect 8168 14028 8861 14056
rect 8168 14016 8174 14028
rect 8849 14025 8861 14028
rect 8895 14025 8907 14059
rect 8849 14019 8907 14025
rect 9214 14016 9220 14068
rect 9272 14056 9278 14068
rect 9325 14059 9383 14065
rect 9325 14056 9337 14059
rect 9272 14028 9337 14056
rect 9272 14016 9278 14028
rect 9325 14025 9337 14028
rect 9371 14025 9383 14059
rect 9325 14019 9383 14025
rect 10962 14016 10968 14068
rect 11020 14056 11026 14068
rect 12066 14056 12072 14068
rect 11020 14028 12072 14056
rect 11020 14016 11026 14028
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 13354 14065 13360 14068
rect 13331 14059 13360 14065
rect 13331 14025 13343 14059
rect 13331 14019 13360 14025
rect 13354 14016 13360 14019
rect 13412 14016 13418 14068
rect 14090 14016 14096 14068
rect 14148 14056 14154 14068
rect 14829 14059 14887 14065
rect 14829 14056 14841 14059
rect 14148 14028 14841 14056
rect 14148 14016 14154 14028
rect 14829 14025 14841 14028
rect 14875 14025 14887 14059
rect 14829 14019 14887 14025
rect 15654 14016 15660 14068
rect 15712 14056 15718 14068
rect 16666 14056 16672 14068
rect 15712 14028 16672 14056
rect 15712 14016 15718 14028
rect 16666 14016 16672 14028
rect 16724 14016 16730 14068
rect 16758 14016 16764 14068
rect 16816 14016 16822 14068
rect 17034 14016 17040 14068
rect 17092 14056 17098 14068
rect 20073 14059 20131 14065
rect 20073 14056 20085 14059
rect 17092 14028 20085 14056
rect 17092 14016 17098 14028
rect 20073 14025 20085 14028
rect 20119 14056 20131 14059
rect 20806 14056 20812 14068
rect 20119 14028 20812 14056
rect 20119 14025 20131 14028
rect 20073 14019 20131 14025
rect 20806 14016 20812 14028
rect 20864 14016 20870 14068
rect 21082 14016 21088 14068
rect 21140 14056 21146 14068
rect 21910 14056 21916 14068
rect 21140 14028 21916 14056
rect 21140 14016 21146 14028
rect 21910 14016 21916 14028
rect 21968 14016 21974 14068
rect 3867 13960 4568 13988
rect 5382 13960 6500 13988
rect 3867 13957 3879 13960
rect 3821 13951 3879 13957
rect 1486 13880 1492 13932
rect 1544 13920 1550 13932
rect 1581 13923 1639 13929
rect 1581 13920 1593 13923
rect 1544 13892 1593 13920
rect 1544 13880 1550 13892
rect 1581 13889 1593 13892
rect 1627 13889 1639 13923
rect 3620 13920 3648 13951
rect 6822 13948 6828 14000
rect 6880 13948 6886 14000
rect 9030 13988 9036 14000
rect 8602 13960 9036 13988
rect 9030 13948 9036 13960
rect 9088 13948 9094 14000
rect 9125 13991 9183 13997
rect 9125 13957 9137 13991
rect 9171 13957 9183 13991
rect 11054 13988 11060 14000
rect 9125 13951 9183 13957
rect 10060 13960 11060 13988
rect 4062 13920 4068 13932
rect 3620 13892 4068 13920
rect 1581 13883 1639 13889
rect 4062 13880 4068 13892
rect 4120 13880 4126 13932
rect 6089 13923 6147 13929
rect 6089 13889 6101 13923
rect 6135 13920 6147 13923
rect 7098 13920 7104 13932
rect 6135 13892 7104 13920
rect 6135 13889 6147 13892
rect 6089 13883 6147 13889
rect 7098 13880 7104 13892
rect 7156 13880 7162 13932
rect 8938 13880 8944 13932
rect 8996 13920 9002 13932
rect 9140 13920 9168 13951
rect 10060 13929 10088 13960
rect 11054 13948 11060 13960
rect 11112 13948 11118 14000
rect 11149 13991 11207 13997
rect 11149 13957 11161 13991
rect 11195 13988 11207 13991
rect 11195 13960 17908 13988
rect 11195 13957 11207 13960
rect 11149 13951 11207 13957
rect 8996 13892 9168 13920
rect 10045 13923 10103 13929
rect 8996 13880 9002 13892
rect 10045 13889 10057 13923
rect 10091 13889 10103 13923
rect 10045 13883 10103 13889
rect 10229 13923 10287 13929
rect 10229 13889 10241 13923
rect 10275 13920 10287 13923
rect 10318 13920 10324 13932
rect 10275 13892 10324 13920
rect 10275 13889 10287 13892
rect 10229 13883 10287 13889
rect 10318 13880 10324 13892
rect 10376 13880 10382 13932
rect 10502 13880 10508 13932
rect 10560 13880 10566 13932
rect 10778 13880 10784 13932
rect 10836 13920 10842 13932
rect 10836 13892 11192 13920
rect 10836 13880 10842 13892
rect 1854 13812 1860 13864
rect 1912 13812 1918 13864
rect 7374 13812 7380 13864
rect 7432 13812 7438 13864
rect 9674 13812 9680 13864
rect 9732 13852 9738 13864
rect 10594 13852 10600 13864
rect 9732 13824 10600 13852
rect 9732 13812 9738 13824
rect 10594 13812 10600 13824
rect 10652 13852 10658 13864
rect 10689 13855 10747 13861
rect 10689 13852 10701 13855
rect 10652 13824 10701 13852
rect 10652 13812 10658 13824
rect 10689 13821 10701 13824
rect 10735 13821 10747 13855
rect 10689 13815 10747 13821
rect 10873 13855 10931 13861
rect 10873 13821 10885 13855
rect 10919 13821 10931 13855
rect 10873 13815 10931 13821
rect 10888 13784 10916 13815
rect 10962 13812 10968 13864
rect 11020 13812 11026 13864
rect 11164 13852 11192 13892
rect 11606 13880 11612 13932
rect 11664 13920 11670 13932
rect 11664 13892 11836 13920
rect 11664 13880 11670 13892
rect 11808 13852 11836 13892
rect 11882 13880 11888 13932
rect 11940 13880 11946 13932
rect 11977 13923 12035 13929
rect 11977 13889 11989 13923
rect 12023 13889 12035 13923
rect 11977 13883 12035 13889
rect 11992 13852 12020 13883
rect 12066 13880 12072 13932
rect 12124 13920 12130 13932
rect 12253 13923 12311 13929
rect 12253 13920 12265 13923
rect 12124 13892 12265 13920
rect 12124 13880 12130 13892
rect 12253 13889 12265 13892
rect 12299 13920 12311 13923
rect 12802 13920 12808 13932
rect 12299 13892 12808 13920
rect 12299 13889 12311 13892
rect 12253 13883 12311 13889
rect 12802 13880 12808 13892
rect 12860 13880 12866 13932
rect 13262 13880 13268 13932
rect 13320 13880 13326 13932
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 14090 13880 14096 13932
rect 14148 13880 14154 13932
rect 14829 13923 14887 13929
rect 14829 13889 14841 13923
rect 14875 13889 14887 13923
rect 14829 13883 14887 13889
rect 12992 13864 13044 13870
rect 12618 13852 12624 13864
rect 11164 13824 11652 13852
rect 11808 13824 12624 13852
rect 11146 13784 11152 13796
rect 3252 13756 3832 13784
rect 10888 13756 11152 13784
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 3252 13716 3280 13756
rect 3804 13725 3832 13756
rect 11146 13744 11152 13756
rect 11204 13784 11210 13796
rect 11330 13784 11336 13796
rect 11204 13756 11336 13784
rect 11204 13744 11210 13756
rect 11330 13744 11336 13756
rect 11388 13744 11394 13796
rect 11624 13793 11652 13824
rect 12618 13812 12624 13824
rect 12676 13852 12682 13864
rect 12676 13824 12992 13852
rect 12676 13812 12682 13824
rect 13998 13812 14004 13864
rect 14056 13852 14062 13864
rect 14844 13852 14872 13883
rect 15010 13880 15016 13932
rect 15068 13880 15074 13932
rect 15194 13880 15200 13932
rect 15252 13880 15258 13932
rect 16025 13923 16083 13929
rect 16025 13889 16037 13923
rect 16071 13920 16083 13923
rect 16114 13920 16120 13932
rect 16071 13892 16120 13920
rect 16071 13889 16083 13892
rect 16025 13883 16083 13889
rect 16114 13880 16120 13892
rect 16172 13880 16178 13932
rect 16942 13880 16948 13932
rect 17000 13880 17006 13932
rect 17126 13880 17132 13932
rect 17184 13880 17190 13932
rect 17221 13923 17279 13929
rect 17221 13889 17233 13923
rect 17267 13889 17279 13923
rect 17221 13883 17279 13889
rect 14918 13852 14924 13864
rect 14056 13824 14924 13852
rect 14056 13812 14062 13824
rect 14918 13812 14924 13824
rect 14976 13852 14982 13864
rect 15933 13855 15991 13861
rect 15933 13852 15945 13855
rect 14976 13824 15945 13852
rect 14976 13812 14982 13824
rect 15933 13821 15945 13824
rect 15979 13852 15991 13855
rect 16666 13852 16672 13864
rect 15979 13824 16672 13852
rect 15979 13821 15991 13824
rect 15933 13815 15991 13821
rect 16666 13812 16672 13824
rect 16724 13812 16730 13864
rect 17236 13852 17264 13883
rect 17586 13880 17592 13932
rect 17644 13880 17650 13932
rect 17880 13929 17908 13960
rect 19426 13948 19432 14000
rect 19484 13988 19490 14000
rect 20625 13991 20683 13997
rect 20625 13988 20637 13991
rect 19484 13960 20637 13988
rect 19484 13948 19490 13960
rect 20625 13957 20637 13960
rect 20671 13957 20683 13991
rect 20625 13951 20683 13957
rect 22005 13991 22063 13997
rect 22005 13957 22017 13991
rect 22051 13988 22063 13991
rect 22554 13988 22560 14000
rect 22051 13960 22560 13988
rect 22051 13957 22063 13960
rect 22005 13951 22063 13957
rect 22554 13948 22560 13960
rect 22612 13948 22618 14000
rect 22833 13991 22891 13997
rect 22833 13957 22845 13991
rect 22879 13988 22891 13991
rect 22879 13960 23612 13988
rect 22879 13957 22891 13960
rect 22833 13951 22891 13957
rect 17865 13923 17923 13929
rect 17865 13889 17877 13923
rect 17911 13920 17923 13923
rect 18322 13920 18328 13932
rect 17911 13892 18328 13920
rect 17911 13889 17923 13892
rect 17865 13883 17923 13889
rect 18322 13880 18328 13892
rect 18380 13880 18386 13932
rect 19334 13880 19340 13932
rect 19392 13880 19398 13932
rect 19536 13920 19748 13926
rect 19889 13923 19947 13929
rect 19889 13920 19901 13923
rect 19444 13898 19901 13920
rect 19444 13892 19564 13898
rect 19720 13892 19901 13898
rect 17310 13852 17316 13864
rect 17236 13824 17316 13852
rect 17310 13812 17316 13824
rect 17368 13852 17374 13864
rect 19444 13852 19472 13892
rect 19889 13889 19901 13892
rect 19935 13920 19947 13923
rect 19978 13920 19984 13932
rect 19935 13892 19984 13920
rect 19935 13889 19947 13892
rect 19889 13883 19947 13889
rect 19978 13880 19984 13892
rect 20036 13880 20042 13932
rect 21545 13923 21603 13929
rect 21545 13889 21557 13923
rect 21591 13920 21603 13923
rect 22094 13920 22100 13932
rect 21591 13892 22100 13920
rect 21591 13889 21603 13892
rect 21545 13883 21603 13889
rect 22094 13880 22100 13892
rect 22152 13880 22158 13932
rect 22186 13880 22192 13932
rect 22244 13880 22250 13932
rect 23477 13923 23535 13929
rect 23477 13889 23489 13923
rect 23523 13889 23535 13923
rect 23584 13920 23612 13960
rect 23750 13948 23756 14000
rect 23808 13948 23814 14000
rect 23845 13991 23903 13997
rect 23845 13957 23857 13991
rect 23891 13988 23903 13991
rect 23934 13988 23940 14000
rect 23891 13960 23940 13988
rect 23891 13957 23903 13960
rect 23845 13951 23903 13957
rect 23860 13920 23888 13951
rect 23934 13948 23940 13960
rect 23992 13948 23998 14000
rect 23584 13892 23888 13920
rect 23477 13883 23535 13889
rect 19705 13855 19763 13861
rect 19705 13852 19717 13855
rect 17368 13824 19472 13852
rect 19536 13824 19717 13852
rect 17368 13812 17374 13824
rect 12992 13806 13044 13812
rect 11609 13787 11667 13793
rect 11609 13753 11621 13787
rect 11655 13753 11667 13787
rect 11974 13784 11980 13796
rect 11609 13747 11667 13753
rect 11808 13756 11980 13784
rect 11808 13728 11836 13756
rect 11974 13744 11980 13756
rect 12032 13744 12038 13796
rect 17126 13744 17132 13796
rect 17184 13784 17190 13796
rect 19536 13784 19564 13824
rect 19705 13821 19717 13824
rect 19751 13852 19763 13855
rect 23492 13852 23520 13883
rect 24026 13852 24032 13864
rect 19751 13824 20760 13852
rect 23492 13824 24032 13852
rect 19751 13821 19763 13824
rect 19705 13815 19763 13821
rect 17184 13756 19564 13784
rect 20732 13784 20760 13824
rect 24026 13812 24032 13824
rect 24084 13852 24090 13864
rect 24305 13855 24363 13861
rect 24305 13852 24317 13855
rect 24084 13824 24317 13852
rect 24084 13812 24090 13824
rect 24305 13821 24317 13824
rect 24351 13821 24363 13855
rect 24305 13815 24363 13821
rect 21542 13784 21548 13796
rect 20732 13756 21548 13784
rect 17184 13744 17190 13756
rect 21542 13744 21548 13756
rect 21600 13744 21606 13796
rect 2004 13688 3280 13716
rect 3789 13719 3847 13725
rect 2004 13676 2010 13688
rect 3789 13685 3801 13719
rect 3835 13685 3847 13719
rect 3789 13679 3847 13685
rect 3970 13676 3976 13728
rect 4028 13716 4034 13728
rect 4341 13719 4399 13725
rect 4341 13716 4353 13719
rect 4028 13688 4353 13716
rect 4028 13676 4034 13688
rect 4341 13685 4353 13688
rect 4387 13685 4399 13719
rect 4341 13679 4399 13685
rect 5831 13719 5889 13725
rect 5831 13685 5843 13719
rect 5877 13716 5889 13719
rect 6178 13716 6184 13728
rect 5877 13688 6184 13716
rect 5877 13685 5889 13688
rect 5831 13679 5889 13685
rect 6178 13676 6184 13688
rect 6236 13676 6242 13728
rect 6641 13719 6699 13725
rect 6641 13685 6653 13719
rect 6687 13716 6699 13719
rect 8754 13716 8760 13728
rect 6687 13688 8760 13716
rect 6687 13685 6699 13688
rect 6641 13679 6699 13685
rect 8754 13676 8760 13688
rect 8812 13716 8818 13728
rect 9306 13716 9312 13728
rect 8812 13688 9312 13716
rect 8812 13676 8818 13688
rect 9306 13676 9312 13688
rect 9364 13676 9370 13728
rect 9490 13676 9496 13728
rect 9548 13676 9554 13728
rect 10134 13676 10140 13728
rect 10192 13676 10198 13728
rect 11790 13676 11796 13728
rect 11848 13676 11854 13728
rect 11882 13676 11888 13728
rect 11940 13716 11946 13728
rect 12345 13719 12403 13725
rect 12345 13716 12357 13719
rect 11940 13688 12357 13716
rect 11940 13676 11946 13688
rect 12345 13685 12357 13688
rect 12391 13716 12403 13719
rect 13814 13716 13820 13728
rect 12391 13688 13820 13716
rect 12391 13685 12403 13688
rect 12345 13679 12403 13685
rect 13814 13676 13820 13688
rect 13872 13676 13878 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 15010 13716 15016 13728
rect 14884 13688 15016 13716
rect 14884 13676 14890 13688
rect 15010 13676 15016 13688
rect 15068 13716 15074 13728
rect 15841 13719 15899 13725
rect 15841 13716 15853 13719
rect 15068 13688 15853 13716
rect 15068 13676 15074 13688
rect 15841 13685 15853 13688
rect 15887 13685 15899 13719
rect 15841 13679 15899 13685
rect 20533 13719 20591 13725
rect 20533 13685 20545 13719
rect 20579 13716 20591 13719
rect 20622 13716 20628 13728
rect 20579 13688 20628 13716
rect 20579 13685 20591 13688
rect 20533 13679 20591 13685
rect 20622 13676 20628 13688
rect 20680 13676 20686 13728
rect 21450 13676 21456 13728
rect 21508 13676 21514 13728
rect 1104 13626 24840 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 20214 13626
rect 20266 13574 20278 13626
rect 20330 13574 20342 13626
rect 20394 13574 20406 13626
rect 20458 13574 20470 13626
rect 20522 13574 24840 13626
rect 1104 13552 24840 13574
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2041 13515 2099 13521
rect 2041 13512 2053 13515
rect 2004 13484 2053 13512
rect 2004 13472 2010 13484
rect 2041 13481 2053 13484
rect 2087 13481 2099 13515
rect 2041 13475 2099 13481
rect 2225 13515 2283 13521
rect 2225 13481 2237 13515
rect 2271 13512 2283 13515
rect 2866 13512 2872 13524
rect 2271 13484 2872 13512
rect 2271 13481 2283 13484
rect 2225 13475 2283 13481
rect 2866 13472 2872 13484
rect 2924 13472 2930 13524
rect 6178 13472 6184 13524
rect 6236 13472 6242 13524
rect 7374 13472 7380 13524
rect 7432 13512 7438 13524
rect 7837 13515 7895 13521
rect 7837 13512 7849 13515
rect 7432 13484 7849 13512
rect 7432 13472 7438 13484
rect 7837 13481 7849 13484
rect 7883 13481 7895 13515
rect 7837 13475 7895 13481
rect 9306 13472 9312 13524
rect 9364 13472 9370 13524
rect 11701 13515 11759 13521
rect 11701 13481 11713 13515
rect 11747 13512 11759 13515
rect 11974 13512 11980 13524
rect 11747 13484 11980 13512
rect 11747 13481 11759 13484
rect 11701 13475 11759 13481
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12805 13515 12863 13521
rect 12805 13481 12817 13515
rect 12851 13512 12863 13515
rect 14458 13512 14464 13524
rect 12851 13484 14464 13512
rect 12851 13481 12863 13484
rect 12805 13475 12863 13481
rect 14458 13472 14464 13484
rect 14516 13472 14522 13524
rect 15194 13472 15200 13524
rect 15252 13512 15258 13524
rect 16114 13512 16120 13524
rect 15252 13484 16120 13512
rect 15252 13472 15258 13484
rect 16114 13472 16120 13484
rect 16172 13512 16178 13524
rect 16577 13515 16635 13521
rect 16577 13512 16589 13515
rect 16172 13484 16589 13512
rect 16172 13472 16178 13484
rect 16577 13481 16589 13484
rect 16623 13481 16635 13515
rect 16577 13475 16635 13481
rect 16942 13472 16948 13524
rect 17000 13472 17006 13524
rect 22462 13512 22468 13524
rect 17236 13484 22468 13512
rect 1854 13404 1860 13456
rect 1912 13444 1918 13456
rect 2501 13447 2559 13453
rect 2501 13444 2513 13447
rect 1912 13416 2513 13444
rect 1912 13404 1918 13416
rect 2501 13413 2513 13416
rect 2547 13413 2559 13447
rect 2501 13407 2559 13413
rect 10870 13404 10876 13456
rect 10928 13444 10934 13456
rect 17236 13444 17264 13484
rect 22462 13472 22468 13484
rect 22520 13512 22526 13524
rect 22520 13484 23244 13512
rect 22520 13472 22526 13484
rect 10928 13416 17264 13444
rect 18785 13447 18843 13453
rect 10928 13404 10934 13416
rect 18785 13413 18797 13447
rect 18831 13444 18843 13447
rect 19426 13444 19432 13456
rect 18831 13416 19432 13444
rect 18831 13413 18843 13416
rect 18785 13407 18843 13413
rect 19426 13404 19432 13416
rect 19484 13404 19490 13456
rect 20993 13447 21051 13453
rect 20993 13413 21005 13447
rect 21039 13444 21051 13447
rect 22186 13444 22192 13456
rect 21039 13416 22192 13444
rect 21039 13413 21051 13416
rect 20993 13407 21051 13413
rect 22186 13404 22192 13416
rect 22244 13444 22250 13456
rect 22649 13447 22707 13453
rect 22649 13444 22661 13447
rect 22244 13416 22661 13444
rect 22244 13404 22250 13416
rect 22649 13413 22661 13416
rect 22695 13413 22707 13447
rect 22649 13407 22707 13413
rect 1946 13336 1952 13388
rect 2004 13376 2010 13388
rect 2222 13376 2228 13388
rect 2004 13348 2228 13376
rect 2004 13336 2010 13348
rect 2222 13336 2228 13348
rect 2280 13336 2286 13388
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13376 3203 13379
rect 3418 13376 3424 13388
rect 3191 13348 3424 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 3418 13336 3424 13348
rect 3476 13376 3482 13388
rect 4890 13376 4896 13388
rect 3476 13348 4896 13376
rect 3476 13336 3482 13348
rect 4890 13336 4896 13348
rect 4948 13376 4954 13388
rect 5537 13379 5595 13385
rect 5537 13376 5549 13379
rect 4948 13348 5549 13376
rect 4948 13336 4954 13348
rect 5537 13345 5549 13348
rect 5583 13345 5595 13379
rect 5537 13339 5595 13345
rect 5721 13379 5779 13385
rect 5721 13345 5733 13379
rect 5767 13376 5779 13379
rect 6730 13376 6736 13388
rect 5767 13348 6736 13376
rect 5767 13345 5779 13348
rect 5721 13339 5779 13345
rect 6730 13336 6736 13348
rect 6788 13336 6794 13388
rect 8110 13336 8116 13388
rect 8168 13376 8174 13388
rect 8481 13379 8539 13385
rect 8168 13348 8248 13376
rect 8168 13336 8174 13348
rect 2130 13308 2136 13320
rect 1872 13280 2136 13308
rect 1872 13252 1900 13280
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 2869 13311 2927 13317
rect 2869 13277 2881 13311
rect 2915 13308 2927 13311
rect 3326 13308 3332 13320
rect 2915 13280 3332 13308
rect 2915 13277 2927 13280
rect 2869 13271 2927 13277
rect 3326 13268 3332 13280
rect 3384 13268 3390 13320
rect 8220 13317 8248 13348
rect 8481 13345 8493 13379
rect 8527 13376 8539 13379
rect 8570 13376 8576 13388
rect 8527 13348 8576 13376
rect 8527 13345 8539 13348
rect 8481 13339 8539 13345
rect 8570 13336 8576 13348
rect 8628 13336 8634 13388
rect 10229 13379 10287 13385
rect 10229 13345 10241 13379
rect 10275 13376 10287 13379
rect 10778 13376 10784 13388
rect 10275 13348 10784 13376
rect 10275 13345 10287 13348
rect 10229 13339 10287 13345
rect 10778 13336 10784 13348
rect 10836 13336 10842 13388
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13376 12587 13379
rect 13170 13376 13176 13388
rect 12575 13348 13176 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 13170 13336 13176 13348
rect 13228 13336 13234 13388
rect 15286 13376 15292 13388
rect 13372 13348 15292 13376
rect 8205 13311 8263 13317
rect 8205 13277 8217 13311
rect 8251 13277 8263 13311
rect 8205 13271 8263 13277
rect 9769 13311 9827 13317
rect 9769 13277 9781 13311
rect 9815 13308 9827 13311
rect 9858 13308 9864 13320
rect 9815 13280 9864 13308
rect 9815 13277 9827 13280
rect 9769 13271 9827 13277
rect 9858 13268 9864 13280
rect 9916 13268 9922 13320
rect 9953 13311 10011 13317
rect 9953 13277 9965 13311
rect 9999 13277 10011 13311
rect 9953 13271 10011 13277
rect 1854 13200 1860 13252
rect 1912 13200 1918 13252
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 5813 13243 5871 13249
rect 5813 13240 5825 13243
rect 4028 13212 5825 13240
rect 4028 13200 4034 13212
rect 5813 13209 5825 13212
rect 5859 13209 5871 13243
rect 5813 13203 5871 13209
rect 8110 13200 8116 13252
rect 8168 13240 8174 13252
rect 8297 13243 8355 13249
rect 8297 13240 8309 13243
rect 8168 13212 8309 13240
rect 8168 13200 8174 13212
rect 8297 13209 8309 13212
rect 8343 13209 8355 13243
rect 8297 13203 8355 13209
rect 8938 13200 8944 13252
rect 8996 13240 9002 13252
rect 9306 13249 9312 13252
rect 9293 13243 9312 13249
rect 8996 13212 9260 13240
rect 8996 13200 9002 13212
rect 1302 13132 1308 13184
rect 1360 13172 1366 13184
rect 1489 13175 1547 13181
rect 1489 13172 1501 13175
rect 1360 13144 1501 13172
rect 1360 13132 1366 13144
rect 1489 13141 1501 13144
rect 1535 13141 1547 13175
rect 1489 13135 1547 13141
rect 2038 13132 2044 13184
rect 2096 13181 2102 13184
rect 2096 13175 2115 13181
rect 2103 13141 2115 13175
rect 2096 13135 2115 13141
rect 2961 13175 3019 13181
rect 2961 13141 2973 13175
rect 3007 13172 3019 13175
rect 3602 13172 3608 13184
rect 3007 13144 3608 13172
rect 3007 13141 3019 13144
rect 2961 13135 3019 13141
rect 2096 13132 2102 13135
rect 3602 13132 3608 13144
rect 3660 13132 3666 13184
rect 9122 13132 9128 13184
rect 9180 13132 9186 13184
rect 9232 13172 9260 13212
rect 9293 13209 9305 13243
rect 9293 13203 9312 13209
rect 9306 13200 9312 13203
rect 9364 13200 9370 13252
rect 9493 13243 9551 13249
rect 9493 13209 9505 13243
rect 9539 13240 9551 13243
rect 9968 13240 9996 13271
rect 10318 13268 10324 13320
rect 10376 13308 10382 13320
rect 11057 13311 11115 13317
rect 11057 13308 11069 13311
rect 10376 13280 11069 13308
rect 10376 13268 10382 13280
rect 11057 13277 11069 13280
rect 11103 13308 11115 13311
rect 11146 13308 11152 13320
rect 11103 13280 11152 13308
rect 11103 13277 11115 13280
rect 11057 13271 11115 13277
rect 11146 13268 11152 13280
rect 11204 13268 11210 13320
rect 11900 13280 12388 13308
rect 9539 13212 9996 13240
rect 9539 13209 9551 13212
rect 9493 13203 9551 13209
rect 9508 13172 9536 13203
rect 10686 13200 10692 13252
rect 10744 13240 10750 13252
rect 11698 13249 11704 13252
rect 10781 13243 10839 13249
rect 10781 13240 10793 13243
rect 10744 13212 10793 13240
rect 10744 13200 10750 13212
rect 10781 13209 10793 13212
rect 10827 13209 10839 13243
rect 10781 13203 10839 13209
rect 11685 13243 11704 13249
rect 11685 13209 11697 13243
rect 11685 13203 11704 13209
rect 11698 13200 11704 13203
rect 11756 13200 11762 13252
rect 11900 13249 11928 13280
rect 11885 13243 11943 13249
rect 11885 13209 11897 13243
rect 11931 13209 11943 13243
rect 12360 13240 12388 13280
rect 12618 13268 12624 13320
rect 12676 13268 12682 13320
rect 12894 13268 12900 13320
rect 12952 13308 12958 13320
rect 13372 13317 13400 13348
rect 15286 13336 15292 13348
rect 15344 13336 15350 13388
rect 15746 13336 15752 13388
rect 15804 13376 15810 13388
rect 15804 13348 16620 13376
rect 15804 13336 15810 13348
rect 13357 13311 13415 13317
rect 13357 13308 13369 13311
rect 12952 13280 13369 13308
rect 12952 13268 12958 13280
rect 13357 13277 13369 13280
rect 13403 13277 13415 13311
rect 13357 13271 13415 13277
rect 13630 13268 13636 13320
rect 13688 13268 13694 13320
rect 13817 13311 13875 13317
rect 13817 13277 13829 13311
rect 13863 13308 13875 13311
rect 13906 13308 13912 13320
rect 13863 13280 13912 13308
rect 13863 13277 13875 13280
rect 13817 13271 13875 13277
rect 13906 13268 13912 13280
rect 13964 13268 13970 13320
rect 15010 13268 15016 13320
rect 15068 13308 15074 13320
rect 15565 13311 15623 13317
rect 15565 13308 15577 13311
rect 15068 13280 15577 13308
rect 15068 13268 15074 13280
rect 15565 13277 15577 13280
rect 15611 13277 15623 13311
rect 15565 13271 15623 13277
rect 15930 13268 15936 13320
rect 15988 13308 15994 13320
rect 16592 13317 16620 13348
rect 16666 13336 16672 13388
rect 16724 13376 16730 13388
rect 17494 13376 17500 13388
rect 16724 13348 17500 13376
rect 16724 13336 16730 13348
rect 17494 13336 17500 13348
rect 17552 13336 17558 13388
rect 18322 13336 18328 13388
rect 18380 13336 18386 13388
rect 18414 13336 18420 13388
rect 18472 13376 18478 13388
rect 19702 13376 19708 13388
rect 18472 13348 19708 13376
rect 18472 13336 18478 13348
rect 19702 13336 19708 13348
rect 19760 13336 19766 13388
rect 20070 13336 20076 13388
rect 20128 13336 20134 13388
rect 21085 13379 21143 13385
rect 21085 13345 21097 13379
rect 21131 13376 21143 13379
rect 21450 13376 21456 13388
rect 21131 13348 21456 13376
rect 21131 13345 21143 13348
rect 21085 13339 21143 13345
rect 21450 13336 21456 13348
rect 21508 13336 21514 13388
rect 23216 13385 23244 13484
rect 23201 13379 23259 13385
rect 23201 13345 23213 13379
rect 23247 13345 23259 13379
rect 23201 13339 23259 13345
rect 16025 13311 16083 13317
rect 16025 13308 16037 13311
rect 15988 13280 16037 13308
rect 15988 13268 15994 13280
rect 16025 13277 16037 13280
rect 16071 13277 16083 13311
rect 16025 13271 16083 13277
rect 16301 13311 16359 13317
rect 16301 13277 16313 13311
rect 16347 13277 16359 13311
rect 16301 13271 16359 13277
rect 16577 13311 16635 13317
rect 16577 13277 16589 13311
rect 16623 13277 16635 13311
rect 16577 13271 16635 13277
rect 12986 13240 12992 13252
rect 12360 13212 12992 13240
rect 11885 13203 11943 13209
rect 12986 13200 12992 13212
rect 13044 13200 13050 13252
rect 13446 13200 13452 13252
rect 13504 13240 13510 13252
rect 16316 13240 16344 13271
rect 17954 13268 17960 13320
rect 18012 13268 18018 13320
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19521 13311 19579 13317
rect 19521 13308 19533 13311
rect 19392 13280 19533 13308
rect 19392 13268 19398 13280
rect 19521 13277 19533 13280
rect 19567 13277 19579 13311
rect 19521 13271 19579 13277
rect 20533 13311 20591 13317
rect 20533 13277 20545 13311
rect 20579 13308 20591 13311
rect 21361 13311 21419 13317
rect 21361 13308 21373 13311
rect 20579 13280 21373 13308
rect 20579 13277 20591 13280
rect 20533 13271 20591 13277
rect 21361 13277 21373 13280
rect 21407 13277 21419 13311
rect 21361 13271 21419 13277
rect 16758 13240 16764 13252
rect 13504 13212 15976 13240
rect 16316 13212 16764 13240
rect 13504 13200 13510 13212
rect 9232 13144 9536 13172
rect 10962 13132 10968 13184
rect 11020 13172 11026 13184
rect 11149 13175 11207 13181
rect 11149 13172 11161 13175
rect 11020 13144 11161 13172
rect 11020 13132 11026 13144
rect 11149 13141 11161 13144
rect 11195 13141 11207 13175
rect 11149 13135 11207 13141
rect 11514 13132 11520 13184
rect 11572 13132 11578 13184
rect 12066 13132 12072 13184
rect 12124 13172 12130 13184
rect 12161 13175 12219 13181
rect 12161 13172 12173 13175
rect 12124 13144 12173 13172
rect 12124 13132 12130 13144
rect 12161 13141 12173 13144
rect 12207 13141 12219 13175
rect 12161 13135 12219 13141
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 15013 13175 15071 13181
rect 15013 13172 15025 13175
rect 14700 13144 15025 13172
rect 14700 13132 14706 13144
rect 15013 13141 15025 13144
rect 15059 13141 15071 13175
rect 15948 13172 15976 13212
rect 16758 13200 16764 13212
rect 16816 13200 16822 13252
rect 18049 13243 18107 13249
rect 18049 13209 18061 13243
rect 18095 13240 18107 13243
rect 18506 13240 18512 13252
rect 18095 13212 18512 13240
rect 18095 13209 18107 13212
rect 18049 13203 18107 13209
rect 18506 13200 18512 13212
rect 18564 13200 18570 13252
rect 18874 13200 18880 13252
rect 18932 13200 18938 13252
rect 19978 13200 19984 13252
rect 20036 13200 20042 13252
rect 20548 13172 20576 13271
rect 22830 13268 22836 13320
rect 22888 13268 22894 13320
rect 23474 13268 23480 13320
rect 23532 13308 23538 13320
rect 23753 13311 23811 13317
rect 23753 13308 23765 13311
rect 23532 13280 23765 13308
rect 23532 13268 23538 13280
rect 23753 13277 23765 13280
rect 23799 13277 23811 13311
rect 23753 13271 23811 13277
rect 20714 13200 20720 13252
rect 20772 13240 20778 13252
rect 23014 13240 23020 13252
rect 20772 13212 23020 13240
rect 20772 13200 20778 13212
rect 23014 13200 23020 13212
rect 23072 13200 23078 13252
rect 23658 13200 23664 13252
rect 23716 13200 23722 13252
rect 15948 13144 20576 13172
rect 15013 13135 15071 13141
rect 21266 13132 21272 13184
rect 21324 13172 21330 13184
rect 22186 13172 22192 13184
rect 21324 13144 22192 13172
rect 21324 13132 21330 13144
rect 22186 13132 22192 13144
rect 22244 13132 22250 13184
rect 24118 13132 24124 13184
rect 24176 13132 24182 13184
rect 1104 13082 24840 13104
rect 1104 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 24214 13082
rect 24266 13030 24278 13082
rect 24330 13030 24342 13082
rect 24394 13030 24406 13082
rect 24458 13030 24470 13082
rect 24522 13030 24840 13082
rect 1104 13008 24840 13030
rect 1673 12971 1731 12977
rect 1673 12937 1685 12971
rect 1719 12968 1731 12971
rect 9766 12968 9772 12980
rect 1719 12940 9772 12968
rect 1719 12937 1731 12940
rect 1673 12931 1731 12937
rect 9766 12928 9772 12940
rect 9824 12928 9830 12980
rect 10594 12928 10600 12980
rect 10652 12968 10658 12980
rect 10965 12971 11023 12977
rect 10965 12968 10977 12971
rect 10652 12940 10977 12968
rect 10652 12928 10658 12940
rect 10965 12937 10977 12940
rect 11011 12937 11023 12971
rect 10965 12931 11023 12937
rect 11698 12928 11704 12980
rect 11756 12968 11762 12980
rect 11882 12968 11888 12980
rect 11756 12940 11888 12968
rect 11756 12928 11762 12940
rect 1854 12860 1860 12912
rect 1912 12900 1918 12912
rect 2041 12903 2099 12909
rect 2041 12900 2053 12903
rect 1912 12872 2053 12900
rect 1912 12860 1918 12872
rect 2041 12869 2053 12872
rect 2087 12869 2099 12903
rect 2041 12863 2099 12869
rect 2130 12860 2136 12912
rect 2188 12900 2194 12912
rect 2241 12903 2299 12909
rect 2241 12900 2253 12903
rect 2188 12872 2253 12900
rect 2188 12860 2194 12872
rect 2241 12869 2253 12872
rect 2287 12900 2299 12903
rect 3053 12903 3111 12909
rect 2287 12872 2774 12900
rect 2287 12869 2299 12872
rect 2241 12863 2299 12869
rect 1302 12792 1308 12844
rect 1360 12832 1366 12844
rect 1489 12835 1547 12841
rect 1489 12832 1501 12835
rect 1360 12804 1501 12832
rect 1360 12792 1366 12804
rect 1489 12801 1501 12804
rect 1535 12801 1547 12835
rect 2746 12832 2774 12872
rect 3053 12869 3065 12903
rect 3099 12900 3111 12903
rect 3234 12900 3240 12912
rect 3099 12872 3240 12900
rect 3099 12869 3111 12872
rect 3053 12863 3111 12869
rect 3234 12860 3240 12872
rect 3292 12860 3298 12912
rect 3865 12903 3923 12909
rect 3865 12869 3877 12903
rect 3911 12900 3923 12903
rect 3911 12872 4016 12900
rect 3911 12869 3923 12872
rect 3865 12863 3923 12869
rect 3988 12832 4016 12872
rect 4062 12860 4068 12912
rect 4120 12860 4126 12912
rect 5718 12860 5724 12912
rect 5776 12860 5782 12912
rect 5902 12860 5908 12912
rect 5960 12909 5966 12912
rect 5960 12903 5979 12909
rect 5967 12900 5979 12903
rect 6546 12900 6552 12912
rect 5967 12872 6552 12900
rect 5967 12869 5979 12872
rect 5960 12863 5979 12869
rect 5960 12860 5966 12863
rect 6546 12860 6552 12872
rect 6604 12860 6610 12912
rect 8570 12900 8576 12912
rect 7944 12872 8576 12900
rect 4614 12832 4620 12844
rect 2746 12804 4620 12832
rect 1489 12795 1547 12801
rect 4614 12792 4620 12804
rect 4672 12832 4678 12844
rect 5920 12832 5948 12860
rect 7944 12841 7972 12872
rect 8570 12860 8576 12872
rect 8628 12860 8634 12912
rect 9490 12860 9496 12912
rect 9548 12860 9554 12912
rect 10229 12903 10287 12909
rect 10229 12869 10241 12903
rect 10275 12900 10287 12903
rect 10318 12900 10324 12912
rect 10275 12872 10324 12900
rect 10275 12869 10287 12872
rect 10229 12863 10287 12869
rect 10318 12860 10324 12872
rect 10376 12860 10382 12912
rect 4672 12804 5948 12832
rect 7929 12835 7987 12841
rect 4672 12792 4678 12804
rect 7929 12801 7941 12835
rect 7975 12801 7987 12835
rect 7929 12795 7987 12801
rect 11606 12792 11612 12844
rect 11664 12792 11670 12844
rect 11698 12792 11704 12844
rect 11756 12792 11762 12844
rect 2222 12724 2228 12776
rect 2280 12764 2286 12776
rect 2280 12736 3096 12764
rect 2280 12724 2286 12736
rect 2409 12699 2467 12705
rect 2409 12665 2421 12699
rect 2455 12696 2467 12699
rect 2774 12696 2780 12708
rect 2455 12668 2780 12696
rect 2455 12665 2467 12668
rect 2409 12659 2467 12665
rect 2774 12656 2780 12668
rect 2832 12656 2838 12708
rect 3068 12696 3096 12736
rect 3142 12724 3148 12776
rect 3200 12724 3206 12776
rect 3329 12767 3387 12773
rect 3329 12733 3341 12767
rect 3375 12764 3387 12767
rect 3418 12764 3424 12776
rect 3375 12736 3424 12764
rect 3375 12733 3387 12736
rect 3329 12727 3387 12733
rect 3418 12724 3424 12736
rect 3476 12724 3482 12776
rect 7098 12724 7104 12776
rect 7156 12764 7162 12776
rect 8205 12767 8263 12773
rect 8205 12764 8217 12767
rect 7156 12736 8217 12764
rect 7156 12724 7162 12736
rect 8205 12733 8217 12736
rect 8251 12733 8263 12767
rect 8205 12727 8263 12733
rect 8481 12767 8539 12773
rect 8481 12733 8493 12767
rect 8527 12764 8539 12767
rect 9490 12764 9496 12776
rect 8527 12736 9496 12764
rect 8527 12733 8539 12736
rect 8481 12727 8539 12733
rect 9490 12724 9496 12736
rect 9548 12724 9554 12776
rect 10505 12767 10563 12773
rect 10505 12733 10517 12767
rect 10551 12733 10563 12767
rect 10505 12727 10563 12733
rect 6730 12696 6736 12708
rect 3068 12668 3924 12696
rect 2222 12588 2228 12640
rect 2280 12588 2286 12640
rect 2314 12588 2320 12640
rect 2372 12628 2378 12640
rect 2685 12631 2743 12637
rect 2685 12628 2697 12631
rect 2372 12600 2697 12628
rect 2372 12588 2378 12600
rect 2685 12597 2697 12600
rect 2731 12597 2743 12631
rect 2685 12591 2743 12597
rect 3694 12588 3700 12640
rect 3752 12588 3758 12640
rect 3896 12637 3924 12668
rect 5920 12668 6736 12696
rect 3881 12631 3939 12637
rect 3881 12597 3893 12631
rect 3927 12628 3939 12631
rect 4706 12628 4712 12640
rect 3927 12600 4712 12628
rect 3927 12597 3939 12600
rect 3881 12591 3939 12597
rect 4706 12588 4712 12600
rect 4764 12628 4770 12640
rect 5810 12628 5816 12640
rect 4764 12600 5816 12628
rect 4764 12588 4770 12600
rect 5810 12588 5816 12600
rect 5868 12628 5874 12640
rect 5920 12637 5948 12668
rect 6730 12656 6736 12668
rect 6788 12656 6794 12708
rect 5905 12631 5963 12637
rect 5905 12628 5917 12631
rect 5868 12600 5917 12628
rect 5868 12588 5874 12600
rect 5905 12597 5917 12600
rect 5951 12597 5963 12631
rect 5905 12591 5963 12597
rect 6089 12631 6147 12637
rect 6089 12597 6101 12631
rect 6135 12628 6147 12631
rect 6178 12628 6184 12640
rect 6135 12600 6184 12628
rect 6135 12597 6147 12600
rect 6089 12591 6147 12597
rect 6178 12588 6184 12600
rect 6236 12588 6242 12640
rect 7745 12631 7803 12637
rect 7745 12597 7757 12631
rect 7791 12628 7803 12631
rect 8662 12628 8668 12640
rect 7791 12600 8668 12628
rect 7791 12597 7803 12600
rect 7745 12591 7803 12597
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 8938 12588 8944 12640
rect 8996 12628 9002 12640
rect 10520 12628 10548 12727
rect 11330 12724 11336 12776
rect 11388 12764 11394 12776
rect 11808 12764 11836 12940
rect 11882 12928 11888 12940
rect 11940 12928 11946 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12621 12971 12679 12977
rect 12621 12968 12633 12971
rect 12124 12940 12633 12968
rect 12124 12928 12130 12940
rect 12621 12937 12633 12940
rect 12667 12937 12679 12971
rect 13906 12968 13912 12980
rect 12621 12931 12679 12937
rect 12912 12940 13912 12968
rect 11974 12860 11980 12912
rect 12032 12900 12038 12912
rect 12912 12900 12940 12940
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 15930 12968 15936 12980
rect 15580 12940 15936 12968
rect 15381 12903 15439 12909
rect 15381 12900 15393 12903
rect 12032 12872 12940 12900
rect 12032 12860 12038 12872
rect 11882 12792 11888 12844
rect 11940 12792 11946 12844
rect 12066 12792 12072 12844
rect 12124 12792 12130 12844
rect 12912 12841 12940 12872
rect 13372 12872 15393 12900
rect 12805 12835 12863 12841
rect 12805 12832 12817 12835
rect 12544 12804 12817 12832
rect 12544 12764 12572 12804
rect 12805 12801 12817 12804
rect 12851 12801 12863 12835
rect 12805 12795 12863 12801
rect 12897 12835 12955 12841
rect 12897 12801 12909 12835
rect 12943 12801 12955 12835
rect 12897 12795 12955 12801
rect 12986 12792 12992 12844
rect 13044 12832 13050 12844
rect 13262 12832 13268 12844
rect 13044 12804 13268 12832
rect 13044 12792 13050 12804
rect 13262 12792 13268 12804
rect 13320 12832 13326 12844
rect 13372 12832 13400 12872
rect 15381 12869 15393 12872
rect 15427 12869 15439 12903
rect 15381 12863 15439 12869
rect 13320 12804 13400 12832
rect 14001 12835 14059 12841
rect 13320 12792 13326 12804
rect 14001 12801 14013 12835
rect 14047 12832 14059 12835
rect 14047 12804 14412 12832
rect 14047 12801 14059 12804
rect 14001 12795 14059 12801
rect 11388 12736 12572 12764
rect 11388 12724 11394 12736
rect 12618 12724 12624 12776
rect 12676 12764 12682 12776
rect 13081 12767 13139 12773
rect 13081 12764 13093 12767
rect 12676 12736 13093 12764
rect 12676 12724 12682 12736
rect 13081 12733 13093 12736
rect 13127 12733 13139 12767
rect 13081 12727 13139 12733
rect 11790 12656 11796 12708
rect 11848 12696 11854 12708
rect 14016 12696 14044 12795
rect 14090 12724 14096 12776
rect 14148 12724 14154 12776
rect 14384 12764 14412 12804
rect 14642 12792 14648 12844
rect 14700 12792 14706 12844
rect 14737 12835 14795 12841
rect 14737 12801 14749 12835
rect 14783 12832 14795 12835
rect 14826 12832 14832 12844
rect 14783 12804 14832 12832
rect 14783 12801 14795 12804
rect 14737 12795 14795 12801
rect 14826 12792 14832 12804
rect 14884 12792 14890 12844
rect 14918 12792 14924 12844
rect 14976 12792 14982 12844
rect 15580 12841 15608 12940
rect 15930 12928 15936 12940
rect 15988 12928 15994 12980
rect 16758 12928 16764 12980
rect 16816 12968 16822 12980
rect 18509 12971 18567 12977
rect 18509 12968 18521 12971
rect 16816 12940 18521 12968
rect 16816 12928 16822 12940
rect 18509 12937 18521 12940
rect 18555 12968 18567 12971
rect 20990 12968 20996 12980
rect 18555 12940 20996 12968
rect 18555 12937 18567 12940
rect 18509 12931 18567 12937
rect 20990 12928 20996 12940
rect 21048 12928 21054 12980
rect 21542 12928 21548 12980
rect 21600 12968 21606 12980
rect 21600 12940 24256 12968
rect 21600 12928 21606 12940
rect 16666 12900 16672 12912
rect 15764 12872 16672 12900
rect 15764 12841 15792 12872
rect 16666 12860 16672 12872
rect 16724 12860 16730 12912
rect 16942 12900 16948 12912
rect 16776 12872 16948 12900
rect 15565 12835 15623 12841
rect 15565 12801 15577 12835
rect 15611 12801 15623 12835
rect 15565 12795 15623 12801
rect 15749 12835 15807 12841
rect 15749 12801 15761 12835
rect 15795 12801 15807 12835
rect 15749 12795 15807 12801
rect 15580 12764 15608 12795
rect 16114 12792 16120 12844
rect 16172 12832 16178 12844
rect 16776 12841 16804 12872
rect 16942 12860 16948 12872
rect 17000 12860 17006 12912
rect 18046 12860 18052 12912
rect 18104 12860 18110 12912
rect 21450 12860 21456 12912
rect 21508 12900 21514 12912
rect 24228 12909 24256 12940
rect 24213 12903 24271 12909
rect 21508 12872 23704 12900
rect 21508 12860 21514 12872
rect 16393 12835 16451 12841
rect 16393 12832 16405 12835
rect 16172 12804 16405 12832
rect 16172 12792 16178 12804
rect 16393 12801 16405 12804
rect 16439 12801 16451 12835
rect 16393 12795 16451 12801
rect 16761 12835 16819 12841
rect 16761 12801 16773 12835
rect 16807 12801 16819 12835
rect 16761 12795 16819 12801
rect 18877 12835 18935 12841
rect 18877 12801 18889 12835
rect 18923 12801 18935 12835
rect 18877 12795 18935 12801
rect 20349 12835 20407 12841
rect 20349 12801 20361 12835
rect 20395 12832 20407 12835
rect 20622 12832 20628 12844
rect 20395 12804 20628 12832
rect 20395 12801 20407 12804
rect 20349 12795 20407 12801
rect 15654 12764 15660 12776
rect 14384 12736 15660 12764
rect 15654 12724 15660 12736
rect 15712 12724 15718 12776
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 16209 12767 16267 12773
rect 16209 12764 16221 12767
rect 15896 12736 16221 12764
rect 15896 12724 15902 12736
rect 16209 12733 16221 12736
rect 16255 12733 16267 12767
rect 17037 12767 17095 12773
rect 17037 12764 17049 12767
rect 16209 12727 16267 12733
rect 16868 12736 17049 12764
rect 11848 12668 14044 12696
rect 11848 12656 11854 12668
rect 15746 12656 15752 12708
rect 15804 12696 15810 12708
rect 16025 12699 16083 12705
rect 16025 12696 16037 12699
rect 15804 12668 16037 12696
rect 15804 12656 15810 12668
rect 16025 12665 16037 12668
rect 16071 12665 16083 12699
rect 16301 12699 16359 12705
rect 16301 12696 16313 12699
rect 16025 12659 16083 12665
rect 16132 12668 16313 12696
rect 8996 12600 10548 12628
rect 14369 12631 14427 12637
rect 8996 12588 9002 12600
rect 14369 12597 14381 12631
rect 14415 12628 14427 12631
rect 14918 12628 14924 12640
rect 14415 12600 14924 12628
rect 14415 12597 14427 12600
rect 14369 12591 14427 12597
rect 14918 12588 14924 12600
rect 14976 12588 14982 12640
rect 15102 12588 15108 12640
rect 15160 12588 15166 12640
rect 15930 12588 15936 12640
rect 15988 12628 15994 12640
rect 16132 12628 16160 12668
rect 16301 12665 16313 12668
rect 16347 12665 16359 12699
rect 16301 12659 16359 12665
rect 15988 12600 16160 12628
rect 16209 12631 16267 12637
rect 15988 12588 15994 12600
rect 16209 12597 16221 12631
rect 16255 12628 16267 12631
rect 16868 12628 16896 12736
rect 17037 12733 17049 12736
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 17770 12724 17776 12776
rect 17828 12764 17834 12776
rect 18892 12764 18920 12795
rect 20622 12792 20628 12804
rect 20680 12792 20686 12844
rect 21082 12792 21088 12844
rect 21140 12832 21146 12844
rect 21634 12832 21640 12844
rect 21140 12804 21640 12832
rect 21140 12792 21146 12804
rect 21634 12792 21640 12804
rect 21692 12792 21698 12844
rect 21928 12841 21956 12872
rect 21913 12835 21971 12841
rect 21913 12801 21925 12835
rect 21959 12832 21971 12835
rect 21959 12804 21993 12832
rect 21959 12801 21971 12804
rect 21913 12795 21971 12801
rect 22094 12792 22100 12844
rect 22152 12832 22158 12844
rect 22557 12835 22615 12841
rect 22557 12832 22569 12835
rect 22152 12804 22569 12832
rect 22152 12792 22158 12804
rect 22557 12801 22569 12804
rect 22603 12801 22615 12835
rect 22557 12795 22615 12801
rect 20717 12767 20775 12773
rect 20717 12764 20729 12767
rect 17828 12736 20729 12764
rect 17828 12724 17834 12736
rect 20717 12733 20729 12736
rect 20763 12733 20775 12767
rect 20717 12727 20775 12733
rect 21266 12724 21272 12776
rect 21324 12724 21330 12776
rect 20349 12699 20407 12705
rect 20349 12665 20361 12699
rect 20395 12696 20407 12699
rect 21177 12699 21235 12705
rect 21177 12696 21189 12699
rect 20395 12668 21189 12696
rect 20395 12665 20407 12668
rect 20349 12659 20407 12665
rect 21177 12665 21189 12668
rect 21223 12696 21235 12699
rect 21358 12696 21364 12708
rect 21223 12668 21364 12696
rect 21223 12665 21235 12668
rect 21177 12659 21235 12665
rect 21358 12656 21364 12668
rect 21416 12656 21422 12708
rect 22572 12696 22600 12795
rect 22830 12792 22836 12844
rect 22888 12792 22894 12844
rect 23676 12841 23704 12872
rect 24213 12869 24225 12903
rect 24259 12869 24271 12903
rect 24213 12863 24271 12869
rect 23661 12835 23719 12841
rect 23661 12801 23673 12835
rect 23707 12801 23719 12835
rect 23661 12795 23719 12801
rect 23937 12835 23995 12841
rect 23937 12801 23949 12835
rect 23983 12801 23995 12835
rect 23937 12795 23995 12801
rect 23106 12724 23112 12776
rect 23164 12724 23170 12776
rect 23201 12699 23259 12705
rect 23201 12696 23213 12699
rect 22572 12668 23213 12696
rect 23201 12665 23213 12668
rect 23247 12665 23259 12699
rect 23201 12659 23259 12665
rect 16255 12600 16896 12628
rect 16255 12597 16267 12600
rect 16209 12591 16267 12597
rect 19794 12588 19800 12640
rect 19852 12628 19858 12640
rect 23952 12628 23980 12795
rect 19852 12600 23980 12628
rect 19852 12588 19858 12600
rect 1104 12538 24840 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 12214 12538
rect 12266 12486 12278 12538
rect 12330 12486 12342 12538
rect 12394 12486 12406 12538
rect 12458 12486 12470 12538
rect 12522 12486 20214 12538
rect 20266 12486 20278 12538
rect 20330 12486 20342 12538
rect 20394 12486 20406 12538
rect 20458 12486 20470 12538
rect 20522 12486 24840 12538
rect 1104 12464 24840 12486
rect 4890 12424 4896 12436
rect 4356 12396 4896 12424
rect 1765 12291 1823 12297
rect 1765 12257 1777 12291
rect 1811 12288 1823 12291
rect 2314 12288 2320 12300
rect 1811 12260 2320 12288
rect 1811 12257 1823 12260
rect 1765 12251 1823 12257
rect 2314 12248 2320 12260
rect 2372 12248 2378 12300
rect 4356 12297 4384 12396
rect 4890 12384 4896 12396
rect 4948 12424 4954 12436
rect 4948 12396 7328 12424
rect 4948 12384 4954 12396
rect 4341 12291 4399 12297
rect 4341 12257 4353 12291
rect 4387 12257 4399 12291
rect 4341 12251 4399 12257
rect 4433 12291 4491 12297
rect 4433 12257 4445 12291
rect 4479 12257 4491 12291
rect 4433 12251 4491 12257
rect 4893 12291 4951 12297
rect 4893 12257 4905 12291
rect 4939 12288 4951 12291
rect 7098 12288 7104 12300
rect 4939 12260 7104 12288
rect 4939 12257 4951 12260
rect 4893 12251 4951 12257
rect 1486 12180 1492 12232
rect 1544 12180 1550 12232
rect 3142 12180 3148 12232
rect 3200 12220 3206 12232
rect 4062 12220 4068 12232
rect 3200 12192 4068 12220
rect 3200 12180 3206 12192
rect 4062 12180 4068 12192
rect 4120 12220 4126 12232
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 4120 12192 4261 12220
rect 4120 12180 4126 12192
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 2774 12112 2780 12164
rect 2832 12112 2838 12164
rect 3418 12112 3424 12164
rect 3476 12152 3482 12164
rect 4448 12152 4476 12251
rect 7098 12248 7104 12260
rect 7156 12248 7162 12300
rect 7300 12229 7328 12396
rect 9490 12384 9496 12436
rect 9548 12424 9554 12436
rect 9585 12427 9643 12433
rect 9585 12424 9597 12427
rect 9548 12396 9597 12424
rect 9548 12384 9554 12396
rect 9585 12393 9597 12396
rect 9631 12393 9643 12427
rect 9585 12387 9643 12393
rect 11974 12384 11980 12436
rect 12032 12424 12038 12436
rect 15381 12427 15439 12433
rect 12032 12396 15240 12424
rect 12032 12384 12038 12396
rect 13998 12356 14004 12368
rect 13280 12328 14004 12356
rect 7466 12248 7472 12300
rect 7524 12288 7530 12300
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 7524 12260 8125 12288
rect 7524 12248 7530 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10962 12288 10968 12300
rect 10091 12260 10968 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10962 12248 10968 12260
rect 11020 12248 11026 12300
rect 11149 12291 11207 12297
rect 11149 12257 11161 12291
rect 11195 12288 11207 12291
rect 11422 12288 11428 12300
rect 11195 12260 11428 12288
rect 11195 12257 11207 12260
rect 11149 12251 11207 12257
rect 11422 12248 11428 12260
rect 11480 12288 11486 12300
rect 12894 12288 12900 12300
rect 11480 12260 12900 12288
rect 11480 12248 11486 12260
rect 11060 12232 11112 12238
rect 7285 12223 7343 12229
rect 7285 12189 7297 12223
rect 7331 12189 7343 12223
rect 7285 12183 7343 12189
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8662 12220 8668 12232
rect 8435 12192 8668 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8662 12180 8668 12192
rect 8720 12180 8726 12232
rect 9766 12180 9772 12232
rect 9824 12220 9830 12232
rect 9861 12223 9919 12229
rect 9861 12220 9873 12223
rect 9824 12192 9873 12220
rect 9824 12180 9830 12192
rect 9861 12189 9873 12192
rect 9907 12189 9919 12223
rect 9861 12183 9919 12189
rect 9950 12180 9956 12232
rect 10008 12220 10014 12232
rect 10321 12223 10379 12229
rect 10321 12220 10333 12223
rect 10008 12192 10333 12220
rect 10008 12180 10014 12192
rect 10321 12189 10333 12192
rect 10367 12189 10379 12223
rect 10321 12183 10379 12189
rect 11238 12222 11244 12232
rect 11112 12194 11244 12222
rect 11238 12180 11244 12194
rect 11296 12180 11302 12232
rect 11882 12180 11888 12232
rect 11940 12220 11946 12232
rect 11977 12223 12035 12229
rect 11977 12220 11989 12223
rect 11940 12192 11989 12220
rect 11940 12180 11946 12192
rect 11977 12189 11989 12192
rect 12023 12189 12035 12223
rect 11977 12183 12035 12189
rect 12066 12180 12072 12232
rect 12124 12220 12130 12232
rect 12544 12229 12572 12260
rect 12894 12248 12900 12260
rect 12952 12248 12958 12300
rect 13280 12297 13308 12328
rect 13998 12316 14004 12328
rect 14056 12316 14062 12368
rect 13265 12291 13323 12297
rect 13265 12257 13277 12291
rect 13311 12257 13323 12291
rect 13265 12251 13323 12257
rect 13357 12291 13415 12297
rect 13357 12257 13369 12291
rect 13403 12288 13415 12291
rect 14826 12288 14832 12300
rect 13403 12260 14832 12288
rect 13403 12257 13415 12260
rect 13357 12251 13415 12257
rect 12253 12223 12311 12229
rect 12253 12220 12265 12223
rect 12124 12192 12265 12220
rect 12124 12180 12130 12192
rect 12253 12189 12265 12192
rect 12299 12189 12311 12223
rect 12253 12183 12311 12189
rect 12529 12223 12587 12229
rect 12529 12189 12541 12223
rect 12575 12189 12587 12223
rect 12529 12183 12587 12189
rect 12618 12180 12624 12232
rect 12676 12180 12682 12232
rect 12802 12180 12808 12232
rect 12860 12220 12866 12232
rect 13372 12220 13400 12251
rect 14826 12248 14832 12260
rect 14884 12248 14890 12300
rect 12860 12192 13400 12220
rect 12860 12180 12866 12192
rect 13446 12180 13452 12232
rect 13504 12180 13510 12232
rect 13538 12180 13544 12232
rect 13596 12180 13602 12232
rect 14642 12180 14648 12232
rect 14700 12220 14706 12232
rect 14737 12223 14795 12229
rect 14737 12220 14749 12223
rect 14700 12192 14749 12220
rect 14700 12180 14706 12192
rect 14737 12189 14749 12192
rect 14783 12189 14795 12223
rect 14737 12183 14795 12189
rect 14918 12180 14924 12232
rect 14976 12180 14982 12232
rect 15010 12180 15016 12232
rect 15068 12180 15074 12232
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12189 15163 12223
rect 15105 12183 15163 12189
rect 11060 12174 11112 12180
rect 3476 12124 4476 12152
rect 3476 12112 3482 12124
rect 3234 12044 3240 12096
rect 3292 12044 3298 12096
rect 3878 12044 3884 12096
rect 3936 12044 3942 12096
rect 4448 12084 4476 12124
rect 5166 12112 5172 12164
rect 5224 12112 5230 12164
rect 6178 12112 6184 12164
rect 6236 12112 6242 12164
rect 7377 12155 7435 12161
rect 7377 12152 7389 12155
rect 6656 12124 7389 12152
rect 5534 12084 5540 12096
rect 4448 12056 5540 12084
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 5810 12044 5816 12096
rect 5868 12084 5874 12096
rect 6656 12093 6684 12124
rect 7377 12121 7389 12124
rect 7423 12121 7435 12155
rect 7377 12115 7435 12121
rect 9490 12112 9496 12164
rect 9548 12112 9554 12164
rect 10134 12112 10140 12164
rect 10192 12152 10198 12164
rect 10410 12152 10416 12164
rect 10192 12124 10416 12152
rect 10192 12112 10198 12124
rect 10410 12112 10416 12124
rect 10468 12112 10474 12164
rect 10594 12112 10600 12164
rect 10652 12112 10658 12164
rect 12437 12155 12495 12161
rect 12437 12121 12449 12155
rect 12483 12152 12495 12155
rect 13262 12152 13268 12164
rect 12483 12124 13268 12152
rect 12483 12121 12495 12124
rect 12437 12115 12495 12121
rect 13262 12112 13268 12124
rect 13320 12112 13326 12164
rect 14826 12112 14832 12164
rect 14884 12152 14890 12164
rect 15120 12152 15148 12183
rect 14884 12124 15148 12152
rect 15212 12152 15240 12396
rect 15381 12393 15393 12427
rect 15427 12424 15439 12427
rect 15746 12424 15752 12436
rect 15427 12396 15752 12424
rect 15427 12393 15439 12396
rect 15381 12387 15439 12393
rect 15746 12384 15752 12396
rect 15804 12384 15810 12436
rect 15838 12384 15844 12436
rect 15896 12384 15902 12436
rect 16114 12384 16120 12436
rect 16172 12424 16178 12436
rect 16301 12427 16359 12433
rect 16301 12424 16313 12427
rect 16172 12396 16313 12424
rect 16172 12384 16178 12396
rect 16301 12393 16313 12396
rect 16347 12393 16359 12427
rect 16301 12387 16359 12393
rect 17129 12427 17187 12433
rect 17129 12393 17141 12427
rect 17175 12424 17187 12427
rect 17586 12424 17592 12436
rect 17175 12396 17592 12424
rect 17175 12393 17187 12396
rect 17129 12387 17187 12393
rect 17586 12384 17592 12396
rect 17644 12424 17650 12436
rect 17773 12427 17831 12433
rect 17773 12424 17785 12427
rect 17644 12396 17785 12424
rect 17644 12384 17650 12396
rect 17773 12393 17785 12396
rect 17819 12393 17831 12427
rect 17773 12387 17831 12393
rect 21450 12384 21456 12436
rect 21508 12384 21514 12436
rect 17313 12359 17371 12365
rect 17313 12325 17325 12359
rect 17359 12356 17371 12359
rect 18046 12356 18052 12368
rect 17359 12328 18052 12356
rect 17359 12325 17371 12328
rect 17313 12319 17371 12325
rect 18046 12316 18052 12328
rect 18104 12316 18110 12368
rect 20070 12316 20076 12368
rect 20128 12356 20134 12368
rect 20128 12328 21312 12356
rect 20128 12316 20134 12328
rect 15930 12248 15936 12300
rect 15988 12248 15994 12300
rect 16114 12248 16120 12300
rect 16172 12288 16178 12300
rect 17126 12288 17132 12300
rect 16172 12260 17132 12288
rect 16172 12248 16178 12260
rect 17126 12248 17132 12260
rect 17184 12248 17190 12300
rect 17678 12248 17684 12300
rect 17736 12288 17742 12300
rect 18601 12291 18659 12297
rect 18601 12288 18613 12291
rect 17736 12260 18613 12288
rect 17736 12248 17742 12260
rect 18601 12257 18613 12260
rect 18647 12257 18659 12291
rect 18601 12251 18659 12257
rect 15286 12180 15292 12232
rect 15344 12220 15350 12232
rect 15657 12223 15715 12229
rect 15657 12220 15669 12223
rect 15344 12192 15669 12220
rect 15344 12180 15350 12192
rect 15657 12189 15669 12192
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 15746 12180 15752 12232
rect 15804 12180 15810 12232
rect 16022 12180 16028 12232
rect 16080 12220 16086 12232
rect 16393 12223 16451 12229
rect 16393 12220 16405 12223
rect 16080 12192 16405 12220
rect 16080 12180 16086 12192
rect 16393 12189 16405 12192
rect 16439 12189 16451 12223
rect 17218 12220 17224 12232
rect 16393 12183 16451 12189
rect 16500 12192 17224 12220
rect 16500 12152 16528 12192
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 18322 12180 18328 12232
rect 18380 12180 18386 12232
rect 15212 12124 16528 12152
rect 16945 12155 17003 12161
rect 14884 12112 14890 12124
rect 6641 12087 6699 12093
rect 6641 12084 6653 12087
rect 5868 12056 6653 12084
rect 5868 12044 5874 12056
rect 6641 12053 6653 12056
rect 6687 12053 6699 12087
rect 6641 12047 6699 12053
rect 6914 12044 6920 12096
rect 6972 12044 6978 12096
rect 8570 12044 8576 12096
rect 8628 12084 8634 12096
rect 10226 12084 10232 12096
rect 8628 12056 10232 12084
rect 8628 12044 8634 12056
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 10318 12044 10324 12096
rect 10376 12044 10382 12096
rect 10962 12044 10968 12096
rect 11020 12084 11026 12096
rect 12066 12084 12072 12096
rect 11020 12056 12072 12084
rect 11020 12044 11026 12056
rect 12066 12044 12072 12056
rect 12124 12044 12130 12096
rect 12802 12044 12808 12096
rect 12860 12044 12866 12096
rect 13722 12044 13728 12096
rect 13780 12044 13786 12096
rect 14090 12044 14096 12096
rect 14148 12084 14154 12096
rect 15010 12084 15016 12096
rect 14148 12056 15016 12084
rect 14148 12044 14154 12056
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15120 12084 15148 12124
rect 16945 12121 16957 12155
rect 16991 12152 17003 12155
rect 17494 12152 17500 12164
rect 16991 12124 17500 12152
rect 16991 12121 17003 12124
rect 16945 12115 17003 12121
rect 17494 12112 17500 12124
rect 17552 12152 17558 12164
rect 17589 12155 17647 12161
rect 17589 12152 17601 12155
rect 17552 12124 17601 12152
rect 17552 12112 17558 12124
rect 17589 12121 17601 12124
rect 17635 12121 17647 12155
rect 18616 12152 18644 12251
rect 19794 12248 19800 12300
rect 19852 12288 19858 12300
rect 21284 12297 21312 12328
rect 23658 12316 23664 12368
rect 23716 12356 23722 12368
rect 23753 12359 23811 12365
rect 23753 12356 23765 12359
rect 23716 12328 23765 12356
rect 23716 12316 23722 12328
rect 23753 12325 23765 12328
rect 23799 12325 23811 12359
rect 23753 12319 23811 12325
rect 21177 12291 21235 12297
rect 21177 12288 21189 12291
rect 19852 12260 21189 12288
rect 19852 12248 19858 12260
rect 19334 12180 19340 12232
rect 19392 12180 19398 12232
rect 19978 12180 19984 12232
rect 20036 12180 20042 12232
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12220 20315 12223
rect 20622 12220 20628 12232
rect 20303 12192 20628 12220
rect 20303 12189 20315 12192
rect 20257 12183 20315 12189
rect 20622 12180 20628 12192
rect 20680 12180 20686 12232
rect 19426 12152 19432 12164
rect 18616 12124 19432 12152
rect 17589 12115 17647 12121
rect 19426 12112 19432 12124
rect 19484 12112 19490 12164
rect 15838 12084 15844 12096
rect 15120 12056 15844 12084
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 17155 12087 17213 12093
rect 17155 12053 17167 12087
rect 17201 12084 17213 12087
rect 17678 12084 17684 12096
rect 17201 12056 17684 12084
rect 17201 12053 17213 12056
rect 17155 12047 17213 12053
rect 17678 12044 17684 12056
rect 17736 12084 17742 12096
rect 17789 12087 17847 12093
rect 17789 12084 17801 12087
rect 17736 12056 17801 12084
rect 17736 12044 17742 12056
rect 17789 12053 17801 12056
rect 17835 12053 17847 12087
rect 17789 12047 17847 12053
rect 17954 12044 17960 12096
rect 18012 12044 18018 12096
rect 20622 12044 20628 12096
rect 20680 12084 20686 12096
rect 20732 12084 20760 12260
rect 21177 12257 21189 12260
rect 21223 12257 21235 12291
rect 21177 12251 21235 12257
rect 21269 12291 21327 12297
rect 21269 12257 21281 12291
rect 21315 12288 21327 12291
rect 22094 12288 22100 12300
rect 21315 12260 22100 12288
rect 21315 12257 21327 12260
rect 21269 12251 21327 12257
rect 22094 12248 22100 12260
rect 22152 12248 22158 12300
rect 20990 12180 20996 12232
rect 21048 12180 21054 12232
rect 21082 12180 21088 12232
rect 21140 12180 21146 12232
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 21729 12223 21787 12229
rect 21729 12220 21741 12223
rect 21508 12192 21741 12220
rect 21508 12180 21514 12192
rect 21729 12189 21741 12192
rect 21775 12189 21787 12223
rect 21729 12183 21787 12189
rect 21910 12180 21916 12232
rect 21968 12180 21974 12232
rect 22462 12180 22468 12232
rect 22520 12180 22526 12232
rect 23842 12180 23848 12232
rect 23900 12180 23906 12232
rect 20680 12056 20760 12084
rect 20680 12044 20686 12056
rect 1104 11994 24840 12016
rect 1104 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 24214 11994
rect 24266 11942 24278 11994
rect 24330 11942 24342 11994
rect 24394 11942 24406 11994
rect 24458 11942 24470 11994
rect 24522 11942 24840 11994
rect 1104 11920 24840 11942
rect 3878 11880 3884 11892
rect 2746 11852 3884 11880
rect 2593 11815 2651 11821
rect 2593 11781 2605 11815
rect 2639 11812 2651 11815
rect 2746 11812 2774 11852
rect 3878 11840 3884 11852
rect 3936 11840 3942 11892
rect 4062 11840 4068 11892
rect 4120 11840 4126 11892
rect 4614 11840 4620 11892
rect 4672 11880 4678 11892
rect 4985 11883 5043 11889
rect 4985 11880 4997 11883
rect 4672 11852 4997 11880
rect 4672 11840 4678 11852
rect 4985 11849 4997 11852
rect 5031 11849 5043 11883
rect 4985 11843 5043 11849
rect 5166 11840 5172 11892
rect 5224 11880 5230 11892
rect 5353 11883 5411 11889
rect 5353 11880 5365 11883
rect 5224 11852 5365 11880
rect 5224 11840 5230 11852
rect 5353 11849 5365 11852
rect 5399 11849 5411 11883
rect 5353 11843 5411 11849
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 5810 11880 5816 11892
rect 5767 11852 5816 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 5810 11840 5816 11852
rect 5868 11840 5874 11892
rect 6638 11889 6644 11892
rect 6625 11883 6644 11889
rect 6625 11849 6637 11883
rect 6625 11843 6644 11849
rect 6638 11840 6644 11843
rect 6696 11840 6702 11892
rect 7466 11880 7472 11892
rect 6748 11852 7472 11880
rect 2639 11784 2774 11812
rect 2639 11781 2651 11784
rect 2593 11775 2651 11781
rect 5534 11772 5540 11824
rect 5592 11812 5598 11824
rect 6748 11812 6776 11852
rect 7466 11840 7472 11852
rect 7524 11840 7530 11892
rect 9490 11840 9496 11892
rect 9548 11880 9554 11892
rect 10505 11883 10563 11889
rect 10505 11880 10517 11883
rect 9548 11852 10517 11880
rect 9548 11840 9554 11852
rect 10505 11849 10517 11852
rect 10551 11849 10563 11883
rect 10505 11843 10563 11849
rect 10594 11840 10600 11892
rect 10652 11880 10658 11892
rect 11698 11880 11704 11892
rect 10652 11852 11704 11880
rect 10652 11840 10658 11852
rect 11698 11840 11704 11852
rect 11756 11880 11762 11892
rect 11756 11852 12434 11880
rect 11756 11840 11762 11852
rect 5592 11784 6776 11812
rect 6825 11815 6883 11821
rect 5592 11772 5598 11784
rect 1302 11704 1308 11756
rect 1360 11744 1366 11756
rect 1489 11747 1547 11753
rect 1489 11744 1501 11747
rect 1360 11716 1501 11744
rect 1360 11704 1366 11716
rect 1489 11713 1501 11716
rect 1535 11744 1547 11747
rect 1949 11747 2007 11753
rect 1949 11744 1961 11747
rect 1535 11716 1961 11744
rect 1535 11713 1547 11716
rect 1489 11707 1547 11713
rect 1949 11713 1961 11716
rect 1995 11713 2007 11747
rect 1949 11707 2007 11713
rect 3694 11704 3700 11756
rect 3752 11704 3758 11756
rect 4801 11747 4859 11753
rect 4801 11713 4813 11747
rect 4847 11744 4859 11747
rect 5626 11744 5632 11756
rect 4847 11716 5632 11744
rect 4847 11713 4859 11716
rect 4801 11707 4859 11713
rect 5626 11704 5632 11716
rect 5684 11704 5690 11756
rect 2317 11679 2375 11685
rect 2317 11676 2329 11679
rect 1504 11648 2329 11676
rect 1504 11620 1532 11648
rect 2317 11645 2329 11648
rect 2363 11645 2375 11679
rect 2317 11639 2375 11645
rect 2424 11648 5764 11676
rect 1486 11568 1492 11620
rect 1544 11568 1550 11620
rect 1673 11611 1731 11617
rect 1673 11577 1685 11611
rect 1719 11608 1731 11611
rect 2424 11608 2452 11648
rect 1719 11580 2452 11608
rect 5736 11608 5764 11648
rect 5810 11636 5816 11688
rect 5868 11636 5874 11688
rect 5920 11685 5948 11784
rect 6825 11781 6837 11815
rect 6871 11781 6883 11815
rect 6825 11775 6883 11781
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6840 11744 6868 11775
rect 7374 11772 7380 11824
rect 7432 11772 7438 11824
rect 9122 11812 9128 11824
rect 8602 11784 9128 11812
rect 9122 11772 9128 11784
rect 9180 11772 9186 11824
rect 9950 11772 9956 11824
rect 10008 11772 10014 11824
rect 10045 11815 10103 11821
rect 10045 11781 10057 11815
rect 10091 11812 10103 11815
rect 10686 11812 10692 11824
rect 10091 11784 10692 11812
rect 10091 11781 10103 11784
rect 10045 11775 10103 11781
rect 10686 11772 10692 11784
rect 10744 11772 10750 11824
rect 6052 11716 6868 11744
rect 9677 11747 9735 11753
rect 6052 11704 6058 11716
rect 9677 11713 9689 11747
rect 9723 11713 9735 11747
rect 9677 11707 9735 11713
rect 5905 11679 5963 11685
rect 5905 11645 5917 11679
rect 5951 11645 5963 11679
rect 5905 11639 5963 11645
rect 6638 11636 6644 11688
rect 6696 11676 6702 11688
rect 7098 11676 7104 11688
rect 6696 11648 7104 11676
rect 6696 11636 6702 11648
rect 7098 11636 7104 11648
rect 7156 11636 7162 11688
rect 7208 11648 8984 11676
rect 7208 11608 7236 11648
rect 5736 11580 7236 11608
rect 1719 11577 1731 11580
rect 1673 11571 1731 11577
rect 5902 11500 5908 11552
rect 5960 11540 5966 11552
rect 6457 11543 6515 11549
rect 6457 11540 6469 11543
rect 5960 11512 6469 11540
rect 5960 11500 5966 11512
rect 6457 11509 6469 11512
rect 6503 11509 6515 11543
rect 6457 11503 6515 11509
rect 6641 11543 6699 11549
rect 6641 11509 6653 11543
rect 6687 11540 6699 11543
rect 6730 11540 6736 11552
rect 6687 11512 6736 11540
rect 6687 11509 6699 11512
rect 6641 11503 6699 11509
rect 6730 11500 6736 11512
rect 6788 11500 6794 11552
rect 7742 11500 7748 11552
rect 7800 11540 7806 11552
rect 8110 11540 8116 11552
rect 7800 11512 8116 11540
rect 7800 11500 7806 11512
rect 8110 11500 8116 11512
rect 8168 11540 8174 11552
rect 8849 11543 8907 11549
rect 8849 11540 8861 11543
rect 8168 11512 8861 11540
rect 8168 11500 8174 11512
rect 8849 11509 8861 11512
rect 8895 11509 8907 11543
rect 8956 11540 8984 11648
rect 9692 11620 9720 11707
rect 10318 11704 10324 11756
rect 10376 11704 10382 11756
rect 11422 11744 11428 11756
rect 10704 11716 11428 11744
rect 9861 11679 9919 11685
rect 9861 11645 9873 11679
rect 9907 11676 9919 11679
rect 10704 11676 10732 11716
rect 11422 11704 11428 11716
rect 11480 11744 11486 11756
rect 11609 11747 11667 11753
rect 11609 11744 11621 11747
rect 11480 11716 11621 11744
rect 11480 11704 11486 11716
rect 11609 11713 11621 11716
rect 11655 11713 11667 11747
rect 11716 11744 11744 11840
rect 12406 11812 12434 11852
rect 13814 11840 13820 11892
rect 13872 11880 13878 11892
rect 15197 11883 15255 11889
rect 15197 11880 15209 11883
rect 13872 11852 15209 11880
rect 13872 11840 13878 11852
rect 12406 11784 13676 11812
rect 11977 11747 12035 11753
rect 11977 11744 11989 11747
rect 11716 11716 11989 11744
rect 11609 11707 11667 11713
rect 11977 11713 11989 11716
rect 12023 11713 12035 11747
rect 11977 11707 12035 11713
rect 12066 11704 12072 11756
rect 12124 11704 12130 11756
rect 13170 11704 13176 11756
rect 13228 11704 13234 11756
rect 13648 11753 13676 11784
rect 14384 11753 14412 11852
rect 15197 11849 15209 11852
rect 15243 11880 15255 11883
rect 15470 11880 15476 11892
rect 15243 11852 15476 11880
rect 15243 11849 15255 11852
rect 15197 11843 15255 11849
rect 15470 11840 15476 11852
rect 15528 11880 15534 11892
rect 16666 11880 16672 11892
rect 15528 11852 16672 11880
rect 15528 11840 15534 11852
rect 16666 11840 16672 11852
rect 16724 11840 16730 11892
rect 19705 11883 19763 11889
rect 19705 11849 19717 11883
rect 19751 11880 19763 11883
rect 19978 11880 19984 11892
rect 19751 11852 19984 11880
rect 19751 11849 19763 11852
rect 19705 11843 19763 11849
rect 19978 11840 19984 11852
rect 20036 11840 20042 11892
rect 20070 11840 20076 11892
rect 20128 11880 20134 11892
rect 20901 11883 20959 11889
rect 20901 11880 20913 11883
rect 20128 11852 20300 11880
rect 20128 11840 20134 11852
rect 14642 11772 14648 11824
rect 14700 11812 14706 11824
rect 14829 11815 14887 11821
rect 14829 11812 14841 11815
rect 14700 11784 14841 11812
rect 14700 11772 14706 11784
rect 14829 11781 14841 11784
rect 14875 11812 14887 11815
rect 14875 11784 15424 11812
rect 14875 11781 14887 11784
rect 14829 11775 14887 11781
rect 13357 11747 13415 11753
rect 13357 11713 13369 11747
rect 13403 11713 13415 11747
rect 13357 11707 13415 11713
rect 13633 11747 13691 11753
rect 13633 11713 13645 11747
rect 13679 11713 13691 11747
rect 13633 11707 13691 11713
rect 14369 11747 14427 11753
rect 14369 11713 14381 11747
rect 14415 11713 14427 11747
rect 14737 11747 14795 11753
rect 14737 11744 14749 11747
rect 14369 11707 14427 11713
rect 14568 11716 14749 11744
rect 9907 11648 10732 11676
rect 9907 11645 9919 11648
rect 9861 11639 9919 11645
rect 10778 11636 10784 11688
rect 10836 11636 10842 11688
rect 10873 11679 10931 11685
rect 10873 11645 10885 11679
rect 10919 11676 10931 11679
rect 11790 11676 11796 11688
rect 10919 11648 11796 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 11790 11636 11796 11648
rect 11848 11636 11854 11688
rect 11882 11636 11888 11688
rect 11940 11676 11946 11688
rect 13372 11676 13400 11707
rect 13446 11676 13452 11688
rect 11940 11648 13452 11676
rect 11940 11636 11946 11648
rect 13446 11636 13452 11648
rect 13504 11636 13510 11688
rect 13541 11679 13599 11685
rect 13541 11645 13553 11679
rect 13587 11676 13599 11679
rect 14458 11676 14464 11688
rect 13587 11648 14464 11676
rect 13587 11645 13599 11648
rect 13541 11639 13599 11645
rect 14458 11636 14464 11648
rect 14516 11676 14522 11688
rect 14568 11676 14596 11716
rect 14737 11713 14749 11716
rect 14783 11713 14795 11747
rect 14737 11707 14795 11713
rect 15102 11704 15108 11756
rect 15160 11704 15166 11756
rect 15396 11753 15424 11784
rect 18506 11772 18512 11824
rect 18564 11772 18570 11824
rect 20272 11821 20300 11852
rect 20640 11852 20913 11880
rect 20257 11815 20315 11821
rect 20257 11781 20269 11815
rect 20303 11781 20315 11815
rect 20257 11775 20315 11781
rect 20374 11815 20432 11821
rect 20374 11781 20386 11815
rect 20420 11812 20432 11815
rect 20640 11812 20668 11852
rect 20901 11849 20913 11852
rect 20947 11849 20959 11883
rect 20901 11843 20959 11849
rect 20990 11840 20996 11892
rect 21048 11880 21054 11892
rect 22465 11883 22523 11889
rect 22465 11880 22477 11883
rect 21048 11852 22477 11880
rect 21048 11840 21054 11852
rect 22465 11849 22477 11852
rect 22511 11849 22523 11883
rect 22465 11843 22523 11849
rect 20420 11784 20668 11812
rect 20420 11781 20432 11784
rect 20374 11775 20432 11781
rect 20806 11772 20812 11824
rect 20864 11812 20870 11824
rect 21726 11812 21732 11824
rect 20864 11784 21732 11812
rect 20864 11772 20870 11784
rect 21726 11772 21732 11784
rect 21784 11812 21790 11824
rect 21784 11784 21956 11812
rect 21784 11772 21790 11784
rect 15381 11747 15439 11753
rect 15381 11713 15393 11747
rect 15427 11713 15439 11747
rect 15381 11707 15439 11713
rect 15838 11704 15844 11756
rect 15896 11704 15902 11756
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 14516 11648 14596 11676
rect 14516 11636 14522 11648
rect 14642 11636 14648 11688
rect 14700 11636 14706 11688
rect 15562 11636 15568 11688
rect 15620 11676 15626 11688
rect 15930 11676 15936 11688
rect 15620 11648 15936 11676
rect 15620 11636 15626 11648
rect 15930 11636 15936 11648
rect 15988 11676 15994 11688
rect 16040 11676 16068 11707
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 20174 11753 20232 11759
rect 20174 11750 20186 11753
rect 19392 11716 19932 11744
rect 19392 11704 19398 11716
rect 15988 11648 16068 11676
rect 15988 11636 15994 11648
rect 16942 11636 16948 11688
rect 17000 11676 17006 11688
rect 17221 11679 17279 11685
rect 17221 11676 17233 11679
rect 17000 11648 17233 11676
rect 17000 11636 17006 11648
rect 17221 11645 17233 11648
rect 17267 11645 17279 11679
rect 17497 11679 17555 11685
rect 17497 11676 17509 11679
rect 17221 11639 17279 11645
rect 17328 11648 17509 11676
rect 9674 11568 9680 11620
rect 9732 11608 9738 11620
rect 11146 11608 11152 11620
rect 9732 11580 11152 11608
rect 9732 11568 9738 11580
rect 11146 11568 11152 11580
rect 11204 11568 11210 11620
rect 11422 11568 11428 11620
rect 11480 11608 11486 11620
rect 11480 11580 12434 11608
rect 11480 11568 11486 11580
rect 11974 11540 11980 11552
rect 8956 11512 11980 11540
rect 8849 11503 8907 11509
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12406 11540 12434 11580
rect 12802 11568 12808 11620
rect 12860 11608 12866 11620
rect 17328 11608 17356 11648
rect 17497 11645 17509 11648
rect 17543 11645 17555 11679
rect 17497 11639 17555 11645
rect 18969 11679 19027 11685
rect 18969 11645 18981 11679
rect 19015 11676 19027 11679
rect 19794 11676 19800 11688
rect 19015 11648 19800 11676
rect 19015 11645 19027 11648
rect 18969 11639 19027 11645
rect 19794 11636 19800 11648
rect 19852 11636 19858 11688
rect 19904 11676 19932 11716
rect 20094 11722 20186 11750
rect 20094 11688 20122 11722
rect 20174 11719 20186 11722
rect 20220 11719 20232 11753
rect 20487 11747 20545 11753
rect 20487 11744 20499 11747
rect 20482 11734 20499 11744
rect 20174 11713 20232 11719
rect 20364 11713 20499 11734
rect 20533 11713 20545 11747
rect 20364 11707 20545 11713
rect 20625 11750 20683 11753
rect 20714 11750 20720 11756
rect 20625 11747 20720 11750
rect 20625 11713 20637 11747
rect 20671 11722 20720 11747
rect 20671 11713 20683 11722
rect 20625 11707 20683 11713
rect 20364 11706 20510 11707
rect 19981 11679 20039 11685
rect 19981 11676 19993 11679
rect 19904 11648 19993 11676
rect 19981 11645 19993 11648
rect 20027 11645 20039 11679
rect 19981 11639 20039 11645
rect 20076 11636 20082 11688
rect 20134 11636 20140 11688
rect 12860 11580 17356 11608
rect 12860 11568 12866 11580
rect 19426 11568 19432 11620
rect 19484 11608 19490 11620
rect 20364 11608 20392 11706
rect 20714 11704 20720 11722
rect 20772 11704 20778 11756
rect 21450 11704 21456 11756
rect 21508 11704 21514 11756
rect 21928 11753 21956 11784
rect 22094 11772 22100 11824
rect 22152 11772 22158 11824
rect 23842 11772 23848 11824
rect 23900 11812 23906 11824
rect 24121 11815 24179 11821
rect 24121 11812 24133 11815
rect 23900 11784 24133 11812
rect 23900 11772 23906 11784
rect 24121 11781 24133 11784
rect 24167 11781 24179 11815
rect 24121 11775 24179 11781
rect 21913 11747 21971 11753
rect 21913 11713 21925 11747
rect 21959 11713 21971 11747
rect 21913 11707 21971 11713
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22281 11747 22339 11753
rect 22281 11713 22293 11747
rect 22327 11744 22339 11747
rect 22738 11744 22744 11756
rect 22327 11716 22744 11744
rect 22327 11713 22339 11716
rect 22281 11707 22339 11713
rect 22738 11704 22744 11716
rect 22796 11704 22802 11756
rect 22925 11747 22983 11753
rect 22925 11713 22937 11747
rect 22971 11744 22983 11747
rect 23014 11744 23020 11756
rect 22971 11716 23020 11744
rect 22971 11713 22983 11716
rect 22925 11707 22983 11713
rect 23014 11704 23020 11716
rect 23072 11704 23078 11756
rect 23382 11704 23388 11756
rect 23440 11744 23446 11756
rect 23569 11747 23627 11753
rect 23569 11744 23581 11747
rect 23440 11716 23581 11744
rect 23440 11704 23446 11716
rect 23569 11713 23581 11716
rect 23615 11713 23627 11747
rect 23569 11707 23627 11713
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11713 24363 11747
rect 24305 11707 24363 11713
rect 21082 11636 21088 11688
rect 21140 11676 21146 11688
rect 21177 11679 21235 11685
rect 21177 11676 21189 11679
rect 21140 11648 21189 11676
rect 21140 11636 21146 11648
rect 21177 11645 21189 11648
rect 21223 11645 21235 11679
rect 21177 11639 21235 11645
rect 21358 11636 21364 11688
rect 21416 11676 21422 11688
rect 24320 11676 24348 11707
rect 21416 11648 24348 11676
rect 21416 11636 21422 11648
rect 22186 11608 22192 11620
rect 19484 11580 22192 11608
rect 19484 11568 19490 11580
rect 22186 11568 22192 11580
rect 22244 11568 22250 11620
rect 14461 11543 14519 11549
rect 14461 11540 14473 11543
rect 12406 11512 14473 11540
rect 14461 11509 14473 11512
rect 14507 11540 14519 11543
rect 15102 11540 15108 11552
rect 14507 11512 15108 11540
rect 14507 11509 14519 11512
rect 14461 11503 14519 11509
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 15565 11543 15623 11549
rect 15565 11509 15577 11543
rect 15611 11540 15623 11543
rect 15930 11540 15936 11552
rect 15611 11512 15936 11540
rect 15611 11509 15623 11512
rect 15565 11503 15623 11509
rect 15930 11500 15936 11512
rect 15988 11500 15994 11552
rect 16022 11500 16028 11552
rect 16080 11500 16086 11552
rect 19613 11543 19671 11549
rect 19613 11509 19625 11543
rect 19659 11540 19671 11543
rect 21266 11540 21272 11552
rect 19659 11512 21272 11540
rect 19659 11509 19671 11512
rect 19613 11503 19671 11509
rect 21266 11500 21272 11512
rect 21324 11500 21330 11552
rect 21361 11543 21419 11549
rect 21361 11509 21373 11543
rect 21407 11540 21419 11543
rect 21542 11540 21548 11552
rect 21407 11512 21548 11540
rect 21407 11509 21419 11512
rect 21361 11503 21419 11509
rect 21542 11500 21548 11512
rect 21600 11500 21606 11552
rect 1104 11450 24840 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 20214 11450
rect 20266 11398 20278 11450
rect 20330 11398 20342 11450
rect 20394 11398 20406 11450
rect 20458 11398 20470 11450
rect 20522 11398 24840 11450
rect 1104 11376 24840 11398
rect 2041 11339 2099 11345
rect 2041 11305 2053 11339
rect 2087 11336 2099 11339
rect 2130 11336 2136 11348
rect 2087 11308 2136 11336
rect 2087 11305 2099 11308
rect 2041 11299 2099 11305
rect 2130 11296 2136 11308
rect 2188 11296 2194 11348
rect 4525 11339 4583 11345
rect 4525 11305 4537 11339
rect 4571 11336 4583 11339
rect 4706 11336 4712 11348
rect 4571 11308 4712 11336
rect 4571 11305 4583 11308
rect 4525 11299 4583 11305
rect 4706 11296 4712 11308
rect 4764 11296 4770 11348
rect 4890 11296 4896 11348
rect 4948 11296 4954 11348
rect 5368 11308 7328 11336
rect 2225 11271 2283 11277
rect 2225 11237 2237 11271
rect 2271 11268 2283 11271
rect 2958 11268 2964 11280
rect 2271 11240 2964 11268
rect 2271 11237 2283 11240
rect 2225 11231 2283 11237
rect 2958 11228 2964 11240
rect 3016 11228 3022 11280
rect 5368 11268 5396 11308
rect 4356 11240 5396 11268
rect 7300 11268 7328 11308
rect 7374 11296 7380 11348
rect 7432 11296 7438 11348
rect 9309 11339 9367 11345
rect 9309 11305 9321 11339
rect 9355 11336 9367 11339
rect 10778 11336 10784 11348
rect 9355 11308 10784 11336
rect 9355 11305 9367 11308
rect 9309 11299 9367 11305
rect 10778 11296 10784 11308
rect 10836 11296 10842 11348
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 13633 11339 13691 11345
rect 13633 11336 13645 11339
rect 13320 11308 13645 11336
rect 13320 11296 13326 11308
rect 13633 11305 13645 11308
rect 13679 11305 13691 11339
rect 13633 11299 13691 11305
rect 19889 11339 19947 11345
rect 19889 11305 19901 11339
rect 19935 11336 19947 11339
rect 22741 11339 22799 11345
rect 19935 11308 21220 11336
rect 19935 11305 19947 11308
rect 19889 11299 19947 11305
rect 21192 11280 21220 11308
rect 22741 11305 22753 11339
rect 22787 11336 22799 11339
rect 23106 11336 23112 11348
rect 22787 11308 23112 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 23106 11296 23112 11308
rect 23164 11296 23170 11348
rect 7834 11268 7840 11280
rect 7300 11240 7840 11268
rect 3142 11160 3148 11212
rect 3200 11200 3206 11212
rect 3418 11200 3424 11212
rect 3200 11172 3424 11200
rect 3200 11160 3206 11172
rect 3418 11160 3424 11172
rect 3476 11160 3482 11212
rect 2961 11135 3019 11141
rect 2961 11101 2973 11135
rect 3007 11132 3019 11135
rect 3234 11132 3240 11144
rect 3007 11104 3240 11132
rect 3007 11101 3019 11104
rect 2961 11095 3019 11101
rect 3234 11092 3240 11104
rect 3292 11092 3298 11144
rect 4356 11141 4384 11240
rect 7834 11228 7840 11240
rect 7892 11268 7898 11280
rect 8389 11271 8447 11277
rect 8389 11268 8401 11271
rect 7892 11240 8401 11268
rect 7892 11228 7898 11240
rect 8389 11237 8401 11240
rect 8435 11268 8447 11271
rect 8754 11268 8760 11280
rect 8435 11240 8760 11268
rect 8435 11237 8447 11240
rect 8389 11231 8447 11237
rect 8754 11228 8760 11240
rect 8812 11228 8818 11280
rect 11241 11271 11299 11277
rect 9048 11240 10180 11268
rect 6365 11203 6423 11209
rect 6365 11169 6377 11203
rect 6411 11200 6423 11203
rect 6914 11200 6920 11212
rect 6411 11172 6920 11200
rect 6411 11169 6423 11172
rect 6365 11163 6423 11169
rect 6914 11160 6920 11172
rect 6972 11160 6978 11212
rect 7466 11160 7472 11212
rect 7524 11200 7530 11212
rect 7926 11200 7932 11212
rect 7524 11172 7932 11200
rect 7524 11160 7530 11172
rect 7926 11160 7932 11172
rect 7984 11160 7990 11212
rect 4341 11135 4399 11141
rect 4341 11101 4353 11135
rect 4387 11101 4399 11135
rect 4341 11095 4399 11101
rect 6638 11092 6644 11144
rect 6696 11092 6702 11144
rect 7742 11092 7748 11144
rect 7800 11092 7806 11144
rect 9048 11141 9076 11240
rect 9950 11200 9956 11212
rect 9324 11172 9956 11200
rect 9324 11141 9352 11172
rect 9950 11160 9956 11172
rect 10008 11160 10014 11212
rect 10152 11200 10180 11240
rect 11241 11237 11253 11271
rect 11287 11237 11299 11271
rect 11241 11231 11299 11237
rect 10410 11200 10416 11212
rect 10152 11172 10416 11200
rect 10410 11160 10416 11172
rect 10468 11200 10474 11212
rect 11057 11203 11115 11209
rect 11057 11200 11069 11203
rect 10468 11172 11069 11200
rect 10468 11160 10474 11172
rect 11057 11169 11069 11172
rect 11103 11169 11115 11203
rect 11256 11200 11284 11231
rect 11698 11228 11704 11280
rect 11756 11268 11762 11280
rect 19702 11268 19708 11280
rect 11756 11240 13400 11268
rect 11756 11228 11762 11240
rect 11606 11200 11612 11212
rect 11256 11172 11612 11200
rect 11057 11163 11115 11169
rect 11606 11160 11612 11172
rect 11664 11200 11670 11212
rect 13170 11200 13176 11212
rect 11664 11172 13176 11200
rect 11664 11160 11670 11172
rect 13170 11160 13176 11172
rect 13228 11200 13234 11212
rect 13228 11172 13308 11200
rect 13228 11160 13234 11172
rect 9033 11135 9091 11141
rect 9033 11101 9045 11135
rect 9079 11101 9091 11135
rect 9033 11095 9091 11101
rect 9309 11135 9367 11141
rect 9309 11101 9321 11135
rect 9355 11101 9367 11135
rect 9309 11095 9367 11101
rect 9674 11092 9680 11144
rect 9732 11132 9738 11144
rect 9769 11135 9827 11141
rect 9769 11132 9781 11135
rect 9732 11104 9781 11132
rect 9732 11092 9738 11104
rect 9769 11101 9781 11104
rect 9815 11101 9827 11135
rect 9769 11095 9827 11101
rect 9858 11092 9864 11144
rect 9916 11092 9922 11144
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10229 11135 10287 11141
rect 10229 11132 10241 11135
rect 10192 11104 10241 11132
rect 10192 11092 10198 11104
rect 10229 11101 10241 11104
rect 10275 11101 10287 11135
rect 10229 11095 10287 11101
rect 10778 11092 10784 11144
rect 10836 11092 10842 11144
rect 11422 11092 11428 11144
rect 11480 11092 11486 11144
rect 11793 11135 11851 11141
rect 11793 11101 11805 11135
rect 11839 11101 11851 11135
rect 11793 11095 11851 11101
rect 1854 11024 1860 11076
rect 1912 11024 1918 11076
rect 2038 11024 2044 11076
rect 2096 11073 2102 11076
rect 2096 11067 2115 11073
rect 2103 11033 2115 11067
rect 2096 11027 2115 11033
rect 2096 11024 2102 11027
rect 5902 11024 5908 11076
rect 5960 11024 5966 11076
rect 8573 11067 8631 11073
rect 8573 11033 8585 11067
rect 8619 11064 8631 11067
rect 8662 11064 8668 11076
rect 8619 11036 8668 11064
rect 8619 11033 8631 11036
rect 8573 11027 8631 11033
rect 8662 11024 8668 11036
rect 8720 11024 8726 11076
rect 9125 11067 9183 11073
rect 9125 11033 9137 11067
rect 9171 11064 9183 11067
rect 9171 11036 9352 11064
rect 9171 11033 9183 11036
rect 9125 11027 9183 11033
rect 1946 10956 1952 11008
rect 2004 10996 2010 11008
rect 2501 10999 2559 11005
rect 2501 10996 2513 10999
rect 2004 10968 2513 10996
rect 2004 10956 2010 10968
rect 2501 10965 2513 10968
rect 2547 10965 2559 10999
rect 2501 10959 2559 10965
rect 2866 10956 2872 11008
rect 2924 10956 2930 11008
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 7837 10999 7895 11005
rect 7837 10996 7849 10999
rect 7064 10968 7849 10996
rect 7064 10956 7070 10968
rect 7837 10965 7849 10968
rect 7883 10996 7895 10999
rect 8110 10996 8116 11008
rect 7883 10968 8116 10996
rect 7883 10965 7895 10968
rect 7837 10959 7895 10965
rect 8110 10956 8116 10968
rect 8168 10956 8174 11008
rect 9324 10996 9352 11036
rect 9398 11024 9404 11076
rect 9456 11064 9462 11076
rect 9585 11067 9643 11073
rect 9585 11064 9597 11067
rect 9456 11036 9597 11064
rect 9456 11024 9462 11036
rect 9585 11033 9597 11036
rect 9631 11033 9643 11067
rect 10594 11064 10600 11076
rect 9585 11027 9643 11033
rect 9692 11036 10600 11064
rect 9692 10996 9720 11036
rect 10594 11024 10600 11036
rect 10652 11024 10658 11076
rect 11146 11024 11152 11076
rect 11204 11064 11210 11076
rect 11808 11064 11836 11095
rect 11882 11092 11888 11144
rect 11940 11132 11946 11144
rect 13280 11141 13308 11172
rect 13372 11141 13400 11240
rect 19628 11240 19708 11268
rect 13446 11160 13452 11212
rect 13504 11160 13510 11212
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 15105 11203 15163 11209
rect 15105 11200 15117 11203
rect 15068 11172 15117 11200
rect 15068 11160 15074 11172
rect 15105 11169 15117 11172
rect 15151 11200 15163 11203
rect 16669 11203 16727 11209
rect 15151 11172 16068 11200
rect 15151 11169 15163 11172
rect 15105 11163 15163 11169
rect 12345 11135 12403 11141
rect 12345 11132 12357 11135
rect 11940 11104 12357 11132
rect 11940 11092 11946 11104
rect 12345 11101 12357 11104
rect 12391 11101 12403 11135
rect 12345 11095 12403 11101
rect 13265 11135 13323 11141
rect 13265 11101 13277 11135
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 13357 11135 13415 11141
rect 13357 11101 13369 11135
rect 13403 11101 13415 11135
rect 13357 11095 13415 11101
rect 13630 11092 13636 11144
rect 13688 11092 13694 11144
rect 13814 11092 13820 11144
rect 13872 11132 13878 11144
rect 15654 11132 15660 11144
rect 13872 11104 15660 11132
rect 13872 11092 13878 11104
rect 15654 11092 15660 11104
rect 15712 11132 15718 11144
rect 16040 11141 16068 11172
rect 16669 11169 16681 11203
rect 16715 11200 16727 11203
rect 16942 11200 16948 11212
rect 16715 11172 16948 11200
rect 16715 11169 16727 11172
rect 16669 11163 16727 11169
rect 16942 11160 16948 11172
rect 17000 11160 17006 11212
rect 19628 11209 19656 11240
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 20622 11228 20628 11280
rect 20680 11228 20686 11280
rect 21174 11228 21180 11280
rect 21232 11268 21238 11280
rect 22002 11268 22008 11280
rect 21232 11240 22008 11268
rect 21232 11228 21238 11240
rect 22002 11228 22008 11240
rect 22060 11228 22066 11280
rect 22094 11228 22100 11280
rect 22152 11228 22158 11280
rect 22281 11271 22339 11277
rect 22281 11237 22293 11271
rect 22327 11237 22339 11271
rect 22281 11231 22339 11237
rect 19613 11203 19671 11209
rect 19613 11169 19625 11203
rect 19659 11200 19671 11203
rect 20640 11200 20668 11228
rect 21085 11203 21143 11209
rect 19659 11172 20576 11200
rect 20640 11172 20760 11200
rect 19659 11169 19671 11172
rect 19613 11163 19671 11169
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 15712 11104 15853 11132
rect 15712 11092 15718 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 16025 11135 16083 11141
rect 16025 11101 16037 11135
rect 16071 11101 16083 11135
rect 16025 11095 16083 11101
rect 16117 11135 16175 11141
rect 16117 11101 16129 11135
rect 16163 11101 16175 11135
rect 16117 11095 16175 11101
rect 11204 11036 11928 11064
rect 11204 11024 11210 11036
rect 11900 11008 11928 11036
rect 12618 11024 12624 11076
rect 12676 11064 12682 11076
rect 12897 11067 12955 11073
rect 12897 11064 12909 11067
rect 12676 11036 12909 11064
rect 12676 11024 12682 11036
rect 12897 11033 12909 11036
rect 12943 11064 12955 11067
rect 13648 11064 13676 11092
rect 12943 11036 13676 11064
rect 15289 11067 15347 11073
rect 12943 11033 12955 11036
rect 12897 11027 12955 11033
rect 15289 11033 15301 11067
rect 15335 11064 15347 11067
rect 15378 11064 15384 11076
rect 15335 11036 15384 11064
rect 15335 11033 15347 11036
rect 15289 11027 15347 11033
rect 15378 11024 15384 11036
rect 15436 11024 15442 11076
rect 9324 10968 9720 10996
rect 10042 10956 10048 11008
rect 10100 10956 10106 11008
rect 10137 10999 10195 11005
rect 10137 10965 10149 10999
rect 10183 10996 10195 10999
rect 10318 10996 10324 11008
rect 10183 10968 10324 10996
rect 10183 10965 10195 10968
rect 10137 10959 10195 10965
rect 10318 10956 10324 10968
rect 10376 10956 10382 11008
rect 11882 10956 11888 11008
rect 11940 10956 11946 11008
rect 15654 10956 15660 11008
rect 15712 10956 15718 11008
rect 15838 10956 15844 11008
rect 15896 10996 15902 11008
rect 16132 10996 16160 11095
rect 18046 11092 18052 11144
rect 18104 11092 18110 11144
rect 19705 11135 19763 11141
rect 19705 11101 19717 11135
rect 19751 11132 19763 11135
rect 19886 11132 19892 11144
rect 19751 11104 19892 11132
rect 19751 11101 19763 11104
rect 19705 11095 19763 11101
rect 19886 11092 19892 11104
rect 19944 11132 19950 11144
rect 20441 11135 20499 11141
rect 20441 11132 20453 11135
rect 19944 11104 20453 11132
rect 19944 11092 19950 11104
rect 20441 11101 20453 11104
rect 20487 11101 20499 11135
rect 20548 11132 20576 11172
rect 20622 11132 20628 11144
rect 20548 11104 20628 11132
rect 20441 11095 20499 11101
rect 20622 11092 20628 11104
rect 20680 11092 20686 11144
rect 20732 11141 20760 11172
rect 21085 11169 21097 11203
rect 21131 11169 21143 11203
rect 22112 11200 22140 11228
rect 21085 11163 21143 11169
rect 21928 11172 22140 11200
rect 22296 11200 22324 11231
rect 23014 11200 23020 11212
rect 22296 11172 23020 11200
rect 20717 11135 20775 11141
rect 20717 11101 20729 11135
rect 20763 11101 20775 11135
rect 20717 11095 20775 11101
rect 20809 11135 20867 11141
rect 20809 11101 20821 11135
rect 20855 11132 20867 11135
rect 20990 11132 20996 11144
rect 20855 11104 20996 11132
rect 20855 11101 20867 11104
rect 20809 11095 20867 11101
rect 16574 11024 16580 11076
rect 16632 11064 16638 11076
rect 16945 11067 17003 11073
rect 16945 11064 16957 11067
rect 16632 11036 16957 11064
rect 16632 11024 16638 11036
rect 16945 11033 16957 11036
rect 16991 11033 17003 11067
rect 16945 11027 17003 11033
rect 18693 11067 18751 11073
rect 18693 11033 18705 11067
rect 18739 11064 18751 11067
rect 20824 11064 20852 11095
rect 20990 11092 20996 11104
rect 21048 11092 21054 11144
rect 21100 11132 21128 11163
rect 21637 11135 21695 11141
rect 21637 11132 21649 11135
rect 21100 11104 21649 11132
rect 21637 11101 21649 11104
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 21726 11092 21732 11144
rect 21784 11132 21790 11144
rect 21928 11141 21956 11172
rect 23014 11160 23020 11172
rect 23072 11160 23078 11212
rect 23845 11203 23903 11209
rect 23845 11200 23857 11203
rect 23124 11172 23857 11200
rect 21913 11135 21971 11141
rect 21784 11104 21829 11132
rect 21784 11092 21790 11104
rect 21913 11101 21925 11135
rect 21959 11101 21971 11135
rect 21913 11095 21971 11101
rect 22143 11135 22201 11141
rect 22143 11101 22155 11135
rect 22189 11132 22201 11135
rect 22557 11135 22615 11141
rect 22189 11104 22508 11132
rect 22189 11101 22201 11104
rect 22143 11095 22201 11101
rect 18739 11036 20852 11064
rect 22005 11067 22063 11073
rect 18739 11033 18751 11036
rect 18693 11027 18751 11033
rect 22005 11033 22017 11067
rect 22051 11033 22063 11067
rect 22480 11064 22508 11104
rect 22557 11101 22569 11135
rect 22603 11132 22615 11135
rect 22830 11132 22836 11144
rect 22603 11104 22836 11132
rect 22603 11101 22615 11104
rect 22557 11095 22615 11101
rect 22830 11092 22836 11104
rect 22888 11132 22894 11144
rect 23124 11132 23152 11172
rect 23845 11169 23857 11172
rect 23891 11169 23903 11203
rect 23845 11163 23903 11169
rect 22888 11104 23152 11132
rect 22888 11092 22894 11104
rect 23658 11092 23664 11144
rect 23716 11132 23722 11144
rect 24029 11135 24087 11141
rect 24029 11132 24041 11135
rect 23716 11104 24041 11132
rect 23716 11092 23722 11104
rect 24029 11101 24041 11104
rect 24075 11101 24087 11135
rect 24029 11095 24087 11101
rect 22480 11036 23336 11064
rect 22005 11027 22063 11033
rect 18708 10996 18736 11027
rect 15896 10968 18736 10996
rect 22020 10996 22048 11027
rect 22186 10996 22192 11008
rect 22020 10968 22192 10996
rect 15896 10956 15902 10968
rect 22186 10956 22192 10968
rect 22244 10996 22250 11008
rect 23106 10996 23112 11008
rect 22244 10968 23112 10996
rect 22244 10956 22250 10968
rect 23106 10956 23112 10968
rect 23164 10956 23170 11008
rect 23308 10996 23336 11036
rect 23382 11024 23388 11076
rect 23440 11064 23446 11076
rect 23477 11067 23535 11073
rect 23477 11064 23489 11067
rect 23440 11036 23489 11064
rect 23440 11024 23446 11036
rect 23477 11033 23489 11036
rect 23523 11033 23535 11067
rect 23477 11027 23535 11033
rect 23566 11024 23572 11076
rect 23624 11024 23630 11076
rect 23658 10996 23664 11008
rect 23308 10968 23664 10996
rect 23658 10956 23664 10968
rect 23716 10956 23722 11008
rect 1104 10906 24840 10928
rect 1104 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 24214 10906
rect 24266 10854 24278 10906
rect 24330 10854 24342 10906
rect 24394 10854 24406 10906
rect 24458 10854 24470 10906
rect 24522 10854 24840 10906
rect 1104 10832 24840 10854
rect 2866 10752 2872 10804
rect 2924 10792 2930 10804
rect 3234 10792 3240 10804
rect 2924 10764 3240 10792
rect 2924 10752 2930 10764
rect 3234 10752 3240 10764
rect 3292 10792 3298 10804
rect 3421 10795 3479 10801
rect 3421 10792 3433 10795
rect 3292 10764 3433 10792
rect 3292 10752 3298 10764
rect 3421 10761 3433 10764
rect 3467 10761 3479 10795
rect 3421 10755 3479 10761
rect 5626 10752 5632 10804
rect 5684 10792 5690 10804
rect 7761 10795 7819 10801
rect 7761 10792 7773 10795
rect 5684 10764 7773 10792
rect 5684 10752 5690 10764
rect 7761 10761 7773 10764
rect 7807 10792 7819 10795
rect 9122 10792 9128 10804
rect 7807 10764 9128 10792
rect 7807 10761 7819 10764
rect 7761 10755 7819 10761
rect 9122 10752 9128 10764
rect 9180 10792 9186 10804
rect 9306 10792 9312 10804
rect 9180 10764 9312 10792
rect 9180 10752 9186 10764
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 10042 10752 10048 10804
rect 10100 10792 10106 10804
rect 10870 10792 10876 10804
rect 10100 10764 10876 10792
rect 10100 10752 10106 10764
rect 10870 10752 10876 10764
rect 10928 10752 10934 10804
rect 15562 10752 15568 10804
rect 15620 10792 15626 10804
rect 15620 10764 15700 10792
rect 15620 10752 15626 10764
rect 1946 10684 1952 10736
rect 2004 10684 2010 10736
rect 2958 10684 2964 10736
rect 3016 10684 3022 10736
rect 5074 10684 5080 10736
rect 5132 10684 5138 10736
rect 6546 10684 6552 10736
rect 6604 10724 6610 10736
rect 7561 10727 7619 10733
rect 7561 10724 7573 10727
rect 6604 10696 7573 10724
rect 6604 10684 6610 10696
rect 7561 10693 7573 10696
rect 7607 10693 7619 10727
rect 7561 10687 7619 10693
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 6687 10628 7420 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 1486 10548 1492 10600
rect 1544 10588 1550 10600
rect 1673 10591 1731 10597
rect 1673 10588 1685 10591
rect 1544 10560 1685 10588
rect 1544 10548 1550 10560
rect 1673 10557 1685 10560
rect 1719 10557 1731 10591
rect 1673 10551 1731 10557
rect 4065 10591 4123 10597
rect 4065 10557 4077 10591
rect 4111 10588 4123 10591
rect 4111 10560 4844 10588
rect 4111 10557 4123 10560
rect 4065 10551 4123 10557
rect 4816 10452 4844 10560
rect 5350 10548 5356 10600
rect 5408 10588 5414 10600
rect 5813 10591 5871 10597
rect 5813 10588 5825 10591
rect 5408 10560 5825 10588
rect 5408 10548 5414 10560
rect 5813 10557 5825 10560
rect 5859 10557 5871 10591
rect 5813 10551 5871 10557
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10557 6147 10591
rect 6089 10551 6147 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10588 6975 10591
rect 7006 10588 7012 10600
rect 6963 10560 7012 10588
rect 6963 10557 6975 10560
rect 6917 10551 6975 10557
rect 6104 10520 6132 10551
rect 7006 10548 7012 10560
rect 7064 10548 7070 10600
rect 6638 10520 6644 10532
rect 6104 10492 6644 10520
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 7392 10520 7420 10628
rect 7576 10588 7604 10687
rect 7926 10684 7932 10736
rect 7984 10724 7990 10736
rect 8205 10727 8263 10733
rect 8205 10724 8217 10727
rect 7984 10696 8217 10724
rect 7984 10684 7990 10696
rect 8205 10693 8217 10696
rect 8251 10693 8263 10727
rect 8205 10687 8263 10693
rect 9858 10684 9864 10736
rect 9916 10724 9922 10736
rect 10962 10724 10968 10736
rect 9916 10696 10968 10724
rect 9916 10684 9922 10696
rect 10962 10684 10968 10696
rect 11020 10684 11026 10736
rect 11790 10684 11796 10736
rect 11848 10724 11854 10736
rect 11885 10727 11943 10733
rect 11885 10724 11897 10727
rect 11848 10696 11897 10724
rect 11848 10684 11854 10696
rect 11885 10693 11897 10696
rect 11931 10693 11943 10727
rect 12894 10724 12900 10736
rect 11885 10687 11943 10693
rect 11992 10696 12900 10724
rect 8110 10616 8116 10668
rect 8168 10656 8174 10668
rect 8389 10659 8447 10665
rect 8389 10656 8401 10659
rect 8168 10628 8401 10656
rect 8168 10616 8174 10628
rect 8389 10625 8401 10628
rect 8435 10625 8447 10659
rect 8389 10619 8447 10625
rect 8481 10659 8539 10665
rect 8481 10625 8493 10659
rect 8527 10656 8539 10659
rect 8570 10656 8576 10668
rect 8527 10628 8576 10656
rect 8527 10625 8539 10628
rect 8481 10619 8539 10625
rect 8570 10616 8576 10628
rect 8628 10616 8634 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 9769 10659 9827 10665
rect 9769 10656 9781 10659
rect 9732 10628 9781 10656
rect 9732 10616 9738 10628
rect 9769 10625 9781 10628
rect 9815 10625 9827 10659
rect 11241 10659 11299 10665
rect 11241 10656 11253 10659
rect 9769 10619 9827 10625
rect 9876 10628 11253 10656
rect 8938 10588 8944 10600
rect 7576 10560 8432 10588
rect 8205 10523 8263 10529
rect 8205 10520 8217 10523
rect 7392 10492 8217 10520
rect 8205 10489 8217 10492
rect 8251 10489 8263 10523
rect 8404 10520 8432 10560
rect 8588 10560 8944 10588
rect 8588 10520 8616 10560
rect 8938 10548 8944 10560
rect 8996 10588 9002 10600
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8996 10560 9137 10588
rect 8996 10548 9002 10560
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9876 10588 9904 10628
rect 11241 10625 11253 10628
rect 11287 10656 11299 10659
rect 11992 10656 12020 10696
rect 12894 10684 12900 10696
rect 12952 10684 12958 10736
rect 15102 10684 15108 10736
rect 15160 10724 15166 10736
rect 15197 10727 15255 10733
rect 15197 10724 15209 10727
rect 15160 10696 15209 10724
rect 15160 10684 15166 10696
rect 15197 10693 15209 10696
rect 15243 10693 15255 10727
rect 15197 10687 15255 10693
rect 11287 10628 12020 10656
rect 12437 10659 12495 10665
rect 11287 10625 11299 10628
rect 11241 10619 11299 10625
rect 12437 10625 12449 10659
rect 12483 10656 12495 10659
rect 12618 10656 12624 10668
rect 12483 10628 12624 10656
rect 12483 10625 12495 10628
rect 12437 10619 12495 10625
rect 12618 10616 12624 10628
rect 12676 10616 12682 10668
rect 12989 10659 13047 10665
rect 12989 10625 13001 10659
rect 13035 10656 13047 10659
rect 13262 10656 13268 10668
rect 13035 10628 13268 10656
rect 13035 10625 13047 10628
rect 12989 10619 13047 10625
rect 13262 10616 13268 10628
rect 13320 10616 13326 10668
rect 13722 10616 13728 10668
rect 13780 10616 13786 10668
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 15286 10656 15292 10668
rect 14507 10628 15292 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 15286 10616 15292 10628
rect 15344 10656 15350 10668
rect 15565 10659 15623 10665
rect 15565 10656 15577 10659
rect 15344 10628 15577 10656
rect 15344 10616 15350 10628
rect 15565 10625 15577 10628
rect 15611 10625 15623 10659
rect 15565 10619 15623 10625
rect 15672 10656 15700 10764
rect 16022 10752 16028 10804
rect 16080 10752 16086 10804
rect 16301 10795 16359 10801
rect 16301 10761 16313 10795
rect 16347 10792 16359 10795
rect 16574 10792 16580 10804
rect 16347 10764 16580 10792
rect 16347 10761 16359 10764
rect 16301 10755 16359 10761
rect 16574 10752 16580 10764
rect 16632 10752 16638 10804
rect 18782 10752 18788 10804
rect 18840 10792 18846 10804
rect 18840 10764 20576 10792
rect 18840 10752 18846 10764
rect 16040 10724 16068 10752
rect 16040 10696 16436 10724
rect 16408 10665 16436 10696
rect 17954 10684 17960 10736
rect 18012 10684 18018 10736
rect 20548 10733 20576 10764
rect 20622 10752 20628 10804
rect 20680 10792 20686 10804
rect 21450 10792 21456 10804
rect 20680 10764 21456 10792
rect 20680 10752 20686 10764
rect 21450 10752 21456 10764
rect 21508 10752 21514 10804
rect 21545 10795 21603 10801
rect 21545 10761 21557 10795
rect 21591 10792 21603 10795
rect 23382 10792 23388 10804
rect 21591 10764 23388 10792
rect 21591 10761 21603 10764
rect 21545 10755 21603 10761
rect 23382 10752 23388 10764
rect 23440 10752 23446 10804
rect 23566 10752 23572 10804
rect 23624 10792 23630 10804
rect 24029 10795 24087 10801
rect 24029 10792 24041 10795
rect 23624 10764 24041 10792
rect 23624 10752 23630 10764
rect 24029 10761 24041 10764
rect 24075 10761 24087 10795
rect 24029 10755 24087 10761
rect 20533 10727 20591 10733
rect 20533 10693 20545 10727
rect 20579 10693 20591 10727
rect 20533 10687 20591 10693
rect 22281 10727 22339 10733
rect 22281 10693 22293 10727
rect 22327 10724 22339 10727
rect 23290 10724 23296 10736
rect 22327 10696 23296 10724
rect 22327 10693 22339 10696
rect 22281 10687 22339 10693
rect 23290 10684 23296 10696
rect 23348 10724 23354 10736
rect 23477 10727 23535 10733
rect 23477 10724 23489 10727
rect 23348 10696 23489 10724
rect 23348 10684 23354 10696
rect 23477 10693 23489 10696
rect 23523 10693 23535 10727
rect 23477 10687 23535 10693
rect 16025 10659 16083 10665
rect 16025 10656 16037 10659
rect 15672 10628 16037 10656
rect 9125 10551 9183 10557
rect 9232 10560 9904 10588
rect 8404 10492 8616 10520
rect 8205 10483 8263 10489
rect 9030 10480 9036 10532
rect 9088 10520 9094 10532
rect 9232 10520 9260 10560
rect 10318 10548 10324 10600
rect 10376 10588 10382 10600
rect 10756 10591 10814 10597
rect 10756 10588 10768 10591
rect 10376 10560 10768 10588
rect 10376 10548 10382 10560
rect 10756 10557 10768 10560
rect 10802 10557 10814 10591
rect 10756 10551 10814 10557
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 12897 10591 12955 10597
rect 12897 10588 12909 10591
rect 11940 10560 12909 10588
rect 11940 10548 11946 10560
rect 12897 10557 12909 10560
rect 12943 10557 12955 10591
rect 15672 10588 15700 10628
rect 16025 10625 16037 10628
rect 16071 10625 16083 10659
rect 16025 10619 16083 10625
rect 16117 10659 16175 10665
rect 16117 10625 16129 10659
rect 16163 10656 16175 10659
rect 16393 10659 16451 10665
rect 16163 10628 16344 10656
rect 16163 10625 16175 10628
rect 16117 10619 16175 10625
rect 12897 10551 12955 10557
rect 15120 10560 15700 10588
rect 9088 10492 9260 10520
rect 9088 10480 9094 10492
rect 9766 10480 9772 10532
rect 9824 10520 9830 10532
rect 10597 10523 10655 10529
rect 10597 10520 10609 10523
rect 9824 10492 10609 10520
rect 9824 10480 9830 10492
rect 10597 10489 10609 10492
rect 10643 10520 10655 10523
rect 15120 10520 15148 10560
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 16209 10591 16267 10597
rect 16209 10588 16221 10591
rect 15988 10560 16221 10588
rect 15988 10548 15994 10560
rect 16209 10557 16221 10560
rect 16255 10557 16267 10591
rect 16209 10551 16267 10557
rect 10643 10492 15148 10520
rect 10643 10489 10655 10492
rect 10597 10483 10655 10489
rect 15194 10480 15200 10532
rect 15252 10520 15258 10532
rect 16316 10520 16344 10628
rect 16393 10625 16405 10659
rect 16439 10625 16451 10659
rect 16393 10619 16451 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10656 21511 10659
rect 21499 10628 22784 10656
rect 21499 10625 21511 10628
rect 21453 10619 21511 10625
rect 16942 10548 16948 10600
rect 17000 10588 17006 10600
rect 17037 10591 17095 10597
rect 17037 10588 17049 10591
rect 17000 10560 17049 10588
rect 17000 10548 17006 10560
rect 17037 10557 17049 10560
rect 17083 10557 17095 10591
rect 17037 10551 17095 10557
rect 17310 10548 17316 10600
rect 17368 10548 17374 10600
rect 21542 10548 21548 10600
rect 21600 10588 21606 10600
rect 22373 10591 22431 10597
rect 22373 10588 22385 10591
rect 21600 10560 22385 10588
rect 21600 10548 21606 10560
rect 22373 10557 22385 10560
rect 22419 10557 22431 10591
rect 22373 10551 22431 10557
rect 22554 10548 22560 10600
rect 22612 10548 22618 10600
rect 22756 10588 22784 10628
rect 23382 10616 23388 10668
rect 23440 10616 23446 10668
rect 23842 10616 23848 10668
rect 23900 10656 23906 10668
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23900 10628 24225 10656
rect 23900 10616 23906 10628
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 23474 10588 23480 10600
rect 22756 10560 23480 10588
rect 23474 10548 23480 10560
rect 23532 10548 23538 10600
rect 23569 10591 23627 10597
rect 23569 10557 23581 10591
rect 23615 10557 23627 10591
rect 23569 10551 23627 10557
rect 15252 10492 16344 10520
rect 15252 10480 15258 10492
rect 22646 10480 22652 10532
rect 22704 10520 22710 10532
rect 23584 10520 23612 10551
rect 22704 10492 23612 10520
rect 22704 10480 22710 10492
rect 5442 10452 5448 10464
rect 4816 10424 5448 10452
rect 5442 10412 5448 10424
rect 5500 10412 5506 10464
rect 5810 10412 5816 10464
rect 5868 10452 5874 10464
rect 6457 10455 6515 10461
rect 6457 10452 6469 10455
rect 5868 10424 6469 10452
rect 5868 10412 5874 10424
rect 6457 10421 6469 10424
rect 6503 10421 6515 10455
rect 6457 10415 6515 10421
rect 6825 10455 6883 10461
rect 6825 10421 6837 10455
rect 6871 10452 6883 10455
rect 7282 10452 7288 10464
rect 6871 10424 7288 10452
rect 6871 10421 6883 10424
rect 6825 10415 6883 10421
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7745 10455 7803 10461
rect 7745 10421 7757 10455
rect 7791 10452 7803 10455
rect 7834 10452 7840 10464
rect 7791 10424 7840 10452
rect 7791 10421 7803 10424
rect 7745 10415 7803 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 7926 10412 7932 10464
rect 7984 10412 7990 10464
rect 13354 10412 13360 10464
rect 13412 10412 13418 10464
rect 21910 10412 21916 10464
rect 21968 10412 21974 10464
rect 22830 10412 22836 10464
rect 22888 10452 22894 10464
rect 23017 10455 23075 10461
rect 23017 10452 23029 10455
rect 22888 10424 23029 10452
rect 22888 10412 22894 10424
rect 23017 10421 23029 10424
rect 23063 10421 23075 10455
rect 23017 10415 23075 10421
rect 1104 10362 24840 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 20214 10362
rect 20266 10310 20278 10362
rect 20330 10310 20342 10362
rect 20394 10310 20406 10362
rect 20458 10310 20470 10362
rect 20522 10310 24840 10362
rect 1104 10288 24840 10310
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 4249 10251 4307 10257
rect 4249 10248 4261 10251
rect 2004 10220 4261 10248
rect 2004 10208 2010 10220
rect 4249 10217 4261 10220
rect 4295 10217 4307 10251
rect 4249 10211 4307 10217
rect 1949 10115 2007 10121
rect 1949 10081 1961 10115
rect 1995 10112 2007 10115
rect 2498 10112 2504 10124
rect 1995 10084 2504 10112
rect 1995 10081 2007 10084
rect 1949 10075 2007 10081
rect 2498 10072 2504 10084
rect 2556 10072 2562 10124
rect 1486 10004 1492 10056
rect 1544 10044 1550 10056
rect 1673 10047 1731 10053
rect 1673 10044 1685 10047
rect 1544 10016 1685 10044
rect 1544 10004 1550 10016
rect 1673 10013 1685 10016
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 2958 9936 2964 9988
rect 3016 9936 3022 9988
rect 4264 9976 4292 10211
rect 4706 10208 4712 10260
rect 4764 10248 4770 10260
rect 4893 10251 4951 10257
rect 4893 10248 4905 10251
rect 4764 10220 4905 10248
rect 4764 10208 4770 10220
rect 4893 10217 4905 10220
rect 4939 10217 4951 10251
rect 4893 10211 4951 10217
rect 5074 10208 5080 10260
rect 5132 10208 5138 10260
rect 5350 10208 5356 10260
rect 5408 10208 5414 10260
rect 7282 10208 7288 10260
rect 7340 10248 7346 10260
rect 8570 10248 8576 10260
rect 7340 10220 8576 10248
rect 7340 10208 7346 10220
rect 8570 10208 8576 10220
rect 8628 10208 8634 10260
rect 12618 10208 12624 10260
rect 12676 10208 12682 10260
rect 13262 10208 13268 10260
rect 13320 10248 13326 10260
rect 13357 10251 13415 10257
rect 13357 10248 13369 10251
rect 13320 10220 13369 10248
rect 13320 10208 13326 10220
rect 13357 10217 13369 10220
rect 13403 10217 13415 10251
rect 13357 10211 13415 10217
rect 15013 10251 15071 10257
rect 15013 10217 15025 10251
rect 15059 10248 15071 10251
rect 17310 10248 17316 10260
rect 15059 10220 17316 10248
rect 15059 10217 15071 10220
rect 15013 10211 15071 10217
rect 17310 10208 17316 10220
rect 17368 10208 17374 10260
rect 17586 10208 17592 10260
rect 17644 10248 17650 10260
rect 17681 10251 17739 10257
rect 17681 10248 17693 10251
rect 17644 10220 17693 10248
rect 17644 10208 17650 10220
rect 17681 10217 17693 10220
rect 17727 10217 17739 10251
rect 17681 10211 17739 10217
rect 17865 10251 17923 10257
rect 17865 10217 17877 10251
rect 17911 10248 17923 10251
rect 18046 10248 18052 10260
rect 17911 10220 18052 10248
rect 17911 10217 17923 10220
rect 17865 10211 17923 10217
rect 6546 10180 6552 10192
rect 4448 10152 6552 10180
rect 4448 10053 4476 10152
rect 6546 10140 6552 10152
rect 6604 10140 6610 10192
rect 13173 10183 13231 10189
rect 13173 10149 13185 10183
rect 13219 10180 13231 10183
rect 13538 10180 13544 10192
rect 13219 10152 13544 10180
rect 13219 10149 13231 10152
rect 13173 10143 13231 10149
rect 13538 10140 13544 10152
rect 13596 10140 13602 10192
rect 14737 10183 14795 10189
rect 14737 10149 14749 10183
rect 14783 10180 14795 10183
rect 15654 10180 15660 10192
rect 14783 10152 15660 10180
rect 14783 10149 14795 10152
rect 14737 10143 14795 10149
rect 15654 10140 15660 10152
rect 15712 10140 15718 10192
rect 17696 10180 17724 10211
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18325 10251 18383 10257
rect 18325 10217 18337 10251
rect 18371 10217 18383 10251
rect 18325 10211 18383 10217
rect 18340 10180 18368 10211
rect 18506 10208 18512 10260
rect 18564 10208 18570 10260
rect 22646 10248 22652 10260
rect 20824 10220 22652 10248
rect 17696 10152 18368 10180
rect 5810 10072 5816 10124
rect 5868 10072 5874 10124
rect 7558 10112 7564 10124
rect 6564 10084 7564 10112
rect 4433 10047 4491 10053
rect 4433 10013 4445 10047
rect 4479 10013 4491 10047
rect 4433 10007 4491 10013
rect 5537 10047 5595 10053
rect 5537 10013 5549 10047
rect 5583 10013 5595 10047
rect 5537 10007 5595 10013
rect 4709 9979 4767 9985
rect 4709 9976 4721 9979
rect 4264 9948 4721 9976
rect 4709 9945 4721 9948
rect 4755 9945 4767 9979
rect 4709 9939 4767 9945
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 3421 9911 3479 9917
rect 3421 9908 3433 9911
rect 2924 9880 3433 9908
rect 2924 9868 2930 9880
rect 3421 9877 3433 9880
rect 3467 9877 3479 9911
rect 3421 9871 3479 9877
rect 4614 9868 4620 9920
rect 4672 9908 4678 9920
rect 4909 9911 4967 9917
rect 4909 9908 4921 9911
rect 4672 9880 4921 9908
rect 4672 9868 4678 9880
rect 4909 9877 4921 9880
rect 4955 9877 4967 9911
rect 4909 9871 4967 9877
rect 5442 9868 5448 9920
rect 5500 9908 5506 9920
rect 5552 9908 5580 10007
rect 5626 10004 5632 10056
rect 5684 10004 5690 10056
rect 5721 10047 5779 10053
rect 5721 10013 5733 10047
rect 5767 10044 5779 10047
rect 6564 10044 6592 10084
rect 7558 10072 7564 10084
rect 7616 10112 7622 10124
rect 8665 10115 8723 10121
rect 8665 10112 8677 10115
rect 7616 10084 8677 10112
rect 7616 10072 7622 10084
rect 8665 10081 8677 10084
rect 8711 10081 8723 10115
rect 8665 10075 8723 10081
rect 10318 10072 10324 10124
rect 10376 10112 10382 10124
rect 10376 10084 10640 10112
rect 10376 10072 10382 10084
rect 5767 10016 6592 10044
rect 5767 10013 5779 10016
rect 5721 10007 5779 10013
rect 6638 10004 6644 10056
rect 6696 10004 6702 10056
rect 9033 10047 9091 10053
rect 9033 10013 9045 10047
rect 9079 10013 9091 10047
rect 10612 10044 10640 10084
rect 10870 10072 10876 10124
rect 10928 10112 10934 10124
rect 13354 10112 13360 10124
rect 10928 10084 13360 10112
rect 10928 10072 10934 10084
rect 11716 10053 11744 10084
rect 13354 10072 13360 10084
rect 13412 10072 13418 10124
rect 13630 10072 13636 10124
rect 13688 10112 13694 10124
rect 13688 10084 14872 10112
rect 13688 10072 13694 10084
rect 11241 10047 11299 10053
rect 11241 10044 11253 10047
rect 10612 10016 11253 10044
rect 9033 10007 9091 10013
rect 11241 10013 11253 10016
rect 11287 10013 11299 10047
rect 11241 10007 11299 10013
rect 11701 10047 11759 10053
rect 11701 10013 11713 10047
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 12069 10047 12127 10053
rect 12069 10013 12081 10047
rect 12115 10013 12127 10047
rect 12069 10007 12127 10013
rect 6914 9936 6920 9988
rect 6972 9936 6978 9988
rect 7926 9936 7932 9988
rect 7984 9936 7990 9988
rect 9048 9976 9076 10007
rect 9214 9976 9220 9988
rect 9048 9948 9220 9976
rect 9214 9936 9220 9948
rect 9272 9936 9278 9988
rect 9306 9936 9312 9988
rect 9364 9936 9370 9988
rect 9766 9936 9772 9988
rect 9824 9936 9830 9988
rect 10962 9936 10968 9988
rect 11020 9976 11026 9988
rect 12084 9976 12112 10007
rect 12894 10004 12900 10056
rect 12952 10004 12958 10056
rect 13998 10004 14004 10056
rect 14056 10044 14062 10056
rect 14844 10053 14872 10084
rect 15286 10072 15292 10124
rect 15344 10112 15350 10124
rect 15344 10084 16344 10112
rect 15344 10072 15350 10084
rect 14553 10047 14611 10053
rect 14553 10044 14565 10047
rect 14056 10016 14565 10044
rect 14056 10004 14062 10016
rect 14553 10013 14565 10016
rect 14599 10013 14611 10047
rect 14553 10007 14611 10013
rect 14645 10047 14703 10053
rect 14645 10013 14657 10047
rect 14691 10044 14703 10047
rect 14829 10047 14887 10053
rect 14691 10016 14780 10044
rect 14691 10013 14703 10016
rect 14645 10007 14703 10013
rect 13541 9979 13599 9985
rect 11020 9948 12434 9976
rect 11020 9936 11026 9948
rect 7098 9908 7104 9920
rect 5500 9880 7104 9908
rect 5500 9868 5506 9880
rect 7098 9868 7104 9880
rect 7156 9868 7162 9920
rect 10226 9868 10232 9920
rect 10284 9908 10290 9920
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10284 9880 10793 9908
rect 10284 9868 10290 9880
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 12406 9908 12434 9948
rect 13541 9945 13553 9979
rect 13587 9976 13599 9979
rect 13814 9976 13820 9988
rect 13587 9948 13820 9976
rect 13587 9945 13599 9948
rect 13541 9939 13599 9945
rect 13814 9936 13820 9948
rect 13872 9936 13878 9988
rect 12618 9908 12624 9920
rect 12406 9880 12624 9908
rect 10781 9871 10839 9877
rect 12618 9868 12624 9880
rect 12676 9868 12682 9920
rect 12894 9868 12900 9920
rect 12952 9908 12958 9920
rect 13331 9911 13389 9917
rect 13331 9908 13343 9911
rect 12952 9880 13343 9908
rect 12952 9868 12958 9880
rect 13331 9877 13343 9880
rect 13377 9877 13389 9911
rect 14752 9908 14780 10016
rect 14829 10013 14841 10047
rect 14875 10013 14887 10047
rect 14829 10007 14887 10013
rect 15378 10004 15384 10056
rect 15436 10004 15442 10056
rect 16316 10053 16344 10084
rect 19886 10072 19892 10124
rect 19944 10112 19950 10124
rect 20824 10121 20852 10220
rect 22646 10208 22652 10220
rect 22704 10208 22710 10260
rect 23290 10208 23296 10260
rect 23348 10248 23354 10260
rect 23385 10251 23443 10257
rect 23385 10248 23397 10251
rect 23348 10220 23397 10248
rect 23348 10208 23354 10220
rect 23385 10217 23397 10220
rect 23431 10217 23443 10251
rect 23385 10211 23443 10217
rect 24026 10208 24032 10260
rect 24084 10248 24090 10260
rect 24121 10251 24179 10257
rect 24121 10248 24133 10251
rect 24084 10220 24133 10248
rect 24084 10208 24090 10220
rect 24121 10217 24133 10220
rect 24167 10217 24179 10251
rect 24121 10211 24179 10217
rect 20809 10115 20867 10121
rect 20809 10112 20821 10115
rect 19944 10084 20821 10112
rect 19944 10072 19950 10084
rect 20809 10081 20821 10084
rect 20855 10081 20867 10115
rect 20809 10075 20867 10081
rect 21637 10115 21695 10121
rect 21637 10081 21649 10115
rect 21683 10112 21695 10115
rect 22462 10112 22468 10124
rect 21683 10084 22468 10112
rect 21683 10081 21695 10084
rect 21637 10075 21695 10081
rect 22462 10072 22468 10084
rect 22520 10112 22526 10124
rect 22922 10112 22928 10124
rect 22520 10084 22928 10112
rect 22520 10072 22526 10084
rect 22922 10072 22928 10084
rect 22980 10072 22986 10124
rect 23106 10072 23112 10124
rect 23164 10112 23170 10124
rect 23164 10084 23796 10112
rect 23164 10072 23170 10084
rect 16307 10047 16365 10053
rect 16307 10013 16319 10047
rect 16353 10013 16365 10047
rect 16307 10007 16365 10013
rect 16485 10047 16543 10053
rect 16485 10013 16497 10047
rect 16531 10044 16543 10047
rect 16666 10044 16672 10056
rect 16531 10016 16672 10044
rect 16531 10013 16543 10016
rect 16485 10007 16543 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 20622 10004 20628 10056
rect 20680 10044 20686 10056
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 20680 10016 20729 10044
rect 20680 10004 20686 10016
rect 20717 10013 20729 10016
rect 20763 10013 20775 10047
rect 20717 10007 20775 10013
rect 23566 10004 23572 10056
rect 23624 10044 23630 10056
rect 23768 10053 23796 10084
rect 23661 10047 23719 10053
rect 23661 10044 23673 10047
rect 23624 10016 23673 10044
rect 23624 10004 23630 10016
rect 23661 10013 23673 10016
rect 23707 10013 23719 10047
rect 23661 10007 23719 10013
rect 23753 10047 23811 10053
rect 23753 10013 23765 10047
rect 23799 10013 23811 10047
rect 23753 10007 23811 10013
rect 23937 10047 23995 10053
rect 23937 10013 23949 10047
rect 23983 10013 23995 10047
rect 23937 10007 23995 10013
rect 15286 9936 15292 9988
rect 15344 9976 15350 9988
rect 16393 9979 16451 9985
rect 16393 9976 16405 9979
rect 15344 9948 16405 9976
rect 15344 9936 15350 9948
rect 16393 9945 16405 9948
rect 16439 9945 16451 9979
rect 16393 9939 16451 9945
rect 17494 9936 17500 9988
rect 17552 9976 17558 9988
rect 18141 9979 18199 9985
rect 18141 9976 18153 9979
rect 17552 9948 18153 9976
rect 17552 9936 17558 9948
rect 18141 9945 18153 9948
rect 18187 9976 18199 9979
rect 19794 9976 19800 9988
rect 18187 9948 19800 9976
rect 18187 9945 18199 9948
rect 18141 9939 18199 9945
rect 19794 9936 19800 9948
rect 19852 9936 19858 9988
rect 21542 9976 21548 9988
rect 20640 9948 21548 9976
rect 15746 9908 15752 9920
rect 14752 9880 15752 9908
rect 13331 9871 13389 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 17678 9868 17684 9920
rect 17736 9917 17742 9920
rect 17736 9911 17755 9917
rect 17743 9908 17755 9911
rect 18341 9911 18399 9917
rect 18341 9908 18353 9911
rect 17743 9880 18353 9908
rect 17743 9877 17755 9880
rect 17736 9871 17755 9877
rect 18341 9877 18353 9880
rect 18387 9908 18399 9911
rect 19610 9908 19616 9920
rect 18387 9880 19616 9908
rect 18387 9877 18399 9880
rect 18341 9871 18399 9877
rect 17736 9868 17742 9871
rect 19610 9868 19616 9880
rect 19668 9868 19674 9920
rect 19978 9868 19984 9920
rect 20036 9908 20042 9920
rect 20640 9917 20668 9948
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 21910 9936 21916 9988
rect 21968 9936 21974 9988
rect 22646 9936 22652 9988
rect 22704 9936 22710 9988
rect 23952 9976 23980 10007
rect 23308 9948 23980 9976
rect 20257 9911 20315 9917
rect 20257 9908 20269 9911
rect 20036 9880 20269 9908
rect 20036 9868 20042 9880
rect 20257 9877 20269 9880
rect 20303 9877 20315 9911
rect 20257 9871 20315 9877
rect 20625 9911 20683 9917
rect 20625 9877 20637 9911
rect 20671 9877 20683 9911
rect 20625 9871 20683 9877
rect 21361 9911 21419 9917
rect 21361 9877 21373 9911
rect 21407 9908 21419 9911
rect 21634 9908 21640 9920
rect 21407 9880 21640 9908
rect 21407 9877 21419 9880
rect 21361 9871 21419 9877
rect 21634 9868 21640 9880
rect 21692 9868 21698 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 23308 9908 23336 9948
rect 22152 9880 23336 9908
rect 22152 9868 22158 9880
rect 1104 9818 24840 9840
rect 1104 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 24214 9818
rect 24266 9766 24278 9818
rect 24330 9766 24342 9818
rect 24394 9766 24406 9818
rect 24458 9766 24470 9818
rect 24522 9766 24840 9818
rect 1104 9744 24840 9766
rect 2225 9707 2283 9713
rect 2225 9673 2237 9707
rect 2271 9673 2283 9707
rect 2225 9667 2283 9673
rect 1854 9596 1860 9648
rect 1912 9596 1918 9648
rect 2038 9596 2044 9648
rect 2096 9645 2102 9648
rect 2096 9639 2115 9645
rect 2103 9605 2115 9639
rect 2240 9636 2268 9667
rect 2498 9664 2504 9716
rect 2556 9664 2562 9716
rect 2866 9664 2872 9716
rect 2924 9664 2930 9716
rect 6914 9664 6920 9716
rect 6972 9664 6978 9716
rect 7466 9664 7472 9716
rect 7524 9704 7530 9716
rect 9030 9704 9036 9716
rect 7524 9676 9036 9704
rect 7524 9664 7530 9676
rect 9030 9664 9036 9676
rect 9088 9664 9094 9716
rect 10226 9664 10232 9716
rect 10284 9704 10290 9716
rect 10284 9676 12572 9704
rect 10284 9664 10290 9676
rect 2958 9636 2964 9648
rect 2240 9608 2964 9636
rect 2096 9599 2115 9605
rect 2096 9596 2102 9599
rect 2958 9596 2964 9608
rect 3016 9596 3022 9648
rect 4982 9596 4988 9648
rect 5040 9596 5046 9648
rect 6270 9596 6276 9648
rect 6328 9636 6334 9648
rect 6328 9608 6684 9636
rect 6328 9596 6334 9608
rect 3234 9568 3240 9580
rect 2976 9540 3240 9568
rect 2976 9509 3004 9540
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 6546 9568 6552 9580
rect 6503 9540 6552 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 6656 9577 6684 9608
rect 8938 9596 8944 9648
rect 8996 9596 9002 9648
rect 9122 9596 9128 9648
rect 9180 9645 9186 9648
rect 9180 9639 9199 9645
rect 9187 9636 9199 9639
rect 9585 9639 9643 9645
rect 9585 9636 9597 9639
rect 9187 9608 9597 9636
rect 9187 9605 9199 9608
rect 9180 9599 9199 9605
rect 9585 9605 9597 9608
rect 9631 9605 9643 9639
rect 9585 9599 9643 9605
rect 9180 9596 9186 9599
rect 6641 9571 6699 9577
rect 6641 9537 6653 9571
rect 6687 9537 6699 9571
rect 6641 9531 6699 9537
rect 7098 9528 7104 9580
rect 7156 9568 7162 9580
rect 7466 9568 7472 9580
rect 7156 9540 7472 9568
rect 7156 9528 7162 9540
rect 7466 9528 7472 9540
rect 7524 9528 7530 9580
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 9858 9568 9864 9580
rect 9815 9540 9864 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 9858 9528 9864 9540
rect 9916 9528 9922 9580
rect 10318 9528 10324 9580
rect 10376 9568 10382 9580
rect 10781 9571 10839 9577
rect 10781 9568 10793 9571
rect 10376 9540 10793 9568
rect 10376 9528 10382 9540
rect 10781 9537 10793 9540
rect 10827 9537 10839 9571
rect 10781 9531 10839 9537
rect 10870 9528 10876 9580
rect 10928 9528 10934 9580
rect 10965 9571 11023 9577
rect 10965 9537 10977 9571
rect 11011 9537 11023 9571
rect 10965 9531 11023 9537
rect 2961 9503 3019 9509
rect 2961 9469 2973 9503
rect 3007 9469 3019 9503
rect 2961 9463 3019 9469
rect 3142 9460 3148 9512
rect 3200 9460 3206 9512
rect 4249 9503 4307 9509
rect 4249 9469 4261 9503
rect 4295 9469 4307 9503
rect 4249 9463 4307 9469
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 5258 9500 5264 9512
rect 4571 9472 5264 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 1486 9392 1492 9444
rect 1544 9432 1550 9444
rect 4264 9432 4292 9463
rect 5258 9460 5264 9472
rect 5316 9460 5322 9512
rect 5902 9460 5908 9512
rect 5960 9500 5966 9512
rect 5997 9503 6055 9509
rect 5997 9500 6009 9503
rect 5960 9472 6009 9500
rect 5960 9460 5966 9472
rect 5997 9469 6009 9472
rect 6043 9500 6055 9503
rect 6362 9500 6368 9512
rect 6043 9472 6368 9500
rect 6043 9469 6055 9472
rect 5997 9463 6055 9469
rect 6362 9460 6368 9472
rect 6420 9460 6426 9512
rect 7377 9503 7435 9509
rect 7377 9469 7389 9503
rect 7423 9500 7435 9503
rect 7558 9500 7564 9512
rect 7423 9472 7564 9500
rect 7423 9469 7435 9472
rect 7377 9463 7435 9469
rect 7558 9460 7564 9472
rect 7616 9500 7622 9512
rect 7834 9500 7840 9512
rect 7616 9472 7840 9500
rect 7616 9460 7622 9472
rect 7834 9460 7840 9472
rect 7892 9460 7898 9512
rect 10410 9460 10416 9512
rect 10468 9500 10474 9512
rect 10980 9500 11008 9531
rect 11514 9528 11520 9580
rect 11572 9568 11578 9580
rect 11793 9571 11851 9577
rect 11793 9568 11805 9571
rect 11572 9540 11805 9568
rect 11572 9528 11578 9540
rect 11793 9537 11805 9540
rect 11839 9537 11851 9571
rect 11793 9531 11851 9537
rect 11885 9571 11943 9577
rect 11885 9537 11897 9571
rect 11931 9568 11943 9571
rect 12066 9568 12072 9580
rect 11931 9540 12072 9568
rect 11931 9537 11943 9540
rect 11885 9531 11943 9537
rect 12066 9528 12072 9540
rect 12124 9528 12130 9580
rect 10468 9472 11008 9500
rect 10468 9460 10474 9472
rect 6638 9432 6644 9444
rect 1544 9404 4292 9432
rect 1544 9392 1550 9404
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 2130 9364 2136 9376
rect 2087 9336 2136 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 2130 9324 2136 9336
rect 2188 9324 2194 9376
rect 4264 9364 4292 9404
rect 5552 9404 6644 9432
rect 5552 9364 5580 9404
rect 6638 9392 6644 9404
rect 6696 9392 6702 9444
rect 9309 9435 9367 9441
rect 9309 9401 9321 9435
rect 9355 9432 9367 9435
rect 9766 9432 9772 9444
rect 9355 9404 9772 9432
rect 9355 9401 9367 9404
rect 9309 9395 9367 9401
rect 9766 9392 9772 9404
rect 9824 9392 9830 9444
rect 4264 9336 5580 9364
rect 5810 9324 5816 9376
rect 5868 9364 5874 9376
rect 6457 9367 6515 9373
rect 6457 9364 6469 9367
rect 5868 9336 6469 9364
rect 5868 9324 5874 9336
rect 6457 9333 6469 9336
rect 6503 9333 6515 9367
rect 6457 9327 6515 9333
rect 7285 9367 7343 9373
rect 7285 9333 7297 9367
rect 7331 9364 7343 9367
rect 7374 9364 7380 9376
rect 7331 9336 7380 9364
rect 7331 9333 7343 9336
rect 7285 9327 7343 9333
rect 7374 9324 7380 9336
rect 7432 9324 7438 9376
rect 8754 9324 8760 9376
rect 8812 9364 8818 9376
rect 9125 9367 9183 9373
rect 9125 9364 9137 9367
rect 8812 9336 9137 9364
rect 8812 9324 8818 9336
rect 9125 9333 9137 9336
rect 9171 9333 9183 9367
rect 9125 9327 9183 9333
rect 10502 9324 10508 9376
rect 10560 9324 10566 9376
rect 10980 9364 11008 9472
rect 11238 9460 11244 9512
rect 11296 9460 11302 9512
rect 12360 9509 12388 9676
rect 12544 9636 12572 9676
rect 12618 9664 12624 9716
rect 12676 9664 12682 9716
rect 13262 9704 13268 9716
rect 12728 9676 13268 9704
rect 12728 9636 12756 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 15565 9707 15623 9713
rect 15565 9673 15577 9707
rect 15611 9704 15623 9707
rect 15746 9704 15752 9716
rect 15611 9676 15752 9704
rect 15611 9673 15623 9676
rect 15565 9667 15623 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 18953 9707 19011 9713
rect 18953 9673 18965 9707
rect 18999 9704 19011 9707
rect 22186 9704 22192 9716
rect 18999 9673 19012 9704
rect 18953 9667 19012 9673
rect 14642 9636 14648 9648
rect 12544 9608 12756 9636
rect 14384 9608 14648 9636
rect 12710 9528 12716 9580
rect 12768 9568 12774 9580
rect 12989 9571 13047 9577
rect 12989 9568 13001 9571
rect 12768 9540 13001 9568
rect 12768 9528 12774 9540
rect 12989 9537 13001 9540
rect 13035 9537 13047 9571
rect 12989 9531 13047 9537
rect 13998 9528 14004 9580
rect 14056 9528 14062 9580
rect 14384 9577 14412 9608
rect 14642 9596 14648 9608
rect 14700 9636 14706 9648
rect 17129 9639 17187 9645
rect 14700 9608 15608 9636
rect 14700 9596 14706 9608
rect 14369 9571 14427 9577
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 14458 9528 14464 9580
rect 14516 9528 14522 9580
rect 14921 9571 14979 9577
rect 14921 9537 14933 9571
rect 14967 9568 14979 9571
rect 15286 9568 15292 9580
rect 14967 9540 15292 9568
rect 14967 9537 14979 9540
rect 14921 9531 14979 9537
rect 15286 9528 15292 9540
rect 15344 9528 15350 9580
rect 15580 9577 15608 9608
rect 17129 9605 17141 9639
rect 17175 9636 17187 9639
rect 18046 9636 18052 9648
rect 17175 9608 18052 9636
rect 17175 9605 17187 9608
rect 17129 9599 17187 9605
rect 18046 9596 18052 9608
rect 18104 9636 18110 9648
rect 18233 9639 18291 9645
rect 18233 9636 18245 9639
rect 18104 9608 18245 9636
rect 18104 9596 18110 9608
rect 18233 9605 18245 9608
rect 18279 9605 18291 9639
rect 18233 9599 18291 9605
rect 18598 9596 18604 9648
rect 18656 9636 18662 9648
rect 18984 9636 19012 9667
rect 20364 9676 22192 9704
rect 18656 9608 19012 9636
rect 19153 9639 19211 9645
rect 18656 9596 18662 9608
rect 19153 9605 19165 9639
rect 19199 9605 19211 9639
rect 20364 9636 20392 9676
rect 22186 9664 22192 9676
rect 22244 9704 22250 9716
rect 22462 9704 22468 9716
rect 22244 9676 22468 9704
rect 22244 9664 22250 9676
rect 22462 9664 22468 9676
rect 22520 9664 22526 9716
rect 22554 9664 22560 9716
rect 22612 9704 22618 9716
rect 23750 9704 23756 9716
rect 22612 9676 23756 9704
rect 22612 9664 22618 9676
rect 23750 9664 23756 9676
rect 23808 9664 23814 9716
rect 22094 9645 22100 9648
rect 19153 9599 19211 9605
rect 19720 9608 20392 9636
rect 22081 9639 22100 9645
rect 15565 9571 15623 9577
rect 15565 9537 15577 9571
rect 15611 9537 15623 9571
rect 15565 9531 15623 9537
rect 12345 9503 12403 9509
rect 12345 9469 12357 9503
rect 12391 9469 12403 9503
rect 12345 9463 12403 9469
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9469 15255 9503
rect 15197 9463 15255 9469
rect 11149 9435 11207 9441
rect 11149 9401 11161 9435
rect 11195 9432 11207 9435
rect 12894 9432 12900 9444
rect 11195 9404 12900 9432
rect 11195 9401 11207 9404
rect 11149 9395 11207 9401
rect 12894 9392 12900 9404
rect 12952 9392 12958 9444
rect 13909 9435 13967 9441
rect 13909 9432 13921 9435
rect 13188 9404 13921 9432
rect 12253 9367 12311 9373
rect 12253 9364 12265 9367
rect 10980 9336 12265 9364
rect 12253 9333 12265 9336
rect 12299 9364 12311 9367
rect 13188 9364 13216 9404
rect 13909 9401 13921 9404
rect 13955 9401 13967 9435
rect 13909 9395 13967 9401
rect 14737 9435 14795 9441
rect 14737 9401 14749 9435
rect 14783 9432 14795 9435
rect 15102 9432 15108 9444
rect 14783 9404 15108 9432
rect 14783 9401 14795 9404
rect 14737 9395 14795 9401
rect 15102 9392 15108 9404
rect 15160 9392 15166 9444
rect 12299 9336 13216 9364
rect 12299 9333 12311 9336
rect 12253 9327 12311 9333
rect 13446 9324 13452 9376
rect 13504 9324 13510 9376
rect 13722 9324 13728 9376
rect 13780 9364 13786 9376
rect 14829 9367 14887 9373
rect 14829 9364 14841 9367
rect 13780 9336 14841 9364
rect 13780 9324 13786 9336
rect 14829 9333 14841 9336
rect 14875 9364 14887 9367
rect 15222 9364 15250 9463
rect 15580 9432 15608 9531
rect 15654 9528 15660 9580
rect 15712 9568 15718 9580
rect 16025 9571 16083 9577
rect 16025 9568 16037 9571
rect 15712 9540 16037 9568
rect 15712 9528 15718 9540
rect 16025 9537 16037 9540
rect 16071 9537 16083 9571
rect 16025 9531 16083 9537
rect 16114 9528 16120 9580
rect 16172 9568 16178 9580
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 16172 9540 16221 9568
rect 16172 9528 16178 9540
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 18141 9571 18199 9577
rect 18141 9537 18153 9571
rect 18187 9568 18199 9571
rect 18690 9568 18696 9580
rect 18187 9540 18696 9568
rect 18187 9537 18199 9540
rect 18141 9531 18199 9537
rect 18690 9528 18696 9540
rect 18748 9528 18754 9580
rect 18874 9528 18880 9580
rect 18932 9568 18938 9580
rect 19168 9568 19196 9599
rect 18932 9540 19196 9568
rect 18932 9528 18938 9540
rect 19334 9528 19340 9580
rect 19392 9568 19398 9580
rect 19720 9577 19748 9608
rect 22081 9605 22093 9639
rect 22081 9599 22100 9605
rect 22094 9596 22100 9599
rect 22152 9596 22158 9648
rect 22281 9639 22339 9645
rect 22281 9605 22293 9639
rect 22327 9605 22339 9639
rect 22281 9599 22339 9605
rect 19705 9571 19763 9577
rect 19705 9568 19717 9571
rect 19392 9540 19717 9568
rect 19392 9528 19398 9540
rect 19705 9537 19717 9540
rect 19751 9537 19763 9571
rect 19705 9531 19763 9537
rect 15746 9460 15752 9512
rect 15804 9460 15810 9512
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 15896 9472 17233 9500
rect 15896 9460 15902 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 17405 9503 17463 9509
rect 17405 9469 17417 9503
rect 17451 9500 17463 9503
rect 18230 9500 18236 9512
rect 17451 9472 18236 9500
rect 17451 9469 17463 9472
rect 17405 9463 17463 9469
rect 18230 9460 18236 9472
rect 18288 9500 18294 9512
rect 18325 9503 18383 9509
rect 18325 9500 18337 9503
rect 18288 9472 18337 9500
rect 18288 9460 18294 9472
rect 18325 9469 18337 9472
rect 18371 9469 18383 9503
rect 18325 9463 18383 9469
rect 19978 9460 19984 9512
rect 20036 9460 20042 9512
rect 16117 9435 16175 9441
rect 16117 9432 16129 9435
rect 15580 9404 16129 9432
rect 16117 9401 16129 9404
rect 16163 9401 16175 9435
rect 21100 9432 21128 9554
rect 21358 9528 21364 9580
rect 21416 9568 21422 9580
rect 22296 9568 22324 9599
rect 21416 9540 22324 9568
rect 22480 9568 22508 9664
rect 22830 9596 22836 9648
rect 22888 9596 22894 9648
rect 23474 9596 23480 9648
rect 23532 9596 23538 9648
rect 22557 9571 22615 9577
rect 22557 9568 22569 9571
rect 22480 9540 22569 9568
rect 21416 9528 21422 9540
rect 22557 9537 22569 9540
rect 22603 9537 22615 9571
rect 22557 9531 22615 9537
rect 21453 9503 21511 9509
rect 21453 9469 21465 9503
rect 21499 9500 21511 9503
rect 21542 9500 21548 9512
rect 21499 9472 21548 9500
rect 21499 9469 21511 9472
rect 21453 9463 21511 9469
rect 21542 9460 21548 9472
rect 21600 9460 21606 9512
rect 23382 9460 23388 9512
rect 23440 9500 23446 9512
rect 24305 9503 24363 9509
rect 24305 9500 24317 9503
rect 23440 9472 24317 9500
rect 23440 9460 23446 9472
rect 24305 9469 24317 9472
rect 24351 9469 24363 9503
rect 24305 9463 24363 9469
rect 21913 9435 21971 9441
rect 21913 9432 21925 9435
rect 21100 9404 21925 9432
rect 16117 9395 16175 9401
rect 21913 9401 21925 9404
rect 21959 9401 21971 9435
rect 21913 9395 21971 9401
rect 14875 9336 15250 9364
rect 14875 9333 14887 9336
rect 14829 9327 14887 9333
rect 16574 9324 16580 9376
rect 16632 9364 16638 9376
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 16632 9336 16773 9364
rect 16632 9324 16638 9336
rect 16761 9333 16773 9336
rect 16807 9333 16819 9367
rect 16761 9327 16819 9333
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 17773 9367 17831 9373
rect 17773 9364 17785 9367
rect 17276 9336 17785 9364
rect 17276 9324 17282 9336
rect 17773 9333 17785 9336
rect 17819 9333 17831 9367
rect 17773 9327 17831 9333
rect 18782 9324 18788 9376
rect 18840 9324 18846 9376
rect 18966 9324 18972 9376
rect 19024 9364 19030 9376
rect 22097 9367 22155 9373
rect 22097 9364 22109 9367
rect 19024 9336 22109 9364
rect 19024 9324 19030 9336
rect 22097 9333 22109 9336
rect 22143 9364 22155 9367
rect 22278 9364 22284 9376
rect 22143 9336 22284 9364
rect 22143 9333 22155 9336
rect 22097 9327 22155 9333
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 1104 9274 24840 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 20214 9274
rect 20266 9222 20278 9274
rect 20330 9222 20342 9274
rect 20394 9222 20406 9274
rect 20458 9222 20470 9274
rect 20522 9222 24840 9274
rect 1104 9200 24840 9222
rect 4798 9120 4804 9172
rect 4856 9120 4862 9172
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 5258 9120 5264 9172
rect 5316 9120 5322 9172
rect 5350 9120 5356 9172
rect 5408 9160 5414 9172
rect 8389 9163 8447 9169
rect 5408 9132 8340 9160
rect 5408 9120 5414 9132
rect 8018 9092 8024 9104
rect 4632 9064 8024 9092
rect 1486 8916 1492 8968
rect 1544 8956 1550 8968
rect 1581 8959 1639 8965
rect 1581 8956 1593 8959
rect 1544 8928 1593 8956
rect 1544 8916 1550 8928
rect 1581 8925 1593 8928
rect 1627 8925 1639 8959
rect 1581 8919 1639 8925
rect 1857 8891 1915 8897
rect 1857 8857 1869 8891
rect 1903 8857 1915 8891
rect 1857 8851 1915 8857
rect 1872 8820 1900 8851
rect 2130 8848 2136 8900
rect 2188 8888 2194 8900
rect 4632 8897 4660 9064
rect 8018 9052 8024 9064
rect 8076 9052 8082 9104
rect 5626 9024 5632 9036
rect 5552 8996 5632 9024
rect 5442 8916 5448 8968
rect 5500 8916 5506 8968
rect 5552 8965 5580 8996
rect 5626 8984 5632 8996
rect 5684 9024 5690 9036
rect 7009 9027 7067 9033
rect 5684 8996 6776 9024
rect 5684 8984 5690 8996
rect 5810 8965 5816 8968
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8925 5595 8959
rect 5537 8919 5595 8925
rect 5767 8959 5816 8965
rect 5767 8925 5779 8959
rect 5813 8925 5816 8959
rect 5767 8919 5816 8925
rect 5810 8916 5816 8919
rect 5868 8916 5874 8968
rect 5905 8959 5963 8965
rect 5905 8925 5917 8959
rect 5951 8956 5963 8959
rect 6181 8959 6239 8965
rect 6181 8956 6193 8959
rect 5951 8928 6193 8956
rect 5951 8925 5963 8928
rect 5905 8919 5963 8925
rect 6181 8925 6193 8928
rect 6227 8925 6239 8959
rect 6181 8919 6239 8925
rect 6362 8916 6368 8968
rect 6420 8916 6426 8968
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 6641 8959 6699 8965
rect 6641 8956 6653 8959
rect 6512 8928 6653 8956
rect 6512 8916 6518 8928
rect 6641 8925 6653 8928
rect 6687 8925 6699 8959
rect 6748 8956 6776 8996
rect 7009 8993 7021 9027
rect 7055 9024 7067 9027
rect 7190 9024 7196 9036
rect 7055 8996 7196 9024
rect 7055 8993 7067 8996
rect 7009 8987 7067 8993
rect 7190 8984 7196 8996
rect 7248 8984 7254 9036
rect 6748 8928 7420 8956
rect 6641 8919 6699 8925
rect 7392 8900 7420 8928
rect 7466 8916 7472 8968
rect 7524 8916 7530 8968
rect 4617 8891 4675 8897
rect 4617 8888 4629 8891
rect 2188 8860 2346 8888
rect 3252 8860 4629 8888
rect 2188 8848 2194 8860
rect 2222 8820 2228 8832
rect 1872 8792 2228 8820
rect 2222 8780 2228 8792
rect 2280 8780 2286 8832
rect 2498 8780 2504 8832
rect 2556 8820 2562 8832
rect 3252 8820 3280 8860
rect 4617 8857 4629 8860
rect 4663 8857 4675 8891
rect 4617 8851 4675 8857
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 4833 8891 4891 8897
rect 4833 8888 4845 8891
rect 4764 8860 4845 8888
rect 4764 8848 4770 8860
rect 4833 8857 4845 8860
rect 4879 8888 4891 8891
rect 5350 8888 5356 8900
rect 4879 8860 5356 8888
rect 4879 8857 4891 8860
rect 4833 8851 4891 8857
rect 5350 8848 5356 8860
rect 5408 8848 5414 8900
rect 5629 8891 5687 8897
rect 5629 8857 5641 8891
rect 5675 8888 5687 8891
rect 5675 8860 7052 8888
rect 5675 8857 5687 8860
rect 5629 8851 5687 8857
rect 2556 8792 3280 8820
rect 2556 8780 2562 8792
rect 3326 8780 3332 8832
rect 3384 8780 3390 8832
rect 5534 8780 5540 8832
rect 5592 8820 5598 8832
rect 6549 8823 6607 8829
rect 6549 8820 6561 8823
rect 5592 8792 6561 8820
rect 5592 8780 5598 8792
rect 6549 8789 6561 8792
rect 6595 8820 6607 8823
rect 6914 8820 6920 8832
rect 6595 8792 6920 8820
rect 6595 8789 6607 8792
rect 6549 8783 6607 8789
rect 6914 8780 6920 8792
rect 6972 8780 6978 8832
rect 7024 8820 7052 8860
rect 7098 8848 7104 8900
rect 7156 8897 7162 8900
rect 7156 8891 7205 8897
rect 7156 8857 7159 8891
rect 7193 8857 7205 8891
rect 7156 8851 7205 8857
rect 7285 8891 7343 8897
rect 7285 8857 7297 8891
rect 7331 8857 7343 8891
rect 7285 8851 7343 8857
rect 7156 8848 7162 8851
rect 7300 8820 7328 8851
rect 7374 8848 7380 8900
rect 7432 8848 7438 8900
rect 7834 8888 7840 8900
rect 7468 8860 7840 8888
rect 7468 8820 7496 8860
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 8018 8848 8024 8900
rect 8076 8888 8082 8900
rect 8205 8891 8263 8897
rect 8205 8888 8217 8891
rect 8076 8860 8217 8888
rect 8076 8848 8082 8860
rect 8205 8857 8217 8860
rect 8251 8857 8263 8891
rect 8312 8888 8340 9132
rect 8389 9129 8401 9163
rect 8435 9160 8447 9163
rect 8662 9160 8668 9172
rect 8435 9132 8668 9160
rect 8435 9129 8447 9132
rect 8389 9123 8447 9129
rect 8662 9120 8668 9132
rect 8720 9120 8726 9172
rect 9306 9120 9312 9172
rect 9364 9160 9370 9172
rect 9493 9163 9551 9169
rect 9493 9160 9505 9163
rect 9364 9132 9505 9160
rect 9364 9120 9370 9132
rect 9493 9129 9505 9132
rect 9539 9129 9551 9163
rect 9493 9123 9551 9129
rect 9723 9163 9781 9169
rect 9723 9129 9735 9163
rect 9769 9160 9781 9163
rect 10502 9160 10508 9172
rect 9769 9132 10508 9160
rect 9769 9129 9781 9132
rect 9723 9123 9781 9129
rect 10502 9120 10508 9132
rect 10560 9120 10566 9172
rect 18046 9120 18052 9172
rect 18104 9120 18110 9172
rect 18509 9163 18567 9169
rect 18509 9129 18521 9163
rect 18555 9160 18567 9163
rect 18966 9160 18972 9172
rect 18555 9132 18972 9160
rect 18555 9129 18567 9132
rect 18509 9123 18567 9129
rect 18966 9120 18972 9132
rect 19024 9120 19030 9172
rect 19794 9120 19800 9172
rect 19852 9160 19858 9172
rect 22097 9163 22155 9169
rect 19852 9132 21864 9160
rect 19852 9120 19858 9132
rect 9585 9095 9643 9101
rect 9585 9061 9597 9095
rect 9631 9092 9643 9095
rect 13446 9092 13452 9104
rect 9631 9064 13452 9092
rect 9631 9061 9643 9064
rect 9585 9055 9643 9061
rect 13446 9052 13452 9064
rect 13504 9052 13510 9104
rect 10321 9027 10379 9033
rect 10321 9024 10333 9027
rect 9876 8996 10333 9024
rect 9398 8916 9404 8968
rect 9456 8916 9462 8968
rect 9876 8965 9904 8996
rect 10321 8993 10333 8996
rect 10367 8993 10379 9027
rect 10321 8987 10379 8993
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 12161 9027 12219 9033
rect 12161 9024 12173 9027
rect 11296 8996 12173 9024
rect 11296 8984 11302 8996
rect 12161 8993 12173 8996
rect 12207 8993 12219 9027
rect 15194 9024 15200 9036
rect 12161 8987 12219 8993
rect 14108 8996 15200 9024
rect 14108 8968 14136 8996
rect 15194 8984 15200 8996
rect 15252 8984 15258 9036
rect 16301 9027 16359 9033
rect 16301 8993 16313 9027
rect 16347 9024 16359 9027
rect 16942 9024 16948 9036
rect 16347 8996 16948 9024
rect 16347 8993 16359 8996
rect 16301 8987 16359 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 19334 8984 19340 9036
rect 19392 8984 19398 9036
rect 19610 8984 19616 9036
rect 19668 9024 19674 9036
rect 21836 9024 21864 9132
rect 22097 9129 22109 9163
rect 22143 9160 22155 9163
rect 22370 9160 22376 9172
rect 22143 9132 22376 9160
rect 22143 9129 22155 9132
rect 22097 9123 22155 9129
rect 22370 9120 22376 9132
rect 22428 9120 22434 9172
rect 22557 9163 22615 9169
rect 22557 9129 22569 9163
rect 22603 9129 22615 9163
rect 22557 9123 22615 9129
rect 21910 9052 21916 9104
rect 21968 9092 21974 9104
rect 22572 9092 22600 9123
rect 22646 9120 22652 9172
rect 22704 9160 22710 9172
rect 22741 9163 22799 9169
rect 22741 9160 22753 9163
rect 22704 9132 22753 9160
rect 22704 9120 22710 9132
rect 22741 9129 22753 9132
rect 22787 9129 22799 9163
rect 22741 9123 22799 9129
rect 23198 9120 23204 9172
rect 23256 9160 23262 9172
rect 23293 9163 23351 9169
rect 23293 9160 23305 9163
rect 23256 9132 23305 9160
rect 23256 9120 23262 9132
rect 23293 9129 23305 9132
rect 23339 9129 23351 9163
rect 23293 9123 23351 9129
rect 23474 9120 23480 9172
rect 23532 9120 23538 9172
rect 23658 9120 23664 9172
rect 23716 9160 23722 9172
rect 23937 9163 23995 9169
rect 23937 9160 23949 9163
rect 23716 9132 23949 9160
rect 23716 9120 23722 9132
rect 23937 9129 23949 9132
rect 23983 9129 23995 9163
rect 23937 9123 23995 9129
rect 23216 9092 23244 9120
rect 21968 9064 23244 9092
rect 21968 9052 21974 9064
rect 19668 8996 21772 9024
rect 21836 8996 22094 9024
rect 19668 8984 19674 8996
rect 9861 8959 9919 8965
rect 9861 8925 9873 8959
rect 9907 8925 9919 8959
rect 9861 8919 9919 8925
rect 10224 8959 10282 8965
rect 10224 8925 10236 8959
rect 10270 8956 10282 8959
rect 10870 8956 10876 8968
rect 10270 8928 10876 8956
rect 10270 8925 10282 8928
rect 10224 8919 10282 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 10965 8959 11023 8965
rect 10965 8925 10977 8959
rect 11011 8956 11023 8959
rect 11054 8956 11060 8968
rect 11011 8928 11060 8956
rect 11011 8925 11023 8928
rect 10965 8919 11023 8925
rect 11054 8916 11060 8928
rect 11112 8956 11118 8968
rect 11885 8959 11943 8965
rect 11885 8956 11897 8959
rect 11112 8928 11897 8956
rect 11112 8916 11118 8928
rect 11885 8925 11897 8928
rect 11931 8956 11943 8959
rect 12066 8956 12072 8968
rect 11931 8928 12072 8956
rect 11931 8925 11943 8928
rect 11885 8919 11943 8925
rect 12066 8916 12072 8928
rect 12124 8916 12130 8968
rect 12710 8916 12716 8968
rect 12768 8956 12774 8968
rect 13081 8959 13139 8965
rect 13081 8956 13093 8959
rect 12768 8928 13093 8956
rect 12768 8916 12774 8928
rect 13081 8925 13093 8928
rect 13127 8925 13139 8959
rect 14090 8956 14096 8968
rect 13081 8919 13139 8925
rect 13556 8928 14096 8956
rect 8421 8891 8479 8897
rect 8421 8888 8433 8891
rect 8312 8860 8433 8888
rect 8205 8851 8263 8857
rect 8421 8857 8433 8860
rect 8467 8888 8479 8891
rect 8467 8860 9904 8888
rect 8467 8857 8479 8860
rect 8421 8851 8479 8857
rect 9876 8832 9904 8860
rect 10318 8848 10324 8900
rect 10376 8848 10382 8900
rect 10410 8848 10416 8900
rect 10468 8848 10474 8900
rect 10502 8848 10508 8900
rect 10560 8888 10566 8900
rect 10597 8891 10655 8897
rect 10597 8888 10609 8891
rect 10560 8860 10609 8888
rect 10560 8848 10566 8860
rect 10597 8857 10609 8860
rect 10643 8857 10655 8891
rect 10597 8851 10655 8857
rect 11517 8891 11575 8897
rect 11517 8857 11529 8891
rect 11563 8888 11575 8891
rect 13556 8888 13584 8928
rect 14090 8916 14096 8928
rect 14148 8916 14154 8968
rect 14182 8916 14188 8968
rect 14240 8916 14246 8968
rect 21450 8916 21456 8968
rect 21508 8956 21514 8968
rect 21637 8959 21695 8965
rect 21637 8956 21649 8959
rect 21508 8928 21649 8956
rect 21508 8916 21514 8928
rect 21637 8925 21649 8928
rect 21683 8925 21695 8959
rect 21637 8919 21695 8925
rect 11563 8860 13584 8888
rect 13633 8891 13691 8897
rect 11563 8857 11575 8860
rect 11517 8851 11575 8857
rect 13633 8857 13645 8891
rect 13679 8857 13691 8891
rect 13633 8851 13691 8857
rect 7024 8792 7496 8820
rect 7653 8823 7711 8829
rect 7653 8789 7665 8823
rect 7699 8820 7711 8823
rect 7742 8820 7748 8832
rect 7699 8792 7748 8820
rect 7699 8789 7711 8792
rect 7653 8783 7711 8789
rect 7742 8780 7748 8792
rect 7800 8780 7806 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 8754 8820 8760 8832
rect 8619 8792 8760 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 8754 8780 8760 8792
rect 8812 8780 8818 8832
rect 9858 8780 9864 8832
rect 9916 8820 9922 8832
rect 12986 8820 12992 8832
rect 9916 8792 12992 8820
rect 9916 8780 9922 8792
rect 12986 8780 12992 8792
rect 13044 8780 13050 8832
rect 13648 8820 13676 8851
rect 14366 8848 14372 8900
rect 14424 8888 14430 8900
rect 14461 8891 14519 8897
rect 14461 8888 14473 8891
rect 14424 8860 14473 8888
rect 14424 8848 14430 8860
rect 14461 8857 14473 8860
rect 14507 8857 14519 8891
rect 14461 8851 14519 8857
rect 15194 8848 15200 8900
rect 15252 8848 15258 8900
rect 16574 8848 16580 8900
rect 16632 8848 16638 8900
rect 18693 8891 18751 8897
rect 17802 8860 18368 8888
rect 14642 8820 14648 8832
rect 13648 8792 14648 8820
rect 14642 8780 14648 8792
rect 14700 8780 14706 8832
rect 14734 8780 14740 8832
rect 14792 8820 14798 8832
rect 18340 8829 18368 8860
rect 18693 8857 18705 8891
rect 18739 8888 18751 8891
rect 18874 8888 18880 8900
rect 18739 8860 18880 8888
rect 18739 8857 18751 8860
rect 18693 8851 18751 8857
rect 18874 8848 18880 8860
rect 18932 8848 18938 8900
rect 19334 8848 19340 8900
rect 19392 8888 19398 8900
rect 19613 8891 19671 8897
rect 19613 8888 19625 8891
rect 19392 8860 19625 8888
rect 19392 8848 19398 8860
rect 19613 8857 19625 8860
rect 19659 8857 19671 8891
rect 19613 8851 19671 8857
rect 20070 8848 20076 8900
rect 20128 8848 20134 8900
rect 15933 8823 15991 8829
rect 15933 8820 15945 8823
rect 14792 8792 15945 8820
rect 14792 8780 14798 8792
rect 15933 8789 15945 8792
rect 15979 8789 15991 8823
rect 15933 8783 15991 8789
rect 18325 8823 18383 8829
rect 18325 8789 18337 8823
rect 18371 8789 18383 8823
rect 18325 8783 18383 8789
rect 18493 8823 18551 8829
rect 18493 8789 18505 8823
rect 18539 8820 18551 8823
rect 18598 8820 18604 8832
rect 18539 8792 18604 8820
rect 18539 8789 18551 8792
rect 18493 8783 18551 8789
rect 18598 8780 18604 8792
rect 18656 8780 18662 8832
rect 19702 8780 19708 8832
rect 19760 8820 19766 8832
rect 20622 8820 20628 8832
rect 19760 8792 20628 8820
rect 19760 8780 19766 8792
rect 20622 8780 20628 8792
rect 20680 8820 20686 8832
rect 21085 8823 21143 8829
rect 21085 8820 21097 8823
rect 20680 8792 21097 8820
rect 20680 8780 20686 8792
rect 21085 8789 21097 8792
rect 21131 8789 21143 8823
rect 21085 8783 21143 8789
rect 21266 8780 21272 8832
rect 21324 8820 21330 8832
rect 21453 8823 21511 8829
rect 21453 8820 21465 8823
rect 21324 8792 21465 8820
rect 21324 8780 21330 8792
rect 21453 8789 21465 8792
rect 21499 8789 21511 8823
rect 21744 8820 21772 8996
rect 21818 8916 21824 8968
rect 21876 8956 21882 8968
rect 21913 8959 21971 8965
rect 21913 8956 21925 8959
rect 21876 8928 21925 8956
rect 21876 8916 21882 8928
rect 21913 8925 21925 8928
rect 21959 8925 21971 8959
rect 21913 8919 21971 8925
rect 22066 8888 22094 8996
rect 24118 8916 24124 8968
rect 24176 8916 24182 8968
rect 22373 8891 22431 8897
rect 22373 8888 22385 8891
rect 22066 8860 22385 8888
rect 22373 8857 22385 8860
rect 22419 8888 22431 8891
rect 23109 8891 23167 8897
rect 23109 8888 23121 8891
rect 22419 8860 23121 8888
rect 22419 8857 22431 8860
rect 22373 8851 22431 8857
rect 23109 8857 23121 8860
rect 23155 8857 23167 8891
rect 23325 8891 23383 8897
rect 23325 8888 23337 8891
rect 23109 8851 23167 8857
rect 23216 8860 23337 8888
rect 22583 8823 22641 8829
rect 22583 8820 22595 8823
rect 21744 8792 22595 8820
rect 21453 8783 21511 8789
rect 22583 8789 22595 8792
rect 22629 8820 22641 8823
rect 23216 8820 23244 8860
rect 23325 8857 23337 8860
rect 23371 8888 23383 8891
rect 24670 8888 24676 8900
rect 23371 8860 24676 8888
rect 23371 8857 23383 8860
rect 23325 8851 23383 8857
rect 24670 8848 24676 8860
rect 24728 8848 24734 8900
rect 22629 8792 23244 8820
rect 22629 8789 22641 8792
rect 22583 8783 22641 8789
rect 1104 8730 24840 8752
rect 1104 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 24214 8730
rect 24266 8678 24278 8730
rect 24330 8678 24342 8730
rect 24394 8678 24406 8730
rect 24458 8678 24470 8730
rect 24522 8678 24840 8730
rect 1104 8656 24840 8678
rect 2130 8576 2136 8628
rect 2188 8576 2194 8628
rect 2222 8576 2228 8628
rect 2280 8616 2286 8628
rect 2409 8619 2467 8625
rect 2409 8616 2421 8619
rect 2280 8588 2421 8616
rect 2280 8576 2286 8588
rect 2409 8585 2421 8588
rect 2455 8585 2467 8619
rect 2409 8579 2467 8585
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 2866 8616 2872 8628
rect 2823 8588 2872 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 2866 8576 2872 8588
rect 2924 8616 2930 8628
rect 3326 8616 3332 8628
rect 2924 8588 3332 8616
rect 2924 8576 2930 8588
rect 3326 8576 3332 8588
rect 3384 8576 3390 8628
rect 4706 8616 4712 8628
rect 3528 8588 4712 8616
rect 1578 8508 1584 8560
rect 1636 8548 1642 8560
rect 1765 8551 1823 8557
rect 1765 8548 1777 8551
rect 1636 8520 1777 8548
rect 1636 8508 1642 8520
rect 1765 8517 1777 8520
rect 1811 8517 1823 8551
rect 1765 8511 1823 8517
rect 1981 8551 2039 8557
rect 1981 8517 1993 8551
rect 2027 8548 2039 8551
rect 3528 8548 3556 8588
rect 4706 8576 4712 8588
rect 4764 8576 4770 8628
rect 6362 8616 6368 8628
rect 5736 8588 6368 8616
rect 2027 8520 3556 8548
rect 2027 8517 2039 8520
rect 1981 8511 2039 8517
rect 2148 8492 2176 8520
rect 3602 8508 3608 8560
rect 3660 8548 3666 8560
rect 5736 8557 5764 8588
rect 6362 8576 6368 8588
rect 6420 8576 6426 8628
rect 6638 8576 6644 8628
rect 6696 8616 6702 8628
rect 9214 8616 9220 8628
rect 6696 8588 9220 8616
rect 6696 8576 6702 8588
rect 5721 8551 5779 8557
rect 3660 8520 5672 8548
rect 3660 8508 3666 8520
rect 2130 8440 2136 8492
rect 2188 8440 2194 8492
rect 2774 8440 2780 8492
rect 2832 8480 2838 8492
rect 2869 8483 2927 8489
rect 2869 8480 2881 8483
rect 2832 8452 2881 8480
rect 2832 8440 2838 8452
rect 2869 8449 2881 8452
rect 2915 8449 2927 8483
rect 2869 8443 2927 8449
rect 3418 8440 3424 8492
rect 3476 8480 3482 8492
rect 3881 8483 3939 8489
rect 3881 8480 3893 8483
rect 3476 8452 3893 8480
rect 3476 8440 3482 8452
rect 3881 8449 3893 8452
rect 3927 8449 3939 8483
rect 5644 8480 5672 8520
rect 5721 8517 5733 8551
rect 5767 8517 5779 8551
rect 5921 8551 5979 8557
rect 5921 8548 5933 8551
rect 5721 8511 5779 8517
rect 5828 8520 5933 8548
rect 5828 8480 5856 8520
rect 5921 8517 5933 8520
rect 5967 8548 5979 8551
rect 6454 8548 6460 8560
rect 5967 8520 6460 8548
rect 5967 8517 5979 8520
rect 5921 8511 5979 8517
rect 6454 8508 6460 8520
rect 6512 8548 6518 8560
rect 7282 8548 7288 8560
rect 6512 8520 7288 8548
rect 6512 8508 6518 8520
rect 7024 8492 7052 8520
rect 7282 8508 7288 8520
rect 7340 8508 7346 8560
rect 5644 8452 5856 8480
rect 3881 8443 3939 8449
rect 6362 8440 6368 8492
rect 6420 8480 6426 8492
rect 6822 8480 6828 8492
rect 6420 8452 6828 8480
rect 6420 8440 6426 8452
rect 6822 8440 6828 8452
rect 6880 8440 6886 8492
rect 6914 8440 6920 8492
rect 6972 8440 6978 8492
rect 7006 8440 7012 8492
rect 7064 8440 7070 8492
rect 7484 8489 7512 8588
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9953 8619 10011 8625
rect 9953 8585 9965 8619
rect 9999 8616 10011 8619
rect 10870 8616 10876 8628
rect 9999 8588 10876 8616
rect 9999 8585 10011 8588
rect 9953 8579 10011 8585
rect 10870 8576 10876 8588
rect 10928 8576 10934 8628
rect 14366 8576 14372 8628
rect 14424 8576 14430 8628
rect 15194 8576 15200 8628
rect 15252 8576 15258 8628
rect 15838 8616 15844 8628
rect 15304 8588 15844 8616
rect 7742 8508 7748 8560
rect 7800 8508 7806 8560
rect 8754 8508 8760 8560
rect 8812 8508 8818 8560
rect 10226 8548 10232 8560
rect 9784 8520 10232 8548
rect 9784 8489 9812 8520
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 10318 8508 10324 8560
rect 10376 8548 10382 8560
rect 15304 8548 15332 8588
rect 15838 8576 15844 8588
rect 15896 8576 15902 8628
rect 18690 8576 18696 8628
rect 18748 8616 18754 8628
rect 18748 8588 18920 8616
rect 18748 8576 18754 8588
rect 10376 8520 10916 8548
rect 10376 8508 10382 8520
rect 7469 8483 7527 8489
rect 7469 8449 7481 8483
rect 7515 8449 7527 8483
rect 7469 8443 7527 8449
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 9953 8483 10011 8489
rect 9953 8449 9965 8483
rect 9999 8449 10011 8483
rect 9953 8443 10011 8449
rect 3053 8415 3111 8421
rect 3053 8381 3065 8415
rect 3099 8412 3111 8415
rect 3142 8412 3148 8424
rect 3099 8384 3148 8412
rect 3099 8381 3111 8384
rect 3053 8375 3111 8381
rect 3142 8372 3148 8384
rect 3200 8372 3206 8424
rect 6733 8415 6791 8421
rect 6733 8381 6745 8415
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 3605 8347 3663 8353
rect 3605 8313 3617 8347
rect 3651 8344 3663 8347
rect 3786 8344 3792 8356
rect 3651 8316 3792 8344
rect 3651 8313 3663 8316
rect 3605 8307 3663 8313
rect 3786 8304 3792 8316
rect 3844 8304 3850 8356
rect 6454 8304 6460 8356
rect 6512 8344 6518 8356
rect 6748 8344 6776 8375
rect 7190 8372 7196 8424
rect 7248 8372 7254 8424
rect 9217 8415 9275 8421
rect 9217 8412 9229 8415
rect 7576 8384 9229 8412
rect 6914 8344 6920 8356
rect 6512 8316 6920 8344
rect 6512 8304 6518 8316
rect 6914 8304 6920 8316
rect 6972 8344 6978 8356
rect 7576 8344 7604 8384
rect 9217 8381 9229 8384
rect 9263 8381 9275 8415
rect 9968 8412 9996 8443
rect 10410 8440 10416 8492
rect 10468 8440 10474 8492
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 10778 8440 10784 8492
rect 10836 8440 10842 8492
rect 10888 8489 10916 8520
rect 11808 8520 15332 8548
rect 15365 8551 15423 8557
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11701 8483 11759 8489
rect 11701 8480 11713 8483
rect 10919 8452 11713 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11701 8449 11713 8452
rect 11747 8449 11759 8483
rect 11701 8443 11759 8449
rect 11054 8412 11060 8424
rect 9968 8384 11060 8412
rect 9217 8375 9275 8381
rect 6972 8316 7604 8344
rect 9232 8344 9260 8375
rect 11054 8372 11060 8384
rect 11112 8372 11118 8424
rect 11808 8412 11836 8520
rect 15365 8517 15377 8551
rect 15411 8517 15423 8551
rect 15365 8511 15423 8517
rect 11882 8440 11888 8492
rect 11940 8440 11946 8492
rect 11974 8440 11980 8492
rect 12032 8480 12038 8492
rect 12069 8483 12127 8489
rect 12069 8480 12081 8483
rect 12032 8452 12081 8480
rect 12032 8440 12038 8452
rect 12069 8449 12081 8452
rect 12115 8449 12127 8483
rect 12069 8443 12127 8449
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12618 8480 12624 8492
rect 12391 8452 12624 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 12802 8440 12808 8492
rect 12860 8480 12866 8492
rect 12897 8483 12955 8489
rect 12897 8480 12909 8483
rect 12860 8452 12909 8480
rect 12860 8440 12866 8452
rect 12897 8449 12909 8452
rect 12943 8449 12955 8483
rect 12897 8443 12955 8449
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 14734 8480 14740 8492
rect 13872 8452 14740 8480
rect 13872 8440 13878 8452
rect 14734 8440 14740 8452
rect 14792 8440 14798 8492
rect 15102 8440 15108 8492
rect 15160 8480 15166 8492
rect 15380 8480 15408 8511
rect 15470 8508 15476 8560
rect 15528 8548 15534 8560
rect 15565 8551 15623 8557
rect 15565 8548 15577 8551
rect 15528 8520 15577 8548
rect 15528 8508 15534 8520
rect 15565 8517 15577 8520
rect 15611 8548 15623 8551
rect 16666 8548 16672 8560
rect 15611 8520 16672 8548
rect 15611 8517 15623 8520
rect 15565 8511 15623 8517
rect 16666 8508 16672 8520
rect 16724 8508 16730 8560
rect 17218 8508 17224 8560
rect 17276 8508 17282 8560
rect 18782 8548 18788 8560
rect 18446 8520 18788 8548
rect 18782 8508 18788 8520
rect 18840 8508 18846 8560
rect 18892 8548 18920 8588
rect 19334 8576 19340 8628
rect 19392 8576 19398 8628
rect 19702 8576 19708 8628
rect 19760 8576 19766 8628
rect 20070 8576 20076 8628
rect 20128 8616 20134 8628
rect 20349 8619 20407 8625
rect 20349 8616 20361 8619
rect 20128 8588 20361 8616
rect 20128 8576 20134 8588
rect 20349 8585 20361 8588
rect 20395 8585 20407 8619
rect 20349 8579 20407 8585
rect 20517 8619 20575 8625
rect 20517 8585 20529 8619
rect 20563 8616 20575 8619
rect 21203 8619 21261 8625
rect 21203 8616 21215 8619
rect 20563 8588 21215 8616
rect 20563 8585 20575 8588
rect 20517 8579 20575 8585
rect 21203 8585 21215 8588
rect 21249 8616 21261 8619
rect 21542 8616 21548 8628
rect 21249 8588 21548 8616
rect 21249 8585 21261 8588
rect 21203 8579 21261 8585
rect 21542 8576 21548 8588
rect 21600 8616 21606 8628
rect 24187 8619 24245 8625
rect 24187 8616 24199 8619
rect 21600 8588 24199 8616
rect 21600 8576 21606 8588
rect 24187 8585 24199 8588
rect 24233 8585 24245 8619
rect 24187 8579 24245 8585
rect 19797 8551 19855 8557
rect 19797 8548 19809 8551
rect 18892 8520 19809 8548
rect 19797 8517 19809 8520
rect 19843 8517 19855 8551
rect 19797 8511 19855 8517
rect 20717 8551 20775 8557
rect 20717 8517 20729 8551
rect 20763 8517 20775 8551
rect 20717 8511 20775 8517
rect 15746 8480 15752 8492
rect 15160 8452 15752 8480
rect 15160 8440 15166 8452
rect 15746 8440 15752 8452
rect 15804 8440 15810 8492
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8449 15899 8483
rect 20732 8480 20760 8511
rect 20990 8508 20996 8560
rect 21048 8548 21054 8560
rect 21726 8548 21732 8560
rect 21048 8520 21732 8548
rect 21048 8508 21054 8520
rect 21726 8508 21732 8520
rect 21784 8508 21790 8560
rect 22186 8548 22192 8560
rect 22020 8520 22192 8548
rect 21082 8480 21088 8492
rect 20732 8452 21088 8480
rect 15841 8443 15899 8449
rect 11164 8384 11836 8412
rect 12989 8415 13047 8421
rect 11164 8344 11192 8384
rect 12989 8381 13001 8415
rect 13035 8381 13047 8415
rect 12989 8375 13047 8381
rect 9232 8316 11192 8344
rect 11609 8347 11667 8353
rect 6972 8304 6978 8316
rect 11609 8313 11621 8347
rect 11655 8344 11667 8347
rect 11698 8344 11704 8356
rect 11655 8316 11704 8344
rect 11655 8313 11667 8316
rect 11609 8307 11667 8313
rect 11698 8304 11704 8316
rect 11756 8304 11762 8356
rect 13004 8344 13032 8375
rect 14090 8372 14096 8424
rect 14148 8372 14154 8424
rect 14642 8372 14648 8424
rect 14700 8412 14706 8424
rect 15856 8412 15884 8443
rect 21082 8440 21088 8452
rect 21140 8480 21146 8492
rect 21358 8480 21364 8492
rect 21140 8452 21364 8480
rect 21140 8440 21146 8452
rect 21358 8440 21364 8452
rect 21416 8440 21422 8492
rect 22020 8489 22048 8520
rect 22186 8508 22192 8520
rect 22244 8508 22250 8560
rect 24397 8551 24455 8557
rect 24397 8517 24409 8551
rect 24443 8548 24455 8551
rect 24670 8548 24676 8560
rect 24443 8520 24676 8548
rect 24443 8517 24455 8520
rect 24397 8511 24455 8517
rect 24670 8508 24676 8520
rect 24728 8508 24734 8560
rect 22005 8483 22063 8489
rect 22005 8449 22017 8483
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 14700 8384 15884 8412
rect 14700 8372 14706 8384
rect 16114 8372 16120 8424
rect 16172 8372 16178 8424
rect 16942 8372 16948 8424
rect 17000 8372 17006 8424
rect 19702 8372 19708 8424
rect 19760 8412 19766 8424
rect 19886 8412 19892 8424
rect 19760 8384 19892 8412
rect 19760 8372 19766 8384
rect 19886 8372 19892 8384
rect 19944 8372 19950 8424
rect 22278 8372 22284 8424
rect 22336 8372 22342 8424
rect 23400 8412 23428 8466
rect 23400 8384 24072 8412
rect 15841 8347 15899 8353
rect 15841 8344 15853 8347
rect 13004 8316 15853 8344
rect 15841 8313 15853 8316
rect 15887 8313 15899 8347
rect 15841 8307 15899 8313
rect 15930 8304 15936 8356
rect 15988 8304 15994 8356
rect 18782 8304 18788 8356
rect 18840 8344 18846 8356
rect 18969 8347 19027 8353
rect 18969 8344 18981 8347
rect 18840 8316 18981 8344
rect 18840 8304 18846 8316
rect 18969 8313 18981 8316
rect 19015 8313 19027 8347
rect 20990 8344 20996 8356
rect 18969 8307 19027 8313
rect 19306 8316 20996 8344
rect 1946 8236 1952 8288
rect 2004 8236 2010 8288
rect 5534 8236 5540 8288
rect 5592 8276 5598 8288
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 5592 8248 5917 8276
rect 5592 8236 5598 8248
rect 5905 8245 5917 8248
rect 5951 8245 5963 8279
rect 5905 8239 5963 8245
rect 6089 8279 6147 8285
rect 6089 8245 6101 8279
rect 6135 8276 6147 8279
rect 6546 8276 6552 8288
rect 6135 8248 6552 8276
rect 6135 8245 6147 8248
rect 6089 8239 6147 8245
rect 6546 8236 6552 8248
rect 6604 8236 6610 8288
rect 7282 8236 7288 8288
rect 7340 8276 7346 8288
rect 10042 8276 10048 8288
rect 7340 8248 10048 8276
rect 7340 8236 7346 8248
rect 10042 8236 10048 8248
rect 10100 8236 10106 8288
rect 13265 8279 13323 8285
rect 13265 8245 13277 8279
rect 13311 8276 13323 8279
rect 13446 8276 13452 8288
rect 13311 8248 13452 8276
rect 13311 8245 13323 8248
rect 13265 8239 13323 8245
rect 13446 8236 13452 8248
rect 13504 8236 13510 8288
rect 13538 8236 13544 8288
rect 13596 8276 13602 8288
rect 13633 8279 13691 8285
rect 13633 8276 13645 8279
rect 13596 8248 13645 8276
rect 13596 8236 13602 8248
rect 13633 8245 13645 8248
rect 13679 8245 13691 8279
rect 13633 8239 13691 8245
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 15381 8279 15439 8285
rect 15381 8276 15393 8279
rect 15068 8248 15393 8276
rect 15068 8236 15074 8248
rect 15381 8245 15393 8248
rect 15427 8276 15439 8279
rect 16574 8276 16580 8288
rect 15427 8248 16580 8276
rect 15427 8245 15439 8248
rect 15381 8239 15439 8245
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 18874 8236 18880 8288
rect 18932 8276 18938 8288
rect 19306 8276 19334 8316
rect 20990 8304 20996 8316
rect 21048 8304 21054 8356
rect 21358 8304 21364 8356
rect 21416 8304 21422 8356
rect 23290 8304 23296 8356
rect 23348 8344 23354 8356
rect 24044 8353 24072 8384
rect 23753 8347 23811 8353
rect 23753 8344 23765 8347
rect 23348 8316 23765 8344
rect 23348 8304 23354 8316
rect 23753 8313 23765 8316
rect 23799 8313 23811 8347
rect 23753 8307 23811 8313
rect 24029 8347 24087 8353
rect 24029 8313 24041 8347
rect 24075 8313 24087 8347
rect 24029 8307 24087 8313
rect 18932 8248 19334 8276
rect 20533 8279 20591 8285
rect 18932 8236 18938 8248
rect 20533 8245 20545 8279
rect 20579 8276 20591 8279
rect 21174 8276 21180 8288
rect 20579 8248 21180 8276
rect 20579 8245 20591 8248
rect 20533 8239 20591 8245
rect 21174 8236 21180 8248
rect 21232 8236 21238 8288
rect 21634 8236 21640 8288
rect 21692 8276 21698 8288
rect 23658 8276 23664 8288
rect 21692 8248 23664 8276
rect 21692 8236 21698 8248
rect 23658 8236 23664 8248
rect 23716 8236 23722 8288
rect 23842 8236 23848 8288
rect 23900 8276 23906 8288
rect 24213 8279 24271 8285
rect 24213 8276 24225 8279
rect 23900 8248 24225 8276
rect 23900 8236 23906 8248
rect 24213 8245 24225 8248
rect 24259 8245 24271 8279
rect 24213 8239 24271 8245
rect 1104 8186 24840 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 20214 8186
rect 20266 8134 20278 8186
rect 20330 8134 20342 8186
rect 20394 8134 20406 8186
rect 20458 8134 20470 8186
rect 20522 8134 24840 8186
rect 1104 8112 24840 8134
rect 1670 8032 1676 8084
rect 1728 8032 1734 8084
rect 3142 8032 3148 8084
rect 3200 8072 3206 8084
rect 6270 8072 6276 8084
rect 3200 8044 6276 8072
rect 3200 8032 3206 8044
rect 6270 8032 6276 8044
rect 6328 8072 6334 8084
rect 6733 8075 6791 8081
rect 6328 8044 6684 8072
rect 6328 8032 6334 8044
rect 6656 8004 6684 8044
rect 6733 8041 6745 8075
rect 6779 8072 6791 8075
rect 7098 8072 7104 8084
rect 6779 8044 7104 8072
rect 6779 8041 6791 8044
rect 6733 8035 6791 8041
rect 7098 8032 7104 8044
rect 7156 8032 7162 8084
rect 7190 8032 7196 8084
rect 7248 8072 7254 8084
rect 7466 8072 7472 8084
rect 7248 8044 7472 8072
rect 7248 8032 7254 8044
rect 7466 8032 7472 8044
rect 7524 8032 7530 8084
rect 7558 8032 7564 8084
rect 7616 8032 7622 8084
rect 10502 8032 10508 8084
rect 10560 8072 10566 8084
rect 10597 8075 10655 8081
rect 10597 8072 10609 8075
rect 10560 8044 10609 8072
rect 10560 8032 10566 8044
rect 10597 8041 10609 8044
rect 10643 8041 10655 8075
rect 10597 8035 10655 8041
rect 11054 8032 11060 8084
rect 11112 8072 11118 8084
rect 11974 8072 11980 8084
rect 11112 8044 11980 8072
rect 11112 8032 11118 8044
rect 11974 8032 11980 8044
rect 12032 8032 12038 8084
rect 12894 8032 12900 8084
rect 12952 8072 12958 8084
rect 12989 8075 13047 8081
rect 12989 8072 13001 8075
rect 12952 8044 13001 8072
rect 12952 8032 12958 8044
rect 12989 8041 13001 8044
rect 13035 8041 13047 8075
rect 12989 8035 13047 8041
rect 13817 8075 13875 8081
rect 13817 8041 13829 8075
rect 13863 8072 13875 8075
rect 15930 8072 15936 8084
rect 13863 8044 15936 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 15930 8032 15936 8044
rect 15988 8032 15994 8084
rect 16574 8032 16580 8084
rect 16632 8072 16638 8084
rect 17129 8075 17187 8081
rect 17129 8072 17141 8075
rect 16632 8044 17141 8072
rect 16632 8032 16638 8044
rect 17129 8041 17141 8044
rect 17175 8072 17187 8075
rect 17678 8072 17684 8084
rect 17175 8044 17684 8072
rect 17175 8041 17187 8044
rect 17129 8035 17187 8041
rect 17678 8032 17684 8044
rect 17736 8072 17742 8084
rect 18785 8075 18843 8081
rect 18785 8072 18797 8075
rect 17736 8044 18797 8072
rect 17736 8032 17742 8044
rect 18785 8041 18797 8044
rect 18831 8072 18843 8075
rect 18966 8072 18972 8084
rect 18831 8044 18972 8072
rect 18831 8041 18843 8044
rect 18785 8035 18843 8041
rect 18966 8032 18972 8044
rect 19024 8032 19030 8084
rect 19518 8032 19524 8084
rect 19576 8072 19582 8084
rect 19576 8044 21128 8072
rect 19576 8032 19582 8044
rect 7282 8004 7288 8016
rect 6656 7976 7288 8004
rect 2866 7896 2872 7948
rect 2924 7896 2930 7948
rect 3053 7939 3111 7945
rect 3053 7905 3065 7939
rect 3099 7936 3111 7939
rect 3142 7936 3148 7948
rect 3099 7908 3148 7936
rect 3099 7905 3111 7908
rect 3053 7899 3111 7905
rect 3142 7896 3148 7908
rect 3200 7896 3206 7948
rect 3602 7896 3608 7948
rect 3660 7936 3666 7948
rect 3881 7939 3939 7945
rect 3881 7936 3893 7939
rect 3660 7908 3893 7936
rect 3660 7896 3666 7908
rect 3881 7905 3893 7908
rect 3927 7936 3939 7939
rect 4062 7936 4068 7948
rect 3927 7908 4068 7936
rect 3927 7905 3939 7908
rect 3881 7899 3939 7905
rect 4062 7896 4068 7908
rect 4120 7896 4126 7948
rect 5905 7939 5963 7945
rect 5905 7905 5917 7939
rect 5951 7936 5963 7939
rect 6638 7936 6644 7948
rect 5951 7908 6644 7936
rect 5951 7905 5963 7908
rect 5905 7899 5963 7905
rect 6638 7896 6644 7908
rect 6696 7896 6702 7948
rect 1394 7828 1400 7880
rect 1452 7868 1458 7880
rect 1489 7871 1547 7877
rect 1489 7868 1501 7871
rect 1452 7840 1501 7868
rect 1452 7828 1458 7840
rect 1489 7837 1501 7840
rect 1535 7837 1547 7871
rect 1489 7831 1547 7837
rect 1504 7800 1532 7831
rect 1670 7828 1676 7880
rect 1728 7868 1734 7880
rect 2133 7871 2191 7877
rect 2133 7868 2145 7871
rect 1728 7840 2145 7868
rect 1728 7828 1734 7840
rect 2133 7837 2145 7840
rect 2179 7868 2191 7871
rect 2682 7868 2688 7880
rect 2179 7840 2688 7868
rect 2179 7837 2191 7840
rect 2133 7831 2191 7837
rect 2682 7828 2688 7840
rect 2740 7828 2746 7880
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7868 6515 7871
rect 6546 7868 6552 7880
rect 6503 7840 6552 7868
rect 6503 7837 6515 7840
rect 6457 7831 6515 7837
rect 6546 7828 6552 7840
rect 6604 7828 6610 7880
rect 6736 7871 6794 7877
rect 6736 7837 6748 7871
rect 6782 7868 6794 7871
rect 6840 7868 6868 7976
rect 7282 7964 7288 7976
rect 7340 7964 7346 8016
rect 7576 8004 7604 8032
rect 7484 7976 7604 8004
rect 7484 7945 7512 7976
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 11146 8004 11152 8016
rect 7800 7976 11152 8004
rect 7800 7964 7806 7976
rect 11146 7964 11152 7976
rect 11204 7964 11210 8016
rect 12253 8007 12311 8013
rect 11256 7976 12204 8004
rect 7469 7939 7527 7945
rect 7469 7905 7481 7939
rect 7515 7905 7527 7939
rect 7469 7899 7527 7905
rect 7926 7896 7932 7948
rect 7984 7936 7990 7948
rect 10137 7939 10195 7945
rect 7984 7908 9352 7936
rect 7984 7896 7990 7908
rect 6782 7840 6868 7868
rect 6782 7837 6794 7840
rect 6736 7831 6794 7837
rect 7098 7828 7104 7880
rect 7156 7868 7162 7880
rect 7193 7871 7251 7877
rect 7193 7868 7205 7871
rect 7156 7840 7205 7868
rect 7156 7828 7162 7840
rect 7193 7837 7205 7840
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 7285 7871 7343 7877
rect 7285 7837 7297 7871
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7865 7435 7871
rect 7834 7868 7840 7880
rect 7576 7865 7840 7868
rect 7423 7840 7840 7865
rect 7423 7837 7604 7840
rect 7377 7831 7435 7837
rect 3421 7803 3479 7809
rect 3421 7800 3433 7803
rect 1504 7772 3433 7800
rect 3421 7769 3433 7772
rect 3467 7769 3479 7803
rect 3421 7763 3479 7769
rect 4614 7760 4620 7812
rect 4672 7760 4678 7812
rect 5629 7803 5687 7809
rect 5629 7769 5641 7803
rect 5675 7800 5687 7803
rect 5675 7772 6684 7800
rect 5675 7769 5687 7772
rect 5629 7763 5687 7769
rect 1762 7692 1768 7744
rect 1820 7732 1826 7744
rect 2041 7735 2099 7741
rect 2041 7732 2053 7735
rect 1820 7704 2053 7732
rect 1820 7692 1826 7704
rect 2041 7701 2053 7704
rect 2087 7701 2099 7735
rect 2041 7695 2099 7701
rect 2406 7692 2412 7744
rect 2464 7692 2470 7744
rect 2777 7735 2835 7741
rect 2777 7701 2789 7735
rect 2823 7732 2835 7735
rect 3234 7732 3240 7744
rect 2823 7704 3240 7732
rect 2823 7701 2835 7704
rect 2777 7695 2835 7701
rect 3234 7692 3240 7704
rect 3292 7692 3298 7744
rect 6454 7692 6460 7744
rect 6512 7732 6518 7744
rect 6549 7735 6607 7741
rect 6549 7732 6561 7735
rect 6512 7704 6561 7732
rect 6512 7692 6518 7704
rect 6549 7701 6561 7704
rect 6595 7701 6607 7735
rect 6656 7732 6684 7772
rect 7009 7735 7067 7741
rect 7009 7732 7021 7735
rect 6656 7704 7021 7732
rect 6549 7695 6607 7701
rect 7009 7701 7021 7704
rect 7055 7701 7067 7735
rect 7300 7732 7328 7831
rect 7834 7828 7840 7840
rect 7892 7868 7898 7880
rect 8110 7868 8116 7880
rect 7892 7840 8116 7868
rect 7892 7828 7898 7840
rect 8110 7828 8116 7840
rect 8168 7868 8174 7880
rect 8404 7877 8432 7908
rect 8297 7871 8355 7877
rect 8297 7868 8309 7871
rect 8168 7840 8309 7868
rect 8168 7828 8174 7840
rect 8297 7837 8309 7840
rect 8343 7837 8355 7871
rect 8297 7831 8355 7837
rect 8389 7871 8447 7877
rect 8389 7837 8401 7871
rect 8435 7837 8447 7871
rect 8389 7831 8447 7837
rect 8481 7871 8539 7877
rect 8481 7837 8493 7871
rect 8527 7837 8539 7871
rect 8481 7831 8539 7837
rect 7650 7732 7656 7744
rect 7300 7704 7656 7732
rect 7009 7695 7067 7701
rect 7650 7692 7656 7704
rect 7708 7732 7714 7744
rect 8496 7732 8524 7831
rect 9030 7828 9036 7880
rect 9088 7828 9094 7880
rect 9324 7877 9352 7908
rect 10137 7905 10149 7939
rect 10183 7936 10195 7939
rect 10505 7939 10563 7945
rect 10505 7936 10517 7939
rect 10183 7908 10517 7936
rect 10183 7905 10195 7908
rect 10137 7899 10195 7905
rect 10505 7905 10517 7908
rect 10551 7905 10563 7939
rect 11256 7936 11284 7976
rect 10505 7899 10563 7905
rect 10704 7908 11284 7936
rect 9217 7871 9275 7877
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9309 7871 9367 7877
rect 9309 7837 9321 7871
rect 9355 7837 9367 7871
rect 9309 7831 9367 7837
rect 9401 7871 9459 7877
rect 9401 7837 9413 7871
rect 9447 7868 9459 7871
rect 9582 7868 9588 7880
rect 9447 7840 9588 7868
rect 9447 7837 9459 7840
rect 9401 7831 9459 7837
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 9232 7800 9260 7831
rect 8711 7772 9260 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 9416 7732 9444 7831
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 10045 7871 10103 7877
rect 10045 7837 10057 7871
rect 10091 7837 10103 7871
rect 10045 7831 10103 7837
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7868 10287 7871
rect 10704 7868 10732 7908
rect 11330 7896 11336 7948
rect 11388 7896 11394 7948
rect 12176 7936 12204 7976
rect 12253 7973 12265 8007
rect 12299 8004 12311 8007
rect 13722 8004 13728 8016
rect 12299 7976 13728 8004
rect 12299 7973 12311 7976
rect 12253 7967 12311 7973
rect 13722 7964 13728 7976
rect 13780 7964 13786 8016
rect 19610 8004 19616 8016
rect 16776 7976 19616 8004
rect 12802 7936 12808 7948
rect 12176 7908 12808 7936
rect 12802 7896 12808 7908
rect 12860 7936 12866 7948
rect 12860 7908 13124 7936
rect 12860 7896 12866 7908
rect 10275 7840 10732 7868
rect 10781 7871 10839 7877
rect 10275 7837 10287 7840
rect 10229 7831 10287 7837
rect 10781 7837 10793 7871
rect 10827 7837 10839 7871
rect 10781 7831 10839 7837
rect 10060 7800 10088 7831
rect 10686 7800 10692 7812
rect 10060 7772 10692 7800
rect 10686 7760 10692 7772
rect 10744 7760 10750 7812
rect 7708 7704 9444 7732
rect 7708 7692 7714 7704
rect 9490 7692 9496 7744
rect 9548 7732 9554 7744
rect 9677 7735 9735 7741
rect 9677 7732 9689 7735
rect 9548 7704 9689 7732
rect 9548 7692 9554 7704
rect 9677 7701 9689 7704
rect 9723 7701 9735 7735
rect 10796 7732 10824 7831
rect 11054 7828 11060 7880
rect 11112 7828 11118 7880
rect 11348 7868 11376 7896
rect 11609 7871 11667 7877
rect 11609 7868 11621 7871
rect 11348 7840 11621 7868
rect 11609 7837 11621 7840
rect 11655 7837 11667 7871
rect 11609 7831 11667 7837
rect 11698 7828 11704 7880
rect 11756 7868 11762 7880
rect 11793 7871 11851 7877
rect 11793 7868 11805 7871
rect 11756 7840 11805 7868
rect 11756 7828 11762 7840
rect 11793 7837 11805 7840
rect 11839 7837 11851 7871
rect 11793 7831 11851 7837
rect 11882 7828 11888 7880
rect 11940 7828 11946 7880
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7868 12035 7871
rect 12618 7868 12624 7880
rect 12023 7840 12624 7868
rect 12023 7837 12035 7840
rect 11977 7831 12035 7837
rect 11333 7803 11391 7809
rect 11333 7769 11345 7803
rect 11379 7800 11391 7803
rect 11992 7800 12020 7831
rect 12618 7828 12624 7840
rect 12676 7828 12682 7880
rect 11379 7772 12020 7800
rect 13096 7800 13124 7908
rect 13188 7908 13400 7936
rect 13188 7880 13216 7908
rect 13170 7828 13176 7880
rect 13228 7828 13234 7880
rect 13265 7871 13323 7877
rect 13265 7837 13277 7871
rect 13311 7837 13323 7871
rect 13372 7868 13400 7908
rect 13446 7896 13452 7948
rect 13504 7936 13510 7948
rect 14461 7939 14519 7945
rect 14461 7936 14473 7939
rect 13504 7908 14473 7936
rect 13504 7896 13510 7908
rect 14461 7905 14473 7908
rect 14507 7905 14519 7939
rect 14461 7899 14519 7905
rect 14918 7896 14924 7948
rect 14976 7936 14982 7948
rect 15470 7936 15476 7948
rect 14976 7908 15476 7936
rect 14976 7896 14982 7908
rect 15470 7896 15476 7908
rect 15528 7896 15534 7948
rect 13633 7871 13691 7877
rect 13633 7868 13645 7871
rect 13372 7840 13645 7868
rect 13265 7831 13323 7837
rect 13633 7837 13645 7840
rect 13679 7868 13691 7871
rect 13722 7868 13728 7880
rect 13679 7840 13728 7868
rect 13679 7837 13691 7840
rect 13633 7831 13691 7837
rect 13280 7800 13308 7831
rect 13722 7828 13728 7840
rect 13780 7828 13786 7880
rect 13817 7871 13875 7877
rect 13817 7837 13829 7871
rect 13863 7868 13875 7871
rect 14090 7868 14096 7880
rect 13863 7840 14096 7868
rect 13863 7837 13875 7840
rect 13817 7831 13875 7837
rect 14090 7828 14096 7840
rect 14148 7828 14154 7880
rect 14182 7828 14188 7880
rect 14240 7828 14246 7880
rect 16776 7877 16804 7976
rect 19610 7964 19616 7976
rect 19668 7964 19674 8016
rect 21100 8004 21128 8044
rect 21174 8032 21180 8084
rect 21232 8072 21238 8084
rect 21232 8044 22094 8072
rect 21232 8032 21238 8044
rect 21910 8004 21916 8016
rect 21100 7976 21916 8004
rect 21910 7964 21916 7976
rect 21968 7964 21974 8016
rect 22066 8004 22094 8044
rect 22278 8032 22284 8084
rect 22336 8072 22342 8084
rect 22925 8075 22983 8081
rect 22925 8072 22937 8075
rect 22336 8044 22937 8072
rect 22336 8032 22342 8044
rect 22925 8041 22937 8044
rect 22971 8041 22983 8075
rect 22925 8035 22983 8041
rect 23842 8004 23848 8016
rect 22066 7976 23848 8004
rect 23842 7964 23848 7976
rect 23900 7964 23906 8016
rect 17494 7896 17500 7948
rect 17552 7936 17558 7948
rect 18230 7936 18236 7948
rect 17552 7908 18236 7936
rect 17552 7896 17558 7908
rect 18230 7896 18236 7908
rect 18288 7896 18294 7948
rect 18690 7896 18696 7948
rect 18748 7936 18754 7948
rect 18748 7908 19656 7936
rect 18748 7896 18754 7908
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7837 16819 7871
rect 16761 7831 16819 7837
rect 17313 7871 17371 7877
rect 17313 7837 17325 7871
rect 17359 7868 17371 7871
rect 17586 7868 17592 7880
rect 17359 7840 17592 7868
rect 17359 7837 17371 7840
rect 17313 7831 17371 7837
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7868 18015 7871
rect 19628 7868 19656 7908
rect 19702 7896 19708 7948
rect 19760 7936 19766 7948
rect 19889 7939 19947 7945
rect 19889 7936 19901 7939
rect 19760 7908 19901 7936
rect 19760 7896 19766 7908
rect 19889 7905 19901 7908
rect 19935 7936 19947 7939
rect 21085 7939 21143 7945
rect 21085 7936 21097 7939
rect 19935 7908 21097 7936
rect 19935 7905 19947 7908
rect 19889 7899 19947 7905
rect 21085 7905 21097 7908
rect 21131 7936 21143 7939
rect 22005 7939 22063 7945
rect 22005 7936 22017 7939
rect 21131 7908 22017 7936
rect 21131 7905 21143 7908
rect 21085 7899 21143 7905
rect 22005 7905 22017 7908
rect 22051 7905 22063 7939
rect 22005 7899 22063 7905
rect 22094 7896 22100 7948
rect 22152 7936 22158 7948
rect 22646 7936 22652 7948
rect 22152 7908 22652 7936
rect 22152 7896 22158 7908
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 23382 7896 23388 7948
rect 23440 7896 23446 7948
rect 23477 7939 23535 7945
rect 23477 7905 23489 7939
rect 23523 7905 23535 7939
rect 23477 7899 23535 7905
rect 22112 7868 22140 7896
rect 18003 7840 19564 7868
rect 19628 7840 22140 7868
rect 22189 7871 22247 7877
rect 18003 7837 18015 7840
rect 17957 7831 18015 7837
rect 13096 7772 13308 7800
rect 11379 7769 11391 7772
rect 11333 7763 11391 7769
rect 11698 7732 11704 7744
rect 10796 7704 11704 7732
rect 9677 7695 9735 7701
rect 11698 7692 11704 7704
rect 11756 7692 11762 7744
rect 13280 7732 13308 7772
rect 14734 7760 14740 7812
rect 14792 7800 14798 7812
rect 14792 7772 14950 7800
rect 14792 7760 14798 7772
rect 15746 7760 15752 7812
rect 15804 7800 15810 7812
rect 18690 7800 18696 7812
rect 15804 7772 16620 7800
rect 15804 7760 15810 7772
rect 15838 7732 15844 7744
rect 13280 7704 15844 7732
rect 15838 7692 15844 7704
rect 15896 7732 15902 7744
rect 16592 7741 16620 7772
rect 17144 7772 18696 7800
rect 17144 7744 17172 7772
rect 18690 7760 18696 7772
rect 18748 7809 18754 7812
rect 18748 7803 18811 7809
rect 18748 7769 18765 7803
rect 18799 7769 18811 7803
rect 18748 7763 18811 7769
rect 18748 7760 18754 7763
rect 18874 7760 18880 7812
rect 18932 7800 18938 7812
rect 18969 7803 19027 7809
rect 18969 7800 18981 7803
rect 18932 7772 18981 7800
rect 18932 7760 18938 7772
rect 18969 7769 18981 7772
rect 19015 7769 19027 7803
rect 18969 7763 19027 7769
rect 15933 7735 15991 7741
rect 15933 7732 15945 7735
rect 15896 7704 15945 7732
rect 15896 7692 15902 7704
rect 15933 7701 15945 7704
rect 15979 7701 15991 7735
rect 15933 7695 15991 7701
rect 16577 7735 16635 7741
rect 16577 7701 16589 7735
rect 16623 7732 16635 7735
rect 17126 7732 17132 7744
rect 16623 7704 17132 7732
rect 16623 7701 16635 7704
rect 16577 7695 16635 7701
rect 17126 7692 17132 7704
rect 17184 7692 17190 7744
rect 17402 7692 17408 7744
rect 17460 7732 17466 7744
rect 17589 7735 17647 7741
rect 17589 7732 17601 7735
rect 17460 7704 17601 7732
rect 17460 7692 17466 7704
rect 17589 7701 17601 7704
rect 17635 7701 17647 7735
rect 17589 7695 17647 7701
rect 18046 7692 18052 7744
rect 18104 7692 18110 7744
rect 18506 7692 18512 7744
rect 18564 7732 18570 7744
rect 18601 7735 18659 7741
rect 18601 7732 18613 7735
rect 18564 7704 18613 7732
rect 18564 7692 18570 7704
rect 18601 7701 18613 7704
rect 18647 7701 18659 7735
rect 18601 7695 18659 7701
rect 19337 7735 19395 7741
rect 19337 7701 19349 7735
rect 19383 7732 19395 7735
rect 19426 7732 19432 7744
rect 19383 7704 19432 7732
rect 19383 7701 19395 7704
rect 19337 7695 19395 7701
rect 19426 7692 19432 7704
rect 19484 7692 19490 7744
rect 19536 7732 19564 7840
rect 22189 7837 22201 7871
rect 22235 7868 22247 7871
rect 23290 7868 23296 7880
rect 22235 7840 23296 7868
rect 22235 7837 22247 7840
rect 22189 7831 22247 7837
rect 23290 7828 23296 7840
rect 23348 7828 23354 7880
rect 23492 7868 23520 7899
rect 23400 7840 23520 7868
rect 19705 7803 19763 7809
rect 19705 7769 19717 7803
rect 19751 7800 19763 7803
rect 20806 7800 20812 7812
rect 19751 7772 20812 7800
rect 19751 7769 19763 7772
rect 19705 7763 19763 7769
rect 20806 7760 20812 7772
rect 20864 7800 20870 7812
rect 20993 7803 21051 7809
rect 20993 7800 21005 7803
rect 20864 7772 21005 7800
rect 20864 7760 20870 7772
rect 20993 7769 21005 7772
rect 21039 7769 21051 7803
rect 20993 7763 21051 7769
rect 22094 7760 22100 7812
rect 22152 7800 22158 7812
rect 22281 7803 22339 7809
rect 22281 7800 22293 7803
rect 22152 7772 22293 7800
rect 22152 7760 22158 7772
rect 22281 7769 22293 7772
rect 22327 7800 22339 7803
rect 22922 7800 22928 7812
rect 22327 7772 22928 7800
rect 22327 7769 22339 7772
rect 22281 7763 22339 7769
rect 22922 7760 22928 7772
rect 22980 7760 22986 7812
rect 23014 7760 23020 7812
rect 23072 7800 23078 7812
rect 23400 7800 23428 7840
rect 23658 7828 23664 7880
rect 23716 7868 23722 7880
rect 24118 7868 24124 7880
rect 23716 7840 24124 7868
rect 23716 7828 23722 7840
rect 24118 7828 24124 7840
rect 24176 7828 24182 7880
rect 23072 7772 23428 7800
rect 23072 7760 23078 7772
rect 19794 7732 19800 7744
rect 19536 7704 19800 7732
rect 19794 7692 19800 7704
rect 19852 7692 19858 7744
rect 20070 7692 20076 7744
rect 20128 7732 20134 7744
rect 20533 7735 20591 7741
rect 20533 7732 20545 7735
rect 20128 7704 20545 7732
rect 20128 7692 20134 7704
rect 20533 7701 20545 7704
rect 20579 7701 20591 7735
rect 20533 7695 20591 7701
rect 20898 7692 20904 7744
rect 20956 7692 20962 7744
rect 21637 7735 21695 7741
rect 21637 7701 21649 7735
rect 21683 7732 21695 7735
rect 21818 7732 21824 7744
rect 21683 7704 21824 7732
rect 21683 7701 21695 7704
rect 21637 7695 21695 7701
rect 21818 7692 21824 7704
rect 21876 7692 21882 7744
rect 22554 7692 22560 7744
rect 22612 7732 22618 7744
rect 22649 7735 22707 7741
rect 22649 7732 22661 7735
rect 22612 7704 22661 7732
rect 22612 7692 22618 7704
rect 22649 7701 22661 7704
rect 22695 7701 22707 7735
rect 22649 7695 22707 7701
rect 22738 7692 22744 7744
rect 22796 7732 22802 7744
rect 23937 7735 23995 7741
rect 23937 7732 23949 7735
rect 22796 7704 23949 7732
rect 22796 7692 22802 7704
rect 23937 7701 23949 7704
rect 23983 7701 23995 7735
rect 23937 7695 23995 7701
rect 1104 7642 24840 7664
rect 1104 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 24214 7642
rect 24266 7590 24278 7642
rect 24330 7590 24342 7642
rect 24394 7590 24406 7642
rect 24458 7590 24470 7642
rect 24522 7590 24840 7642
rect 1104 7568 24840 7590
rect 2406 7528 2412 7540
rect 1780 7500 2412 7528
rect 1780 7469 1808 7500
rect 2406 7488 2412 7500
rect 2464 7488 2470 7540
rect 3234 7488 3240 7540
rect 3292 7528 3298 7540
rect 4525 7531 4583 7537
rect 3292 7500 4476 7528
rect 3292 7488 3298 7500
rect 1765 7463 1823 7469
rect 1765 7429 1777 7463
rect 1811 7429 1823 7463
rect 1765 7423 1823 7429
rect 4157 7463 4215 7469
rect 4157 7429 4169 7463
rect 4203 7429 4215 7463
rect 4357 7463 4415 7469
rect 4357 7460 4369 7463
rect 4157 7423 4215 7429
rect 4356 7429 4369 7460
rect 4403 7429 4415 7463
rect 4448 7460 4476 7500
rect 4525 7497 4537 7531
rect 4571 7528 4583 7531
rect 4614 7528 4620 7540
rect 4571 7500 4620 7528
rect 4571 7497 4583 7500
rect 4525 7491 4583 7497
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 7282 7488 7288 7540
rect 7340 7488 7346 7540
rect 7926 7488 7932 7540
rect 7984 7488 7990 7540
rect 8110 7488 8116 7540
rect 8168 7528 8174 7540
rect 12710 7528 12716 7540
rect 8168 7500 12716 7528
rect 8168 7488 8174 7500
rect 12710 7488 12716 7500
rect 12768 7488 12774 7540
rect 12986 7537 12992 7540
rect 12805 7531 12863 7537
rect 12805 7497 12817 7531
rect 12851 7497 12863 7531
rect 12805 7491 12863 7497
rect 12973 7531 12992 7537
rect 12973 7497 12985 7531
rect 13044 7528 13050 7540
rect 14645 7531 14703 7537
rect 13044 7500 14596 7528
rect 12973 7491 12992 7497
rect 5810 7460 5816 7472
rect 4448 7432 5816 7460
rect 4356 7423 4415 7429
rect 2866 7352 2872 7404
rect 2924 7352 2930 7404
rect 3786 7392 3792 7404
rect 3747 7364 3792 7392
rect 3786 7352 3792 7364
rect 3844 7352 3850 7404
rect 3881 7395 3939 7401
rect 3881 7361 3893 7395
rect 3927 7392 3939 7395
rect 3970 7392 3976 7404
rect 3927 7364 3976 7392
rect 3927 7361 3939 7364
rect 3881 7355 3939 7361
rect 3970 7352 3976 7364
rect 4028 7352 4034 7404
rect 1486 7284 1492 7336
rect 1544 7284 1550 7336
rect 2498 7284 2504 7336
rect 2556 7324 2562 7336
rect 4172 7324 4200 7423
rect 4356 7392 4384 7423
rect 5810 7420 5816 7432
rect 5868 7420 5874 7472
rect 6457 7463 6515 7469
rect 6457 7460 6469 7463
rect 5920 7432 6469 7460
rect 5920 7404 5948 7432
rect 6457 7429 6469 7432
rect 6503 7429 6515 7463
rect 6457 7423 6515 7429
rect 6546 7420 6552 7472
rect 6604 7460 6610 7472
rect 7453 7463 7511 7469
rect 7453 7460 7465 7463
rect 6604 7432 7465 7460
rect 6604 7420 6610 7432
rect 7453 7429 7465 7432
rect 7499 7460 7511 7463
rect 7499 7429 7512 7460
rect 7453 7423 7512 7429
rect 4706 7392 4712 7404
rect 4356 7364 4712 7392
rect 4706 7352 4712 7364
rect 4764 7392 4770 7404
rect 5074 7392 5080 7404
rect 4764 7364 5080 7392
rect 4764 7352 4770 7364
rect 5074 7352 5080 7364
rect 5132 7352 5138 7404
rect 5166 7352 5172 7404
rect 5224 7352 5230 7404
rect 5902 7352 5908 7404
rect 5960 7352 5966 7404
rect 6086 7352 6092 7404
rect 6144 7352 6150 7404
rect 6638 7352 6644 7404
rect 6696 7352 6702 7404
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7392 6791 7395
rect 6822 7392 6828 7404
rect 6779 7364 6828 7392
rect 6779 7361 6791 7364
rect 6733 7355 6791 7361
rect 2556 7296 4200 7324
rect 2556 7284 2562 7296
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 6748 7324 6776 7355
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 7484 7392 7512 7423
rect 7650 7420 7656 7472
rect 7708 7420 7714 7472
rect 8662 7460 8668 7472
rect 8220 7432 8668 7460
rect 8113 7395 8171 7401
rect 8113 7392 8125 7395
rect 7484 7364 8125 7392
rect 8113 7361 8125 7364
rect 8159 7361 8171 7395
rect 8113 7355 8171 7361
rect 5684 7296 6776 7324
rect 5684 7284 5690 7296
rect 3142 7216 3148 7268
rect 3200 7256 3206 7268
rect 3513 7259 3571 7265
rect 3513 7256 3525 7259
rect 3200 7228 3525 7256
rect 3200 7216 3206 7228
rect 3513 7225 3525 7228
rect 3559 7225 3571 7259
rect 4798 7256 4804 7268
rect 3513 7219 3571 7225
rect 4356 7228 4804 7256
rect 1946 7148 1952 7200
rect 2004 7188 2010 7200
rect 4356 7197 4384 7228
rect 4798 7216 4804 7228
rect 4856 7256 4862 7268
rect 6362 7256 6368 7268
rect 4856 7228 6368 7256
rect 4856 7216 4862 7228
rect 6362 7216 6368 7228
rect 6420 7256 6426 7268
rect 8220 7256 8248 7432
rect 8662 7420 8668 7432
rect 8720 7460 8726 7472
rect 8720 7432 8984 7460
rect 8720 7420 8726 7432
rect 8573 7395 8631 7401
rect 8573 7361 8585 7395
rect 8619 7392 8631 7395
rect 8754 7392 8760 7404
rect 8619 7364 8760 7392
rect 8619 7361 8631 7364
rect 8573 7355 8631 7361
rect 8754 7352 8760 7364
rect 8812 7352 8818 7404
rect 8297 7327 8355 7333
rect 8297 7293 8309 7327
rect 8343 7293 8355 7327
rect 8297 7287 8355 7293
rect 6420 7228 8248 7256
rect 6420 7216 6426 7228
rect 4341 7191 4399 7197
rect 4341 7188 4353 7191
rect 2004 7160 4353 7188
rect 2004 7148 2010 7160
rect 4341 7157 4353 7160
rect 4387 7157 4399 7191
rect 4341 7151 4399 7157
rect 4890 7148 4896 7200
rect 4948 7148 4954 7200
rect 5350 7148 5356 7200
rect 5408 7148 5414 7200
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5776 7160 5917 7188
rect 5776 7148 5782 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 5905 7151 5963 7157
rect 6457 7191 6515 7197
rect 6457 7157 6469 7191
rect 6503 7188 6515 7191
rect 6730 7188 6736 7200
rect 6503 7160 6736 7188
rect 6503 7157 6515 7160
rect 6457 7151 6515 7157
rect 6730 7148 6736 7160
rect 6788 7148 6794 7200
rect 6914 7148 6920 7200
rect 6972 7188 6978 7200
rect 7469 7191 7527 7197
rect 7469 7188 7481 7191
rect 6972 7160 7481 7188
rect 6972 7148 6978 7160
rect 7469 7157 7481 7160
rect 7515 7188 7527 7191
rect 8312 7188 8340 7287
rect 8570 7188 8576 7200
rect 7515 7160 8576 7188
rect 7515 7157 7527 7160
rect 7469 7151 7527 7157
rect 8570 7148 8576 7160
rect 8628 7148 8634 7200
rect 8662 7148 8668 7200
rect 8720 7148 8726 7200
rect 8956 7188 8984 7432
rect 9490 7420 9496 7472
rect 9548 7420 9554 7472
rect 12820 7460 12848 7491
rect 12986 7488 12992 7491
rect 13044 7488 13050 7500
rect 10718 7432 12848 7460
rect 13173 7463 13231 7469
rect 13173 7429 13185 7463
rect 13219 7429 13231 7463
rect 13173 7423 13231 7429
rect 13188 7392 13216 7423
rect 14274 7420 14280 7472
rect 14332 7420 14338 7472
rect 14458 7420 14464 7472
rect 14516 7469 14522 7472
rect 14516 7463 14535 7469
rect 14523 7429 14535 7463
rect 14568 7460 14596 7500
rect 14645 7497 14657 7531
rect 14691 7528 14703 7531
rect 14734 7528 14740 7540
rect 14691 7500 14740 7528
rect 14691 7497 14703 7500
rect 14645 7491 14703 7497
rect 14734 7488 14740 7500
rect 14792 7488 14798 7540
rect 15723 7531 15781 7537
rect 15723 7528 15735 7531
rect 14844 7500 15735 7528
rect 14844 7460 14872 7500
rect 15723 7497 15735 7500
rect 15769 7497 15781 7531
rect 16853 7531 16911 7537
rect 15723 7491 15781 7497
rect 15856 7500 16252 7528
rect 14568 7432 14872 7460
rect 14516 7423 14535 7429
rect 14516 7420 14522 7423
rect 14918 7420 14924 7472
rect 14976 7420 14982 7472
rect 15102 7420 15108 7472
rect 15160 7469 15166 7472
rect 15160 7463 15179 7469
rect 15167 7429 15179 7463
rect 15160 7423 15179 7429
rect 15160 7420 15166 7423
rect 15378 7420 15384 7472
rect 15436 7460 15442 7472
rect 15856 7460 15884 7500
rect 15436 7432 15884 7460
rect 15933 7463 15991 7469
rect 15436 7420 15442 7432
rect 15933 7429 15945 7463
rect 15979 7460 15991 7463
rect 16022 7460 16028 7472
rect 15979 7432 16028 7460
rect 15979 7429 15991 7432
rect 15933 7423 15991 7429
rect 16022 7420 16028 7432
rect 16080 7420 16086 7472
rect 12636 7364 13216 7392
rect 9214 7284 9220 7336
rect 9272 7284 9278 7336
rect 9582 7284 9588 7336
rect 9640 7324 9646 7336
rect 9858 7324 9864 7336
rect 9640 7296 9864 7324
rect 9640 7284 9646 7296
rect 9858 7284 9864 7296
rect 9916 7324 9922 7336
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 9916 7296 11253 7324
rect 9916 7284 9922 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11241 7287 11299 7293
rect 11606 7284 11612 7336
rect 11664 7284 11670 7336
rect 11882 7284 11888 7336
rect 11940 7284 11946 7336
rect 10502 7216 10508 7268
rect 10560 7256 10566 7268
rect 12636 7256 12664 7364
rect 13538 7352 13544 7404
rect 13596 7352 13602 7404
rect 13633 7395 13691 7401
rect 13633 7361 13645 7395
rect 13679 7392 13691 7395
rect 13722 7392 13728 7404
rect 13679 7364 13728 7392
rect 13679 7361 13691 7364
rect 13633 7355 13691 7361
rect 13722 7352 13728 7364
rect 13780 7352 13786 7404
rect 13817 7395 13875 7401
rect 13817 7361 13829 7395
rect 13863 7392 13875 7395
rect 16114 7392 16120 7404
rect 13863 7364 16120 7392
rect 13863 7361 13875 7364
rect 13817 7355 13875 7361
rect 16114 7352 16120 7364
rect 16172 7352 16178 7404
rect 16224 7401 16252 7500
rect 16853 7497 16865 7531
rect 16899 7528 16911 7531
rect 18877 7531 18935 7537
rect 16899 7500 18828 7528
rect 16899 7497 16911 7500
rect 16853 7491 16911 7497
rect 17402 7420 17408 7472
rect 17460 7420 17466 7472
rect 18800 7460 18828 7500
rect 18877 7497 18889 7531
rect 18923 7528 18935 7531
rect 19794 7528 19800 7540
rect 18923 7500 19800 7528
rect 18923 7497 18935 7500
rect 18877 7491 18935 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 20806 7488 20812 7540
rect 20864 7528 20870 7540
rect 20901 7531 20959 7537
rect 20901 7528 20913 7531
rect 20864 7500 20913 7528
rect 20864 7488 20870 7500
rect 20901 7497 20913 7500
rect 20947 7497 20959 7531
rect 20901 7491 20959 7497
rect 21177 7531 21235 7537
rect 21177 7497 21189 7531
rect 21223 7497 21235 7531
rect 21177 7491 21235 7497
rect 19334 7460 19340 7472
rect 18800 7432 19340 7460
rect 19334 7420 19340 7432
rect 19392 7420 19398 7472
rect 19426 7420 19432 7472
rect 19484 7420 19490 7472
rect 21192 7460 21220 7491
rect 20654 7432 21220 7460
rect 21345 7463 21403 7469
rect 21345 7429 21357 7463
rect 21391 7460 21403 7463
rect 21545 7463 21603 7469
rect 21391 7432 21496 7460
rect 21391 7429 21403 7432
rect 21345 7423 21403 7429
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 16393 7395 16451 7401
rect 16393 7361 16405 7395
rect 16439 7361 16451 7395
rect 16393 7355 16451 7361
rect 12710 7284 12716 7336
rect 12768 7324 12774 7336
rect 15102 7324 15108 7336
rect 12768 7296 15108 7324
rect 12768 7284 12774 7296
rect 15102 7284 15108 7296
rect 15160 7284 15166 7336
rect 15286 7284 15292 7336
rect 15344 7324 15350 7336
rect 16408 7324 16436 7355
rect 18506 7352 18512 7404
rect 18564 7352 18570 7404
rect 15344 7296 16436 7324
rect 15344 7284 15350 7296
rect 16942 7284 16948 7336
rect 17000 7324 17006 7336
rect 17129 7327 17187 7333
rect 17129 7324 17141 7327
rect 17000 7296 17141 7324
rect 17000 7284 17006 7296
rect 17129 7293 17141 7296
rect 17175 7324 17187 7327
rect 19153 7327 19211 7333
rect 19153 7324 19165 7327
rect 17175 7296 19165 7324
rect 17175 7293 17187 7296
rect 17129 7287 17187 7293
rect 19153 7293 19165 7296
rect 19199 7324 19211 7327
rect 21468 7324 21496 7432
rect 21545 7429 21557 7463
rect 21591 7460 21603 7463
rect 21726 7460 21732 7472
rect 21591 7432 21732 7460
rect 21591 7429 21603 7432
rect 21545 7423 21603 7429
rect 21726 7420 21732 7432
rect 21784 7420 21790 7472
rect 22554 7420 22560 7472
rect 22612 7420 22618 7472
rect 24026 7460 24032 7472
rect 23782 7432 24032 7460
rect 24026 7420 24032 7432
rect 24084 7420 24090 7472
rect 22186 7352 22192 7404
rect 22244 7392 22250 7404
rect 22281 7395 22339 7401
rect 22281 7392 22293 7395
rect 22244 7364 22293 7392
rect 22244 7352 22250 7364
rect 22281 7361 22293 7364
rect 22327 7361 22339 7395
rect 22281 7355 22339 7361
rect 22646 7324 22652 7336
rect 19199 7296 19288 7324
rect 21468 7296 22652 7324
rect 19199 7293 19211 7296
rect 19153 7287 19211 7293
rect 10560 7228 12664 7256
rect 13004 7228 15792 7256
rect 10560 7216 10566 7228
rect 13004 7197 13032 7228
rect 12989 7191 13047 7197
rect 12989 7188 13001 7191
rect 8956 7160 13001 7188
rect 12989 7157 13001 7160
rect 13035 7157 13047 7191
rect 12989 7151 13047 7157
rect 14461 7191 14519 7197
rect 14461 7157 14473 7191
rect 14507 7188 14519 7191
rect 15010 7188 15016 7200
rect 14507 7160 15016 7188
rect 14507 7157 14519 7160
rect 14461 7151 14519 7157
rect 15010 7148 15016 7160
rect 15068 7188 15074 7200
rect 15105 7191 15163 7197
rect 15105 7188 15117 7191
rect 15068 7160 15117 7188
rect 15068 7148 15074 7160
rect 15105 7157 15117 7160
rect 15151 7157 15163 7191
rect 15105 7151 15163 7157
rect 15194 7148 15200 7200
rect 15252 7188 15258 7200
rect 15289 7191 15347 7197
rect 15289 7188 15301 7191
rect 15252 7160 15301 7188
rect 15252 7148 15258 7160
rect 15289 7157 15301 7160
rect 15335 7157 15347 7191
rect 15289 7151 15347 7157
rect 15562 7148 15568 7200
rect 15620 7148 15626 7200
rect 15764 7197 15792 7228
rect 19260 7200 19288 7296
rect 22646 7284 22652 7296
rect 22704 7284 22710 7336
rect 22922 7284 22928 7336
rect 22980 7324 22986 7336
rect 24029 7327 24087 7333
rect 24029 7324 24041 7327
rect 22980 7296 24041 7324
rect 22980 7284 22986 7296
rect 24029 7293 24041 7296
rect 24075 7293 24087 7327
rect 24029 7287 24087 7293
rect 21376 7228 22048 7256
rect 15749 7191 15807 7197
rect 15749 7157 15761 7191
rect 15795 7157 15807 7191
rect 15749 7151 15807 7157
rect 15930 7148 15936 7200
rect 15988 7188 15994 7200
rect 16301 7191 16359 7197
rect 16301 7188 16313 7191
rect 15988 7160 16313 7188
rect 15988 7148 15994 7160
rect 16301 7157 16313 7160
rect 16347 7157 16359 7191
rect 16301 7151 16359 7157
rect 19242 7148 19248 7200
rect 19300 7148 19306 7200
rect 21376 7197 21404 7228
rect 21361 7191 21419 7197
rect 21361 7157 21373 7191
rect 21407 7157 21419 7191
rect 21361 7151 21419 7157
rect 21450 7148 21456 7200
rect 21508 7188 21514 7200
rect 21913 7191 21971 7197
rect 21913 7188 21925 7191
rect 21508 7160 21925 7188
rect 21508 7148 21514 7160
rect 21913 7157 21925 7160
rect 21959 7157 21971 7191
rect 22020 7188 22048 7228
rect 22370 7188 22376 7200
rect 22020 7160 22376 7188
rect 21913 7151 21971 7157
rect 22370 7148 22376 7160
rect 22428 7188 22434 7200
rect 23290 7188 23296 7200
rect 22428 7160 23296 7188
rect 22428 7148 22434 7160
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 24397 7191 24455 7197
rect 24397 7157 24409 7191
rect 24443 7188 24455 7191
rect 24578 7188 24584 7200
rect 24443 7160 24584 7188
rect 24443 7157 24455 7160
rect 24397 7151 24455 7157
rect 24578 7148 24584 7160
rect 24636 7148 24642 7200
rect 1104 7098 24840 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 20214 7098
rect 20266 7046 20278 7098
rect 20330 7046 20342 7098
rect 20394 7046 20406 7098
rect 20458 7046 20470 7098
rect 20522 7046 24840 7098
rect 1104 7024 24840 7046
rect 1857 6987 1915 6993
rect 1857 6953 1869 6987
rect 1903 6984 1915 6987
rect 1946 6984 1952 6996
rect 1903 6956 1952 6984
rect 1903 6953 1915 6956
rect 1857 6947 1915 6953
rect 1946 6944 1952 6956
rect 2004 6944 2010 6996
rect 6086 6944 6092 6996
rect 6144 6984 6150 6996
rect 6181 6987 6239 6993
rect 6181 6984 6193 6987
rect 6144 6956 6193 6984
rect 6144 6944 6150 6956
rect 6181 6953 6193 6956
rect 6227 6953 6239 6987
rect 6181 6947 6239 6953
rect 7653 6987 7711 6993
rect 7653 6953 7665 6987
rect 7699 6984 7711 6987
rect 8018 6984 8024 6996
rect 7699 6956 8024 6984
rect 7699 6953 7711 6956
rect 7653 6947 7711 6953
rect 8018 6944 8024 6956
rect 8076 6984 8082 6996
rect 10502 6984 10508 6996
rect 8076 6956 10508 6984
rect 8076 6944 8082 6956
rect 10502 6944 10508 6956
rect 10560 6944 10566 6996
rect 16022 6984 16028 6996
rect 10612 6956 16028 6984
rect 2685 6919 2743 6925
rect 2685 6885 2697 6919
rect 2731 6916 2743 6919
rect 3050 6916 3056 6928
rect 2731 6888 3056 6916
rect 2731 6885 2743 6888
rect 2685 6879 2743 6885
rect 3050 6876 3056 6888
rect 3108 6876 3114 6928
rect 3421 6919 3479 6925
rect 3421 6885 3433 6919
rect 3467 6885 3479 6919
rect 3421 6879 3479 6885
rect 2317 6851 2375 6857
rect 2317 6817 2329 6851
rect 2363 6848 2375 6851
rect 3436 6848 3464 6879
rect 5810 6876 5816 6928
rect 5868 6916 5874 6928
rect 5997 6919 6055 6925
rect 5997 6916 6009 6919
rect 5868 6888 6009 6916
rect 5868 6876 5874 6888
rect 5997 6885 6009 6888
rect 6043 6885 6055 6919
rect 6549 6919 6607 6925
rect 6549 6916 6561 6919
rect 5997 6879 6055 6885
rect 6380 6888 6561 6916
rect 2363 6820 3464 6848
rect 2363 6817 2375 6820
rect 2317 6811 2375 6817
rect 2498 6780 2504 6792
rect 1688 6752 2504 6780
rect 1578 6672 1584 6724
rect 1636 6712 1642 6724
rect 1688 6721 1716 6752
rect 2498 6740 2504 6752
rect 2556 6740 2562 6792
rect 3436 6780 3464 6820
rect 3786 6808 3792 6860
rect 3844 6848 3850 6860
rect 4157 6851 4215 6857
rect 4157 6848 4169 6851
rect 3844 6820 4169 6848
rect 3844 6808 3850 6820
rect 4157 6817 4169 6820
rect 4203 6817 4215 6851
rect 5626 6848 5632 6860
rect 4157 6811 4215 6817
rect 5184 6820 5632 6848
rect 5184 6789 5212 6820
rect 5626 6808 5632 6820
rect 5684 6808 5690 6860
rect 5721 6851 5779 6857
rect 5721 6817 5733 6851
rect 5767 6848 5779 6851
rect 6086 6848 6092 6860
rect 5767 6820 6092 6848
rect 5767 6817 5779 6820
rect 5721 6811 5779 6817
rect 6086 6808 6092 6820
rect 6144 6848 6150 6860
rect 6380 6848 6408 6888
rect 6549 6885 6561 6888
rect 6595 6885 6607 6919
rect 6549 6879 6607 6885
rect 9674 6876 9680 6928
rect 9732 6916 9738 6928
rect 10612 6916 10640 6956
rect 16022 6944 16028 6956
rect 16080 6944 16086 6996
rect 17957 6987 18015 6993
rect 17957 6953 17969 6987
rect 18003 6984 18015 6987
rect 18046 6984 18052 6996
rect 18003 6956 18052 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18417 6987 18475 6993
rect 18417 6953 18429 6987
rect 18463 6984 18475 6987
rect 18966 6984 18972 6996
rect 18463 6956 18972 6984
rect 18463 6953 18475 6956
rect 18417 6947 18475 6953
rect 18966 6944 18972 6956
rect 19024 6944 19030 6996
rect 19610 6944 19616 6996
rect 19668 6944 19674 6996
rect 20070 6944 20076 6996
rect 20128 6984 20134 6996
rect 20330 6987 20388 6993
rect 20330 6984 20342 6987
rect 20128 6956 20342 6984
rect 20128 6944 20134 6956
rect 20330 6953 20342 6956
rect 20376 6953 20388 6987
rect 20330 6947 20388 6953
rect 20898 6944 20904 6996
rect 20956 6984 20962 6996
rect 21821 6987 21879 6993
rect 21821 6984 21833 6987
rect 20956 6956 21833 6984
rect 20956 6944 20962 6956
rect 21821 6953 21833 6956
rect 21867 6953 21879 6987
rect 21821 6947 21879 6953
rect 9732 6888 10640 6916
rect 9732 6876 9738 6888
rect 12066 6876 12072 6928
rect 12124 6916 12130 6928
rect 12161 6919 12219 6925
rect 12161 6916 12173 6919
rect 12124 6888 12173 6916
rect 12124 6876 12130 6888
rect 12161 6885 12173 6888
rect 12207 6885 12219 6919
rect 13722 6916 13728 6928
rect 12161 6879 12219 6885
rect 12268 6888 13728 6916
rect 6144 6820 6408 6848
rect 6457 6851 6515 6857
rect 6144 6808 6150 6820
rect 6457 6817 6469 6851
rect 6503 6817 6515 6851
rect 6457 6811 6515 6817
rect 3881 6783 3939 6789
rect 3881 6780 3893 6783
rect 3436 6752 3893 6780
rect 3881 6749 3893 6752
rect 3927 6749 3939 6783
rect 3881 6743 3939 6749
rect 5169 6783 5227 6789
rect 5169 6749 5181 6783
rect 5215 6749 5227 6783
rect 5169 6743 5227 6749
rect 5261 6783 5319 6789
rect 5261 6749 5273 6783
rect 5307 6749 5319 6783
rect 5261 6743 5319 6749
rect 5353 6783 5411 6789
rect 5353 6749 5365 6783
rect 5399 6780 5411 6783
rect 5902 6780 5908 6792
rect 5399 6752 5908 6780
rect 5399 6749 5411 6752
rect 5353 6743 5411 6749
rect 1673 6715 1731 6721
rect 1673 6712 1685 6715
rect 1636 6684 1685 6712
rect 1636 6672 1642 6684
rect 1673 6681 1685 6684
rect 1719 6681 1731 6715
rect 1673 6675 1731 6681
rect 1889 6715 1947 6721
rect 1889 6681 1901 6715
rect 1935 6712 1947 6715
rect 2130 6712 2136 6724
rect 1935 6684 2136 6712
rect 1935 6681 1947 6684
rect 1889 6675 1947 6681
rect 2130 6672 2136 6684
rect 2188 6672 2194 6724
rect 2866 6712 2872 6724
rect 2424 6684 2872 6712
rect 2041 6647 2099 6653
rect 2041 6613 2053 6647
rect 2087 6644 2099 6647
rect 2424 6644 2452 6684
rect 2866 6672 2872 6684
rect 2924 6672 2930 6724
rect 3050 6672 3056 6724
rect 3108 6712 3114 6724
rect 3108 6684 3648 6712
rect 3108 6672 3114 6684
rect 2087 6616 2452 6644
rect 2087 6613 2099 6616
rect 2041 6607 2099 6613
rect 2774 6604 2780 6656
rect 2832 6604 2838 6656
rect 3510 6604 3516 6656
rect 3568 6604 3574 6656
rect 3620 6644 3648 6684
rect 3786 6672 3792 6724
rect 3844 6712 3850 6724
rect 3896 6712 3924 6743
rect 3844 6684 3924 6712
rect 5276 6712 5304 6743
rect 5902 6740 5908 6752
rect 5960 6780 5966 6792
rect 6472 6780 6500 6811
rect 6730 6808 6736 6860
rect 6788 6848 6794 6860
rect 10321 6851 10379 6857
rect 6788 6820 8524 6848
rect 6788 6808 6794 6820
rect 5960 6752 6500 6780
rect 7745 6783 7803 6789
rect 5960 6740 5966 6752
rect 7745 6749 7757 6783
rect 7791 6749 7803 6783
rect 7745 6743 7803 6749
rect 5276 6684 5672 6712
rect 3844 6672 3850 6684
rect 3970 6644 3976 6656
rect 3620 6616 3976 6644
rect 3970 6604 3976 6616
rect 4028 6604 4034 6656
rect 4985 6647 5043 6653
rect 4985 6613 4997 6647
rect 5031 6644 5043 6647
rect 5534 6644 5540 6656
rect 5031 6616 5540 6644
rect 5031 6613 5043 6616
rect 4985 6607 5043 6613
rect 5534 6604 5540 6616
rect 5592 6604 5598 6656
rect 5644 6644 5672 6684
rect 5810 6672 5816 6724
rect 5868 6712 5874 6724
rect 6546 6712 6552 6724
rect 5868 6684 6552 6712
rect 5868 6672 5874 6684
rect 6546 6672 6552 6684
rect 6604 6712 6610 6724
rect 6917 6715 6975 6721
rect 6917 6712 6929 6715
rect 6604 6684 6929 6712
rect 6604 6672 6610 6684
rect 6917 6681 6929 6684
rect 6963 6681 6975 6715
rect 7760 6712 7788 6743
rect 7834 6740 7840 6792
rect 7892 6780 7898 6792
rect 8496 6789 8524 6820
rect 10321 6817 10333 6851
rect 10367 6848 10379 6851
rect 11146 6848 11152 6860
rect 10367 6820 11152 6848
rect 10367 6817 10379 6820
rect 10321 6811 10379 6817
rect 11146 6808 11152 6820
rect 11204 6808 11210 6860
rect 11698 6808 11704 6860
rect 11756 6848 11762 6860
rect 12268 6848 12296 6888
rect 13722 6876 13728 6888
rect 13780 6876 13786 6928
rect 15470 6876 15476 6928
rect 15528 6916 15534 6928
rect 15930 6916 15936 6928
rect 15528 6888 15936 6916
rect 15528 6876 15534 6888
rect 15930 6876 15936 6888
rect 15988 6876 15994 6928
rect 17586 6876 17592 6928
rect 17644 6916 17650 6928
rect 19518 6916 19524 6928
rect 17644 6888 19524 6916
rect 17644 6876 17650 6888
rect 19518 6876 19524 6888
rect 19576 6876 19582 6928
rect 21836 6916 21864 6947
rect 21836 6888 22232 6916
rect 11756 6820 12296 6848
rect 11756 6808 11762 6820
rect 12618 6808 12624 6860
rect 12676 6848 12682 6860
rect 13173 6851 13231 6857
rect 13173 6848 13185 6851
rect 12676 6820 13185 6848
rect 12676 6808 12682 6820
rect 13173 6817 13185 6820
rect 13219 6817 13231 6851
rect 16209 6851 16267 6857
rect 16209 6848 16221 6851
rect 13173 6811 13231 6817
rect 14108 6820 16221 6848
rect 14108 6792 14136 6820
rect 16209 6817 16221 6820
rect 16255 6848 16267 6851
rect 16942 6848 16948 6860
rect 16255 6820 16948 6848
rect 16255 6817 16267 6820
rect 16209 6811 16267 6817
rect 16942 6808 16948 6820
rect 17000 6808 17006 6860
rect 17034 6808 17040 6860
rect 17092 6848 17098 6860
rect 22094 6848 22100 6860
rect 17092 6820 22100 6848
rect 17092 6808 17098 6820
rect 22094 6808 22100 6820
rect 22152 6808 22158 6860
rect 8205 6783 8263 6789
rect 8205 6780 8217 6783
rect 7892 6752 8217 6780
rect 7892 6740 7898 6752
rect 8205 6749 8217 6752
rect 8251 6749 8263 6783
rect 8205 6743 8263 6749
rect 8481 6783 8539 6789
rect 8481 6749 8493 6783
rect 8527 6749 8539 6783
rect 8481 6743 8539 6749
rect 9033 6783 9091 6789
rect 9033 6749 9045 6783
rect 9079 6780 9091 6783
rect 9674 6780 9680 6792
rect 9079 6752 9680 6780
rect 9079 6749 9091 6752
rect 9033 6743 9091 6749
rect 9674 6740 9680 6752
rect 9732 6740 9738 6792
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 8846 6712 8852 6724
rect 7760 6684 8852 6712
rect 6917 6675 6975 6681
rect 8846 6672 8852 6684
rect 8904 6672 8910 6724
rect 9306 6672 9312 6724
rect 9364 6712 9370 6724
rect 9493 6715 9551 6721
rect 9493 6712 9505 6715
rect 9364 6684 9505 6712
rect 9364 6672 9370 6684
rect 9493 6681 9505 6684
rect 9539 6681 9551 6715
rect 9968 6712 9996 6743
rect 10226 6740 10232 6792
rect 10284 6740 10290 6792
rect 10410 6740 10416 6792
rect 10468 6740 10474 6792
rect 10962 6740 10968 6792
rect 11020 6740 11026 6792
rect 11333 6783 11391 6789
rect 11333 6749 11345 6783
rect 11379 6780 11391 6783
rect 11606 6780 11612 6792
rect 11379 6752 11612 6780
rect 11379 6749 11391 6752
rect 11333 6743 11391 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 11790 6740 11796 6792
rect 11848 6780 11854 6792
rect 11977 6783 12035 6789
rect 11977 6780 11989 6783
rect 11848 6752 11989 6780
rect 11848 6740 11854 6752
rect 11977 6749 11989 6752
rect 12023 6780 12035 6783
rect 12529 6783 12587 6789
rect 12023 6752 12434 6780
rect 12023 6749 12035 6752
rect 11977 6743 12035 6749
rect 10594 6712 10600 6724
rect 9968 6684 10600 6712
rect 9493 6675 9551 6681
rect 10594 6672 10600 6684
rect 10652 6672 10658 6724
rect 12406 6712 12434 6752
rect 12529 6749 12541 6783
rect 12575 6780 12587 6783
rect 12802 6780 12808 6792
rect 12575 6752 12808 6780
rect 12575 6749 12587 6752
rect 12529 6743 12587 6749
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 12897 6783 12955 6789
rect 12897 6749 12909 6783
rect 12943 6749 12955 6783
rect 12897 6743 12955 6749
rect 12912 6712 12940 6743
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 14185 6783 14243 6789
rect 14185 6780 14197 6783
rect 14148 6752 14197 6780
rect 14148 6740 14154 6752
rect 14185 6749 14197 6752
rect 14231 6749 14243 6783
rect 14185 6743 14243 6749
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 18874 6780 18880 6792
rect 18288 6752 18880 6780
rect 18288 6740 18294 6752
rect 12406 6684 12940 6712
rect 12986 6672 12992 6724
rect 13044 6712 13050 6724
rect 13354 6712 13360 6724
rect 13044 6684 13360 6712
rect 13044 6672 13050 6684
rect 13354 6672 13360 6684
rect 13412 6672 13418 6724
rect 14458 6672 14464 6724
rect 14516 6672 14522 6724
rect 15194 6672 15200 6724
rect 15252 6672 15258 6724
rect 16485 6715 16543 6721
rect 16485 6681 16497 6715
rect 16531 6712 16543 6715
rect 16758 6712 16764 6724
rect 16531 6684 16764 6712
rect 16531 6681 16543 6684
rect 16485 6675 16543 6681
rect 16758 6672 16764 6684
rect 16816 6672 16822 6724
rect 18616 6721 18644 6752
rect 18874 6740 18880 6752
rect 18932 6740 18938 6792
rect 19334 6740 19340 6792
rect 19392 6780 19398 6792
rect 19978 6780 19984 6792
rect 19392 6752 19984 6780
rect 19392 6740 19398 6752
rect 19978 6740 19984 6752
rect 20036 6780 20042 6792
rect 20073 6783 20131 6789
rect 20073 6780 20085 6783
rect 20036 6752 20085 6780
rect 20036 6740 20042 6752
rect 20073 6749 20085 6752
rect 20119 6749 20131 6783
rect 22204 6780 22232 6888
rect 22278 6808 22284 6860
rect 22336 6848 22342 6860
rect 22741 6851 22799 6857
rect 22741 6848 22753 6851
rect 22336 6820 22753 6848
rect 22336 6808 22342 6820
rect 22741 6817 22753 6820
rect 22787 6848 22799 6851
rect 23014 6848 23020 6860
rect 22787 6820 23020 6848
rect 22787 6817 22799 6820
rect 22741 6811 22799 6817
rect 23014 6808 23020 6820
rect 23072 6808 23078 6860
rect 23750 6808 23756 6860
rect 23808 6808 23814 6860
rect 23569 6783 23627 6789
rect 23569 6780 23581 6783
rect 22204 6752 23581 6780
rect 20073 6743 20131 6749
rect 23569 6749 23581 6752
rect 23615 6749 23627 6783
rect 23569 6743 23627 6749
rect 18601 6715 18659 6721
rect 17710 6684 18276 6712
rect 6638 6644 6644 6656
rect 5644 6616 6644 6644
rect 6638 6604 6644 6616
rect 6696 6604 6702 6656
rect 8110 6604 8116 6656
rect 8168 6644 8174 6656
rect 8297 6647 8355 6653
rect 8297 6644 8309 6647
rect 8168 6616 8309 6644
rect 8168 6604 8174 6616
rect 8297 6613 8309 6616
rect 8343 6613 8355 6647
rect 8297 6607 8355 6613
rect 8665 6647 8723 6653
rect 8665 6613 8677 6647
rect 8711 6644 8723 6647
rect 8754 6644 8760 6656
rect 8711 6616 8760 6644
rect 8711 6613 8723 6616
rect 8665 6607 8723 6613
rect 8754 6604 8760 6616
rect 8812 6604 8818 6656
rect 15933 6647 15991 6653
rect 15933 6613 15945 6647
rect 15979 6644 15991 6647
rect 17218 6644 17224 6656
rect 15979 6616 17224 6644
rect 15979 6613 15991 6616
rect 15933 6607 15991 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 18248 6653 18276 6684
rect 18601 6681 18613 6715
rect 18647 6681 18659 6715
rect 18601 6675 18659 6681
rect 19705 6715 19763 6721
rect 19705 6681 19717 6715
rect 19751 6712 19763 6715
rect 19886 6712 19892 6724
rect 19751 6684 19892 6712
rect 19751 6681 19763 6684
rect 19705 6675 19763 6681
rect 19886 6672 19892 6684
rect 19944 6672 19950 6724
rect 21358 6672 21364 6724
rect 21416 6672 21422 6724
rect 22465 6715 22523 6721
rect 22465 6712 22477 6715
rect 21652 6684 22477 6712
rect 18414 6653 18420 6656
rect 18233 6647 18291 6653
rect 18233 6613 18245 6647
rect 18279 6613 18291 6647
rect 18233 6607 18291 6613
rect 18391 6647 18420 6653
rect 18391 6613 18403 6647
rect 18391 6607 18420 6613
rect 18414 6604 18420 6607
rect 18472 6604 18478 6656
rect 18966 6604 18972 6656
rect 19024 6604 19030 6656
rect 20070 6604 20076 6656
rect 20128 6644 20134 6656
rect 21652 6644 21680 6684
rect 22465 6681 22477 6684
rect 22511 6681 22523 6715
rect 22465 6675 22523 6681
rect 20128 6616 21680 6644
rect 20128 6604 20134 6616
rect 22002 6604 22008 6656
rect 22060 6644 22066 6656
rect 22097 6647 22155 6653
rect 22097 6644 22109 6647
rect 22060 6616 22109 6644
rect 22060 6604 22066 6616
rect 22097 6613 22109 6616
rect 22143 6613 22155 6647
rect 22097 6607 22155 6613
rect 22557 6647 22615 6653
rect 22557 6613 22569 6647
rect 22603 6644 22615 6647
rect 23014 6644 23020 6656
rect 22603 6616 23020 6644
rect 22603 6613 22615 6616
rect 22557 6607 22615 6613
rect 23014 6604 23020 6616
rect 23072 6604 23078 6656
rect 23106 6604 23112 6656
rect 23164 6604 23170 6656
rect 23290 6604 23296 6656
rect 23348 6644 23354 6656
rect 23477 6647 23535 6653
rect 23477 6644 23489 6647
rect 23348 6616 23489 6644
rect 23348 6604 23354 6616
rect 23477 6613 23489 6616
rect 23523 6613 23535 6647
rect 23477 6607 23535 6613
rect 1104 6554 24840 6576
rect 1104 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 24214 6554
rect 24266 6502 24278 6554
rect 24330 6502 24342 6554
rect 24394 6502 24406 6554
rect 24458 6502 24470 6554
rect 24522 6502 24840 6554
rect 1104 6480 24840 6502
rect 1688 6412 4660 6440
rect 1688 6313 1716 6412
rect 1964 6344 2728 6372
rect 1964 6313 1992 6344
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6273 1731 6307
rect 1673 6267 1731 6273
rect 1949 6307 2007 6313
rect 1949 6273 1961 6307
rect 1995 6273 2007 6307
rect 1949 6267 2007 6273
rect 1581 6239 1639 6245
rect 1581 6205 1593 6239
rect 1627 6236 1639 6239
rect 1964 6236 1992 6267
rect 2314 6264 2320 6316
rect 2372 6264 2378 6316
rect 2593 6307 2651 6313
rect 2593 6273 2605 6307
rect 2639 6273 2651 6307
rect 2700 6304 2728 6344
rect 2774 6332 2780 6384
rect 2832 6372 2838 6384
rect 2832 6344 3832 6372
rect 2832 6332 2838 6344
rect 2869 6307 2927 6313
rect 2869 6304 2881 6307
rect 2700 6276 2881 6304
rect 2593 6267 2651 6273
rect 2869 6273 2881 6276
rect 2915 6273 2927 6307
rect 2869 6267 2927 6273
rect 1627 6208 1992 6236
rect 1627 6205 1639 6208
rect 1581 6199 1639 6205
rect 2406 6196 2412 6248
rect 2464 6196 2470 6248
rect 2608 6236 2636 6267
rect 3510 6264 3516 6316
rect 3568 6304 3574 6316
rect 3804 6313 3832 6344
rect 3697 6307 3755 6313
rect 3697 6304 3709 6307
rect 3568 6276 3709 6304
rect 3568 6264 3574 6276
rect 3697 6273 3709 6276
rect 3743 6273 3755 6307
rect 3697 6267 3755 6273
rect 3789 6307 3847 6313
rect 3789 6273 3801 6307
rect 3835 6273 3847 6307
rect 4632 6304 4660 6412
rect 6638 6400 6644 6452
rect 6696 6440 6702 6452
rect 6825 6443 6883 6449
rect 6825 6440 6837 6443
rect 6696 6412 6837 6440
rect 6696 6400 6702 6412
rect 6825 6409 6837 6412
rect 6871 6409 6883 6443
rect 6825 6403 6883 6409
rect 7285 6443 7343 6449
rect 7285 6409 7297 6443
rect 7331 6440 7343 6443
rect 7558 6440 7564 6452
rect 7331 6412 7564 6440
rect 7331 6409 7343 6412
rect 7285 6403 7343 6409
rect 7558 6400 7564 6412
rect 7616 6400 7622 6452
rect 8110 6440 8116 6452
rect 7668 6412 8116 6440
rect 6730 6332 6736 6384
rect 6788 6372 6794 6384
rect 7668 6381 7696 6412
rect 8110 6400 8116 6412
rect 8168 6440 8174 6452
rect 8297 6443 8355 6449
rect 8297 6440 8309 6443
rect 8168 6412 8309 6440
rect 8168 6400 8174 6412
rect 8297 6409 8309 6412
rect 8343 6409 8355 6443
rect 8297 6403 8355 6409
rect 8570 6400 8576 6452
rect 8628 6440 8634 6452
rect 8938 6440 8944 6452
rect 8628 6412 8944 6440
rect 8628 6400 8634 6412
rect 8938 6400 8944 6412
rect 8996 6440 9002 6452
rect 9398 6440 9404 6452
rect 8996 6412 9404 6440
rect 8996 6400 9002 6412
rect 9398 6400 9404 6412
rect 9456 6400 9462 6452
rect 9677 6443 9735 6449
rect 9677 6409 9689 6443
rect 9723 6440 9735 6443
rect 10226 6440 10232 6452
rect 9723 6412 10232 6440
rect 9723 6409 9735 6412
rect 9677 6403 9735 6409
rect 10226 6400 10232 6412
rect 10284 6400 10290 6452
rect 14090 6440 14096 6452
rect 11808 6412 14096 6440
rect 7653 6375 7711 6381
rect 6788 6344 7604 6372
rect 6788 6332 6794 6344
rect 4709 6307 4767 6313
rect 4709 6304 4721 6307
rect 4632 6276 4721 6304
rect 3789 6267 3847 6273
rect 4709 6273 4721 6276
rect 4755 6273 4767 6307
rect 4709 6267 4767 6273
rect 3142 6236 3148 6248
rect 2608 6208 3148 6236
rect 3142 6196 3148 6208
rect 3200 6196 3206 6248
rect 3712 6168 3740 6267
rect 4724 6236 4752 6267
rect 4982 6264 4988 6316
rect 5040 6264 5046 6316
rect 5350 6264 5356 6316
rect 5408 6304 5414 6316
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5408 6276 5549 6304
rect 5408 6264 5414 6276
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 5537 6267 5595 6273
rect 5994 6264 6000 6316
rect 6052 6304 6058 6316
rect 6457 6307 6515 6313
rect 6457 6304 6469 6307
rect 6052 6276 6469 6304
rect 6052 6264 6058 6276
rect 6457 6273 6469 6276
rect 6503 6273 6515 6307
rect 6457 6267 6515 6273
rect 6546 6264 6552 6316
rect 6604 6304 6610 6316
rect 6604 6276 6649 6304
rect 6604 6264 6610 6276
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7101 6307 7159 6313
rect 7101 6304 7113 6307
rect 7064 6276 7113 6304
rect 7064 6264 7070 6276
rect 7101 6273 7113 6276
rect 7147 6273 7159 6307
rect 7101 6267 7159 6273
rect 7190 6264 7196 6316
rect 7248 6304 7254 6316
rect 7576 6313 7604 6344
rect 7653 6341 7665 6375
rect 7699 6341 7711 6375
rect 7653 6335 7711 6341
rect 7834 6332 7840 6384
rect 7892 6332 7898 6384
rect 9214 6332 9220 6384
rect 9272 6372 9278 6384
rect 11808 6372 11836 6412
rect 14090 6400 14096 6412
rect 14148 6400 14154 6452
rect 14458 6400 14464 6452
rect 14516 6440 14522 6452
rect 14645 6443 14703 6449
rect 14645 6440 14657 6443
rect 14516 6412 14657 6440
rect 14516 6400 14522 6412
rect 14645 6409 14657 6412
rect 14691 6409 14703 6443
rect 15562 6440 15568 6452
rect 14645 6403 14703 6409
rect 14936 6412 15568 6440
rect 14936 6372 14964 6412
rect 15562 6400 15568 6412
rect 15620 6400 15626 6452
rect 16758 6400 16764 6452
rect 16816 6400 16822 6452
rect 17218 6400 17224 6452
rect 17276 6400 17282 6452
rect 17862 6400 17868 6452
rect 17920 6400 17926 6452
rect 19153 6443 19211 6449
rect 19153 6409 19165 6443
rect 19199 6440 19211 6443
rect 20714 6440 20720 6452
rect 19199 6412 20720 6440
rect 19199 6409 19211 6412
rect 19153 6403 19211 6409
rect 20714 6400 20720 6412
rect 20772 6400 20778 6452
rect 22094 6440 22100 6452
rect 20824 6412 22100 6440
rect 9272 6344 11836 6372
rect 13294 6344 14964 6372
rect 15013 6375 15071 6381
rect 9272 6332 9278 6344
rect 7285 6307 7343 6313
rect 7285 6304 7297 6307
rect 7248 6276 7297 6304
rect 7248 6264 7254 6276
rect 7285 6273 7297 6276
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7561 6307 7619 6313
rect 7561 6273 7573 6307
rect 7607 6273 7619 6307
rect 7561 6267 7619 6273
rect 8573 6307 8631 6313
rect 8573 6273 8585 6307
rect 8619 6304 8631 6307
rect 8619 6276 9352 6304
rect 8619 6273 8631 6276
rect 8573 6267 8631 6273
rect 9324 6248 9352 6276
rect 9398 6264 9404 6316
rect 9456 6264 9462 6316
rect 9674 6264 9680 6316
rect 9732 6304 9738 6316
rect 10443 6307 10501 6313
rect 10443 6304 10455 6307
rect 9732 6276 10455 6304
rect 9732 6264 9738 6276
rect 10443 6273 10455 6276
rect 10489 6273 10501 6307
rect 10443 6267 10501 6273
rect 10594 6264 10600 6316
rect 10652 6264 10658 6316
rect 10962 6264 10968 6316
rect 11020 6264 11026 6316
rect 11808 6313 11836 6344
rect 15013 6341 15025 6375
rect 15059 6372 15071 6375
rect 17236 6372 17264 6400
rect 18046 6372 18052 6384
rect 15059 6344 17264 6372
rect 17696 6344 18052 6372
rect 15059 6341 15071 6344
rect 15013 6335 15071 6341
rect 11793 6307 11851 6313
rect 11793 6273 11805 6307
rect 11839 6273 11851 6307
rect 11793 6267 11851 6273
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13412 6276 13584 6304
rect 13412 6264 13418 6276
rect 5626 6236 5632 6248
rect 4724 6208 5632 6236
rect 5626 6196 5632 6208
rect 5684 6236 5690 6248
rect 5902 6236 5908 6248
rect 5684 6208 5908 6236
rect 5684 6196 5690 6208
rect 5902 6196 5908 6208
rect 5960 6196 5966 6248
rect 8481 6239 8539 6245
rect 8481 6205 8493 6239
rect 8527 6205 8539 6239
rect 8481 6199 8539 6205
rect 5166 6168 5172 6180
rect 3712 6140 5172 6168
rect 5166 6128 5172 6140
rect 5224 6128 5230 6180
rect 5442 6128 5448 6180
rect 5500 6128 5506 6180
rect 8496 6168 8524 6199
rect 9306 6196 9312 6248
rect 9364 6196 9370 6248
rect 9953 6239 10011 6245
rect 9953 6236 9965 6239
rect 9416 6208 9965 6236
rect 9416 6168 9444 6208
rect 9953 6205 9965 6208
rect 9999 6236 10011 6239
rect 10229 6239 10287 6245
rect 10229 6236 10241 6239
rect 9999 6208 10241 6236
rect 9999 6205 10011 6208
rect 9953 6199 10011 6205
rect 10229 6205 10241 6208
rect 10275 6205 10287 6239
rect 10229 6199 10287 6205
rect 8496 6140 9444 6168
rect 8588 6112 8616 6140
rect 3050 6060 3056 6112
rect 3108 6060 3114 6112
rect 6086 6060 6092 6112
rect 6144 6060 6150 6112
rect 7558 6060 7564 6112
rect 7616 6060 7622 6112
rect 8570 6060 8576 6112
rect 8628 6060 8634 6112
rect 9030 6060 9036 6112
rect 9088 6100 9094 6112
rect 10980 6100 11008 6264
rect 12066 6196 12072 6248
rect 12124 6196 12130 6248
rect 13556 6245 13584 6276
rect 14366 6264 14372 6316
rect 14424 6304 14430 6316
rect 15102 6304 15108 6316
rect 14424 6276 15108 6304
rect 14424 6264 14430 6276
rect 15102 6264 15108 6276
rect 15160 6264 15166 6316
rect 15657 6307 15715 6313
rect 15657 6304 15669 6307
rect 15212 6276 15669 6304
rect 13541 6239 13599 6245
rect 13541 6205 13553 6239
rect 13587 6236 13599 6239
rect 13817 6239 13875 6245
rect 13817 6236 13829 6239
rect 13587 6208 13829 6236
rect 13587 6205 13599 6208
rect 13541 6199 13599 6205
rect 13817 6205 13829 6208
rect 13863 6205 13875 6239
rect 13817 6199 13875 6205
rect 13906 6196 13912 6248
rect 13964 6236 13970 6248
rect 15212 6236 15240 6276
rect 15657 6273 15669 6276
rect 15703 6273 15715 6307
rect 15657 6267 15715 6273
rect 15838 6264 15844 6316
rect 15896 6264 15902 6316
rect 16393 6307 16451 6313
rect 16393 6273 16405 6307
rect 16439 6304 16451 6307
rect 16942 6304 16948 6316
rect 16439 6276 16948 6304
rect 16439 6273 16451 6276
rect 16393 6267 16451 6273
rect 16942 6264 16948 6276
rect 17000 6264 17006 6316
rect 17129 6307 17187 6313
rect 17129 6273 17141 6307
rect 17175 6304 17187 6307
rect 17696 6304 17724 6344
rect 18046 6332 18052 6344
rect 18104 6332 18110 6384
rect 20824 6372 20852 6412
rect 22094 6400 22100 6412
rect 22152 6400 22158 6452
rect 23106 6440 23112 6452
rect 22296 6412 23112 6440
rect 19720 6344 20852 6372
rect 19720 6316 19748 6344
rect 21082 6332 21088 6384
rect 21140 6372 21146 6384
rect 21177 6375 21235 6381
rect 21177 6372 21189 6375
rect 21140 6344 21189 6372
rect 21140 6332 21146 6344
rect 21177 6341 21189 6344
rect 21223 6341 21235 6375
rect 21177 6335 21235 6341
rect 21393 6375 21451 6381
rect 21393 6341 21405 6375
rect 21439 6372 21451 6375
rect 21542 6372 21548 6384
rect 21439 6344 21548 6372
rect 21439 6341 21451 6344
rect 21393 6335 21451 6341
rect 21542 6332 21548 6344
rect 21600 6332 21606 6384
rect 22296 6381 22324 6412
rect 23106 6400 23112 6412
rect 23164 6400 23170 6452
rect 24026 6400 24032 6452
rect 24084 6400 24090 6452
rect 22281 6375 22339 6381
rect 22281 6341 22293 6375
rect 22327 6341 22339 6375
rect 23934 6372 23940 6384
rect 23506 6344 23940 6372
rect 22281 6335 22339 6341
rect 23934 6332 23940 6344
rect 23992 6332 23998 6384
rect 24181 6375 24239 6381
rect 24181 6372 24193 6375
rect 24044 6344 24193 6372
rect 17175 6276 17724 6304
rect 17175 6273 17187 6276
rect 17129 6267 17187 6273
rect 17954 6264 17960 6316
rect 18012 6264 18018 6316
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 13964 6208 15240 6236
rect 15289 6239 15347 6245
rect 13964 6196 13970 6208
rect 15289 6205 15301 6239
rect 15335 6236 15347 6239
rect 17405 6239 17463 6245
rect 17405 6236 17417 6239
rect 15335 6208 17417 6236
rect 15335 6205 15347 6208
rect 15289 6199 15347 6205
rect 17405 6205 17417 6208
rect 17451 6236 17463 6239
rect 17494 6236 17500 6248
rect 17451 6208 17500 6236
rect 17451 6205 17463 6208
rect 17405 6199 17463 6205
rect 17494 6196 17500 6208
rect 17552 6196 17558 6248
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18340 6236 18368 6267
rect 18506 6264 18512 6316
rect 18564 6264 18570 6316
rect 19702 6304 19708 6316
rect 18892 6276 19708 6304
rect 18892 6245 18920 6276
rect 19702 6264 19708 6276
rect 19760 6264 19766 6316
rect 20717 6307 20775 6313
rect 20717 6273 20729 6307
rect 20763 6304 20775 6307
rect 20806 6304 20812 6316
rect 20763 6276 20812 6304
rect 20763 6273 20775 6276
rect 20717 6267 20775 6273
rect 20806 6264 20812 6276
rect 20864 6264 20870 6316
rect 17828 6208 18368 6236
rect 18877 6239 18935 6245
rect 17828 6196 17834 6208
rect 18877 6205 18889 6239
rect 18923 6205 18935 6239
rect 18877 6199 18935 6205
rect 19058 6196 19064 6248
rect 19116 6196 19122 6248
rect 19334 6196 19340 6248
rect 19392 6236 19398 6248
rect 19794 6236 19800 6248
rect 19392 6208 19800 6236
rect 19392 6196 19398 6208
rect 19794 6196 19800 6208
rect 19852 6236 19858 6248
rect 20165 6239 20223 6245
rect 20165 6236 20177 6239
rect 19852 6208 20177 6236
rect 19852 6196 19858 6208
rect 20165 6205 20177 6208
rect 20211 6205 20223 6239
rect 20165 6199 20223 6205
rect 22005 6239 22063 6245
rect 22005 6205 22017 6239
rect 22051 6236 22063 6239
rect 22370 6236 22376 6248
rect 22051 6208 22376 6236
rect 22051 6205 22063 6208
rect 22005 6199 22063 6205
rect 22370 6196 22376 6208
rect 22428 6196 22434 6248
rect 22646 6196 22652 6248
rect 22704 6236 22710 6248
rect 24044 6236 24072 6344
rect 24181 6341 24193 6344
rect 24227 6341 24239 6375
rect 24181 6335 24239 6341
rect 24397 6375 24455 6381
rect 24397 6341 24409 6375
rect 24443 6372 24455 6375
rect 24670 6372 24676 6384
rect 24443 6344 24676 6372
rect 24443 6341 24455 6344
rect 24397 6335 24455 6341
rect 24670 6332 24676 6344
rect 24728 6332 24734 6384
rect 22704 6208 24072 6236
rect 22704 6196 22710 6208
rect 13998 6128 14004 6180
rect 14056 6168 14062 6180
rect 15657 6171 15715 6177
rect 15657 6168 15669 6171
rect 14056 6140 15669 6168
rect 14056 6128 14062 6140
rect 15657 6137 15669 6140
rect 15703 6137 15715 6171
rect 15657 6131 15715 6137
rect 16850 6128 16856 6180
rect 16908 6168 16914 6180
rect 18325 6171 18383 6177
rect 18325 6168 18337 6171
rect 16908 6140 18337 6168
rect 16908 6128 16914 6140
rect 18325 6137 18337 6140
rect 18371 6137 18383 6171
rect 18325 6131 18383 6137
rect 18966 6128 18972 6180
rect 19024 6168 19030 6180
rect 19024 6140 22094 6168
rect 19024 6128 19030 6140
rect 9088 6072 11008 6100
rect 11057 6103 11115 6109
rect 9088 6060 9094 6072
rect 11057 6069 11069 6103
rect 11103 6100 11115 6103
rect 13354 6100 13360 6112
rect 11103 6072 13360 6100
rect 11103 6069 11115 6072
rect 11057 6063 11115 6069
rect 13354 6060 13360 6072
rect 13412 6060 13418 6112
rect 14274 6060 14280 6112
rect 14332 6060 14338 6112
rect 16209 6103 16267 6109
rect 16209 6069 16221 6103
rect 16255 6100 16267 6103
rect 16666 6100 16672 6112
rect 16255 6072 16672 6100
rect 16255 6069 16267 6072
rect 16209 6063 16267 6069
rect 16666 6060 16672 6072
rect 16724 6060 16730 6112
rect 16942 6060 16948 6112
rect 17000 6100 17006 6112
rect 19334 6100 19340 6112
rect 17000 6072 19340 6100
rect 17000 6060 17006 6072
rect 19334 6060 19340 6072
rect 19392 6060 19398 6112
rect 19518 6060 19524 6112
rect 19576 6060 19582 6112
rect 21174 6060 21180 6112
rect 21232 6100 21238 6112
rect 21361 6103 21419 6109
rect 21361 6100 21373 6103
rect 21232 6072 21373 6100
rect 21232 6060 21238 6072
rect 21361 6069 21373 6072
rect 21407 6069 21419 6103
rect 21361 6063 21419 6069
rect 21545 6103 21603 6109
rect 21545 6069 21557 6103
rect 21591 6100 21603 6103
rect 21634 6100 21640 6112
rect 21591 6072 21640 6100
rect 21591 6069 21603 6072
rect 21545 6063 21603 6069
rect 21634 6060 21640 6072
rect 21692 6060 21698 6112
rect 22066 6100 22094 6140
rect 23382 6128 23388 6180
rect 23440 6168 23446 6180
rect 23440 6140 24256 6168
rect 23440 6128 23446 6140
rect 22278 6100 22284 6112
rect 22066 6072 22284 6100
rect 22278 6060 22284 6072
rect 22336 6060 22342 6112
rect 23290 6060 23296 6112
rect 23348 6100 23354 6112
rect 24228 6109 24256 6140
rect 23753 6103 23811 6109
rect 23753 6100 23765 6103
rect 23348 6072 23765 6100
rect 23348 6060 23354 6072
rect 23753 6069 23765 6072
rect 23799 6069 23811 6103
rect 23753 6063 23811 6069
rect 24213 6103 24271 6109
rect 24213 6069 24225 6103
rect 24259 6069 24271 6103
rect 24213 6063 24271 6069
rect 1104 6010 24840 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 20214 6010
rect 20266 5958 20278 6010
rect 20330 5958 20342 6010
rect 20394 5958 20406 6010
rect 20458 5958 20470 6010
rect 20522 5958 24840 6010
rect 1104 5936 24840 5958
rect 2314 5856 2320 5908
rect 2372 5896 2378 5908
rect 4065 5899 4123 5905
rect 4065 5896 4077 5899
rect 2372 5868 4077 5896
rect 2372 5856 2378 5868
rect 4065 5865 4077 5868
rect 4111 5896 4123 5899
rect 4982 5896 4988 5908
rect 4111 5868 4988 5896
rect 4111 5865 4123 5868
rect 4065 5859 4123 5865
rect 4982 5856 4988 5868
rect 5040 5856 5046 5908
rect 5442 5856 5448 5908
rect 5500 5896 5506 5908
rect 5500 5868 6868 5896
rect 5500 5856 5506 5868
rect 3970 5788 3976 5840
rect 4028 5788 4034 5840
rect 2222 5720 2228 5772
rect 2280 5720 2286 5772
rect 3988 5760 4016 5788
rect 4249 5763 4307 5769
rect 4249 5760 4261 5763
rect 2746 5732 3280 5760
rect 3988 5732 4261 5760
rect 1762 5652 1768 5704
rect 1820 5652 1826 5704
rect 2038 5652 2044 5704
rect 2096 5692 2102 5704
rect 2133 5695 2191 5701
rect 2133 5692 2145 5695
rect 2096 5664 2145 5692
rect 2096 5652 2102 5664
rect 2133 5661 2145 5664
rect 2179 5692 2191 5695
rect 2746 5692 2774 5732
rect 2179 5664 2774 5692
rect 2961 5695 3019 5701
rect 2179 5661 2191 5664
rect 2133 5655 2191 5661
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 3050 5692 3056 5704
rect 3007 5664 3056 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3050 5652 3056 5664
rect 3108 5652 3114 5704
rect 3145 5695 3203 5701
rect 3145 5661 3157 5695
rect 3191 5661 3203 5695
rect 3145 5655 3203 5661
rect 1780 5556 1808 5652
rect 2406 5584 2412 5636
rect 2464 5624 2470 5636
rect 3160 5624 3188 5655
rect 2464 5596 3188 5624
rect 3252 5624 3280 5732
rect 4249 5729 4261 5732
rect 4295 5729 4307 5763
rect 5000 5760 5028 5856
rect 5534 5788 5540 5840
rect 5592 5828 5598 5840
rect 5592 5800 6592 5828
rect 5592 5788 5598 5800
rect 4249 5723 4307 5729
rect 4724 5732 4936 5760
rect 5000 5732 5120 5760
rect 3786 5652 3792 5704
rect 3844 5692 3850 5704
rect 3973 5695 4031 5701
rect 3973 5692 3985 5695
rect 3844 5664 3985 5692
rect 3844 5652 3850 5664
rect 3973 5661 3985 5664
rect 4019 5661 4031 5695
rect 3973 5655 4031 5661
rect 4062 5652 4068 5704
rect 4120 5692 4126 5704
rect 4724 5692 4752 5732
rect 4120 5664 4752 5692
rect 4801 5695 4859 5701
rect 4120 5652 4126 5664
rect 4801 5661 4813 5695
rect 4847 5661 4859 5695
rect 4908 5692 4936 5732
rect 4985 5695 5043 5701
rect 4985 5692 4997 5695
rect 4908 5664 4997 5692
rect 4801 5655 4859 5661
rect 4985 5661 4997 5664
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 4080 5624 4108 5652
rect 4816 5624 4844 5655
rect 3252 5596 4108 5624
rect 4264 5596 4844 5624
rect 5092 5624 5120 5732
rect 5736 5732 6408 5760
rect 5736 5704 5764 5732
rect 5166 5652 5172 5704
rect 5224 5692 5230 5704
rect 5445 5695 5503 5701
rect 5445 5692 5457 5695
rect 5224 5664 5457 5692
rect 5224 5652 5230 5664
rect 5445 5661 5457 5664
rect 5491 5661 5503 5695
rect 5445 5655 5503 5661
rect 5534 5652 5540 5704
rect 5592 5692 5598 5704
rect 5592 5664 5637 5692
rect 5592 5652 5598 5664
rect 5718 5652 5724 5704
rect 5776 5652 5782 5704
rect 5902 5652 5908 5704
rect 5960 5701 5966 5704
rect 6380 5701 6408 5732
rect 6564 5701 6592 5800
rect 6840 5769 6868 5868
rect 7834 5856 7840 5908
rect 7892 5896 7898 5908
rect 8205 5899 8263 5905
rect 8205 5896 8217 5899
rect 7892 5868 8217 5896
rect 7892 5856 7898 5868
rect 7944 5769 7972 5868
rect 8205 5865 8217 5868
rect 8251 5865 8263 5899
rect 9306 5896 9312 5908
rect 8205 5859 8263 5865
rect 8404 5868 9312 5896
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5729 6883 5763
rect 7285 5763 7343 5769
rect 7285 5760 7297 5763
rect 6825 5723 6883 5729
rect 6932 5732 7297 5760
rect 5960 5692 5968 5701
rect 6365 5695 6423 5701
rect 5960 5664 6005 5692
rect 5960 5655 5968 5664
rect 6365 5661 6377 5695
rect 6411 5661 6423 5695
rect 6365 5655 6423 5661
rect 6549 5695 6607 5701
rect 6549 5661 6561 5695
rect 6595 5661 6607 5695
rect 6549 5655 6607 5661
rect 5960 5652 5966 5655
rect 6730 5652 6736 5704
rect 6788 5692 6794 5704
rect 6932 5692 6960 5732
rect 7285 5729 7297 5732
rect 7331 5729 7343 5763
rect 7285 5723 7343 5729
rect 7929 5763 7987 5769
rect 7929 5729 7941 5763
rect 7975 5729 7987 5763
rect 7929 5723 7987 5729
rect 6788 5664 6960 5692
rect 7009 5695 7067 5701
rect 6788 5652 6794 5664
rect 7009 5661 7021 5695
rect 7055 5661 7067 5695
rect 7009 5655 7067 5661
rect 7653 5695 7711 5701
rect 7653 5661 7665 5695
rect 7699 5692 7711 5695
rect 8110 5692 8116 5704
rect 7699 5664 8116 5692
rect 7699 5661 7711 5664
rect 7653 5655 7711 5661
rect 5813 5627 5871 5633
rect 5813 5624 5825 5627
rect 5092 5596 5825 5624
rect 2464 5584 2470 5596
rect 4264 5556 4292 5596
rect 5813 5593 5825 5596
rect 5859 5593 5871 5627
rect 5813 5587 5871 5593
rect 6454 5584 6460 5636
rect 6512 5624 6518 5636
rect 7024 5624 7052 5655
rect 8110 5652 8116 5664
rect 8168 5652 8174 5704
rect 8404 5701 8432 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 12066 5856 12072 5908
rect 12124 5896 12130 5908
rect 12253 5899 12311 5905
rect 12253 5896 12265 5899
rect 12124 5868 12265 5896
rect 12124 5856 12130 5868
rect 12253 5865 12265 5868
rect 12299 5865 12311 5899
rect 12253 5859 12311 5865
rect 16853 5899 16911 5905
rect 16853 5865 16865 5899
rect 16899 5896 16911 5899
rect 17126 5896 17132 5908
rect 16899 5868 17132 5896
rect 16899 5865 16911 5868
rect 16853 5859 16911 5865
rect 17126 5856 17132 5868
rect 17184 5896 17190 5908
rect 17678 5896 17684 5908
rect 17184 5868 17684 5896
rect 17184 5856 17190 5868
rect 17678 5856 17684 5868
rect 17736 5896 17742 5908
rect 17773 5899 17831 5905
rect 17773 5896 17785 5899
rect 17736 5868 17785 5896
rect 17736 5856 17742 5868
rect 17773 5865 17785 5868
rect 17819 5865 17831 5899
rect 17773 5859 17831 5865
rect 19429 5899 19487 5905
rect 19429 5865 19441 5899
rect 19475 5896 19487 5899
rect 19610 5896 19616 5908
rect 19475 5868 19616 5896
rect 19475 5865 19487 5868
rect 19429 5859 19487 5865
rect 19610 5856 19616 5868
rect 19668 5856 19674 5908
rect 19889 5899 19947 5905
rect 19889 5865 19901 5899
rect 19935 5896 19947 5899
rect 20070 5896 20076 5908
rect 19935 5868 20076 5896
rect 19935 5865 19947 5868
rect 19889 5859 19947 5865
rect 20070 5856 20076 5868
rect 20128 5856 20134 5908
rect 20622 5896 20628 5908
rect 20180 5868 20628 5896
rect 8570 5788 8576 5840
rect 8628 5788 8634 5840
rect 8846 5788 8852 5840
rect 8904 5828 8910 5840
rect 11698 5828 11704 5840
rect 8904 5800 11704 5828
rect 8904 5788 8910 5800
rect 11698 5788 11704 5800
rect 11756 5788 11762 5840
rect 11974 5788 11980 5840
rect 12032 5828 12038 5840
rect 14185 5831 14243 5837
rect 14185 5828 14197 5831
rect 12032 5800 14197 5828
rect 12032 5788 12038 5800
rect 14185 5797 14197 5800
rect 14231 5797 14243 5831
rect 15654 5828 15660 5840
rect 14185 5791 14243 5797
rect 15028 5800 15660 5828
rect 8588 5760 8616 5788
rect 10318 5760 10324 5772
rect 8496 5732 8616 5760
rect 9232 5732 10324 5760
rect 8496 5701 8524 5732
rect 8389 5695 8447 5701
rect 8389 5661 8401 5695
rect 8435 5661 8447 5695
rect 8389 5655 8447 5661
rect 8481 5695 8539 5701
rect 8481 5661 8493 5695
rect 8527 5661 8539 5695
rect 8481 5655 8539 5661
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5692 8631 5695
rect 8938 5692 8944 5704
rect 8619 5664 8944 5692
rect 8619 5661 8631 5664
rect 8573 5655 8631 5661
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9232 5701 9260 5732
rect 10318 5720 10324 5732
rect 10376 5720 10382 5772
rect 11882 5720 11888 5772
rect 11940 5760 11946 5772
rect 15028 5760 15056 5800
rect 15654 5788 15660 5800
rect 15712 5788 15718 5840
rect 17402 5788 17408 5840
rect 17460 5828 17466 5840
rect 18322 5828 18328 5840
rect 17460 5800 18328 5828
rect 17460 5788 17466 5800
rect 18322 5788 18328 5800
rect 18380 5828 18386 5840
rect 20180 5828 20208 5868
rect 20622 5856 20628 5868
rect 20680 5856 20686 5908
rect 20990 5856 20996 5908
rect 21048 5896 21054 5908
rect 21913 5899 21971 5905
rect 21913 5896 21925 5899
rect 21048 5868 21925 5896
rect 21048 5856 21054 5868
rect 21913 5865 21925 5868
rect 21959 5865 21971 5899
rect 21913 5859 21971 5865
rect 22002 5828 22008 5840
rect 18380 5800 20208 5828
rect 21560 5800 22008 5828
rect 18380 5788 18386 5800
rect 11940 5732 13216 5760
rect 11940 5720 11946 5732
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9217 5695 9275 5701
rect 9217 5661 9229 5695
rect 9263 5661 9275 5695
rect 9217 5655 9275 5661
rect 6512 5596 7052 5624
rect 7193 5627 7251 5633
rect 6512 5584 6518 5596
rect 7193 5593 7205 5627
rect 7239 5624 7251 5627
rect 7834 5624 7840 5636
rect 7239 5596 7840 5624
rect 7239 5593 7251 5596
rect 7193 5587 7251 5593
rect 7834 5584 7840 5596
rect 7892 5584 7898 5636
rect 9048 5624 9076 5655
rect 9490 5652 9496 5704
rect 9548 5652 9554 5704
rect 10226 5652 10232 5704
rect 10284 5692 10290 5704
rect 10689 5695 10747 5701
rect 10689 5692 10701 5695
rect 10284 5664 10701 5692
rect 10284 5652 10290 5664
rect 10689 5661 10701 5664
rect 10735 5661 10747 5695
rect 10689 5655 10747 5661
rect 10781 5695 10839 5701
rect 10781 5661 10793 5695
rect 10827 5661 10839 5695
rect 10781 5655 10839 5661
rect 9508 5624 9536 5652
rect 9048 5596 9536 5624
rect 10594 5584 10600 5636
rect 10652 5624 10658 5636
rect 10796 5624 10824 5655
rect 10870 5652 10876 5704
rect 10928 5652 10934 5704
rect 11606 5692 11612 5704
rect 11567 5664 11612 5692
rect 11606 5652 11612 5664
rect 11664 5652 11670 5704
rect 11701 5695 11759 5701
rect 11701 5661 11713 5695
rect 11747 5692 11759 5695
rect 11974 5692 11980 5704
rect 11747 5664 11980 5692
rect 11747 5661 11759 5664
rect 11701 5655 11759 5661
rect 11974 5652 11980 5664
rect 12032 5652 12038 5704
rect 12437 5695 12495 5701
rect 12437 5661 12449 5695
rect 12483 5661 12495 5695
rect 12437 5655 12495 5661
rect 12529 5695 12587 5701
rect 12529 5661 12541 5695
rect 12575 5692 12587 5695
rect 12618 5692 12624 5704
rect 12575 5664 12624 5692
rect 12575 5661 12587 5664
rect 12529 5655 12587 5661
rect 10652 5596 10824 5624
rect 12452 5624 12480 5655
rect 12618 5652 12624 5664
rect 12676 5652 12682 5704
rect 13188 5701 13216 5732
rect 13464 5732 15056 5760
rect 15136 5732 15516 5760
rect 12805 5695 12863 5701
rect 12805 5661 12817 5695
rect 12851 5692 12863 5695
rect 13173 5695 13231 5701
rect 12851 5664 13124 5692
rect 12851 5661 12863 5664
rect 12805 5655 12863 5661
rect 12710 5624 12716 5636
rect 12452 5596 12716 5624
rect 10652 5584 10658 5596
rect 12710 5584 12716 5596
rect 12768 5584 12774 5636
rect 12897 5627 12955 5633
rect 12897 5593 12909 5627
rect 12943 5624 12955 5627
rect 12986 5624 12992 5636
rect 12943 5596 12992 5624
rect 12943 5593 12955 5596
rect 12897 5587 12955 5593
rect 12986 5584 12992 5596
rect 13044 5584 13050 5636
rect 13096 5624 13124 5664
rect 13173 5661 13185 5695
rect 13219 5661 13231 5695
rect 13173 5655 13231 5661
rect 13354 5652 13360 5704
rect 13412 5652 13418 5704
rect 13464 5624 13492 5732
rect 13541 5695 13599 5701
rect 13541 5661 13553 5695
rect 13587 5692 13599 5695
rect 13722 5692 13728 5704
rect 13587 5664 13728 5692
rect 13587 5661 13599 5664
rect 13541 5655 13599 5661
rect 13722 5652 13728 5664
rect 13780 5652 13786 5704
rect 14274 5652 14280 5704
rect 14332 5692 14338 5704
rect 15043 5695 15101 5701
rect 15043 5692 15055 5695
rect 14332 5664 15055 5692
rect 14332 5652 14338 5664
rect 15043 5661 15055 5664
rect 15089 5692 15101 5695
rect 15136 5692 15164 5732
rect 15488 5701 15516 5732
rect 15746 5720 15752 5772
rect 15804 5720 15810 5772
rect 17310 5720 17316 5772
rect 17368 5760 17374 5772
rect 20070 5760 20076 5772
rect 17368 5732 20076 5760
rect 17368 5720 17374 5732
rect 20070 5720 20076 5732
rect 20128 5720 20134 5772
rect 21266 5760 21272 5772
rect 20180 5732 21272 5760
rect 15089 5664 15164 5692
rect 15197 5695 15255 5701
rect 15089 5661 15101 5664
rect 15043 5655 15101 5661
rect 15197 5661 15209 5695
rect 15243 5661 15255 5695
rect 15197 5655 15255 5661
rect 15473 5695 15531 5701
rect 15473 5661 15485 5695
rect 15519 5661 15531 5695
rect 15473 5655 15531 5661
rect 16393 5695 16451 5701
rect 16393 5661 16405 5695
rect 16439 5692 16451 5695
rect 16574 5692 16580 5704
rect 16439 5664 16580 5692
rect 16439 5661 16451 5664
rect 16393 5655 16451 5661
rect 13096 5596 13492 5624
rect 14369 5627 14427 5633
rect 14369 5593 14381 5627
rect 14415 5593 14427 5627
rect 15212 5624 15240 5655
rect 16408 5624 16436 5655
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 18230 5652 18236 5704
rect 18288 5652 18294 5704
rect 18969 5695 19027 5701
rect 18969 5661 18981 5695
rect 19015 5692 19027 5695
rect 19242 5692 19248 5704
rect 19015 5664 19248 5692
rect 19015 5661 19027 5664
rect 18969 5655 19027 5661
rect 19242 5652 19248 5664
rect 19300 5652 19306 5704
rect 19521 5695 19579 5701
rect 19521 5661 19533 5695
rect 19567 5692 19579 5695
rect 19794 5692 19800 5704
rect 19567 5664 19800 5692
rect 19567 5661 19579 5664
rect 19521 5655 19579 5661
rect 19794 5652 19800 5664
rect 19852 5692 19858 5704
rect 20180 5692 20208 5732
rect 21266 5720 21272 5732
rect 21324 5720 21330 5772
rect 21361 5763 21419 5769
rect 21361 5729 21373 5763
rect 21407 5760 21419 5763
rect 21560 5760 21588 5800
rect 22002 5788 22008 5800
rect 22060 5788 22066 5840
rect 21407 5732 21588 5760
rect 21637 5763 21695 5769
rect 21407 5729 21419 5732
rect 21361 5723 21419 5729
rect 21637 5729 21649 5763
rect 21683 5760 21695 5763
rect 21910 5760 21916 5772
rect 21683 5732 21916 5760
rect 21683 5729 21695 5732
rect 21637 5723 21695 5729
rect 21910 5720 21916 5732
rect 21968 5760 21974 5772
rect 22370 5760 22376 5772
rect 21968 5732 22376 5760
rect 21968 5720 21974 5732
rect 22370 5720 22376 5732
rect 22428 5720 22434 5772
rect 23014 5720 23020 5772
rect 23072 5760 23078 5772
rect 24121 5763 24179 5769
rect 24121 5760 24133 5763
rect 23072 5732 24133 5760
rect 23072 5720 23078 5732
rect 24121 5729 24133 5732
rect 24167 5729 24179 5763
rect 24121 5723 24179 5729
rect 19852 5664 20208 5692
rect 22097 5695 22155 5701
rect 19852 5652 19858 5664
rect 22097 5661 22109 5695
rect 22143 5692 22155 5695
rect 22278 5692 22284 5704
rect 22143 5664 22284 5692
rect 22143 5661 22155 5664
rect 22097 5655 22155 5661
rect 22278 5652 22284 5664
rect 22336 5652 22342 5704
rect 15212 5596 16436 5624
rect 14369 5587 14427 5593
rect 1780 5528 4292 5556
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 4801 5559 4859 5565
rect 4801 5556 4813 5559
rect 4672 5528 4813 5556
rect 4672 5516 4678 5528
rect 4801 5525 4813 5528
rect 4847 5525 4859 5559
rect 4801 5519 4859 5525
rect 6089 5559 6147 5565
rect 6089 5525 6101 5559
rect 6135 5556 6147 5559
rect 7374 5556 7380 5568
rect 6135 5528 7380 5556
rect 6135 5525 6147 5528
rect 6089 5519 6147 5525
rect 7374 5516 7380 5528
rect 7432 5516 7438 5568
rect 9217 5559 9275 5565
rect 9217 5525 9229 5559
rect 9263 5556 9275 5559
rect 9582 5556 9588 5568
rect 9263 5528 9588 5556
rect 9263 5525 9275 5528
rect 9217 5519 9275 5525
rect 9582 5516 9588 5528
rect 9640 5516 9646 5568
rect 10045 5559 10103 5565
rect 10045 5525 10057 5559
rect 10091 5556 10103 5559
rect 10778 5556 10784 5568
rect 10091 5528 10784 5556
rect 10091 5525 10103 5528
rect 10045 5519 10103 5525
rect 10778 5516 10784 5528
rect 10836 5516 10842 5568
rect 10962 5516 10968 5568
rect 11020 5556 11026 5568
rect 11057 5559 11115 5565
rect 11057 5556 11069 5559
rect 11020 5528 11069 5556
rect 11020 5516 11026 5528
rect 11057 5525 11069 5528
rect 11103 5525 11115 5559
rect 11057 5519 11115 5525
rect 11333 5559 11391 5565
rect 11333 5525 11345 5559
rect 11379 5556 11391 5559
rect 11698 5556 11704 5568
rect 11379 5528 11704 5556
rect 11379 5525 11391 5528
rect 11333 5519 11391 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 12802 5516 12808 5568
rect 12860 5556 12866 5568
rect 13170 5556 13176 5568
rect 12860 5528 13176 5556
rect 12860 5516 12866 5528
rect 13170 5516 13176 5528
rect 13228 5556 13234 5568
rect 14384 5556 14412 5587
rect 16666 5584 16672 5636
rect 16724 5584 16730 5636
rect 16942 5633 16948 5636
rect 16885 5627 16948 5633
rect 16885 5593 16897 5627
rect 16931 5593 16948 5627
rect 16885 5587 16948 5593
rect 16942 5584 16948 5587
rect 17000 5584 17006 5636
rect 17402 5584 17408 5636
rect 17460 5624 17466 5636
rect 17589 5627 17647 5633
rect 17589 5624 17601 5627
rect 17460 5596 17601 5624
rect 17460 5584 17466 5596
rect 17589 5593 17601 5596
rect 17635 5593 17647 5627
rect 17589 5587 17647 5593
rect 18432 5596 20116 5624
rect 13228 5528 14412 5556
rect 13228 5516 13234 5528
rect 14826 5516 14832 5568
rect 14884 5516 14890 5568
rect 17034 5516 17040 5568
rect 17092 5516 17098 5568
rect 17218 5516 17224 5568
rect 17276 5556 17282 5568
rect 17789 5559 17847 5565
rect 17789 5556 17801 5559
rect 17276 5528 17801 5556
rect 17276 5516 17282 5528
rect 17789 5525 17801 5528
rect 17835 5525 17847 5559
rect 17789 5519 17847 5525
rect 17954 5516 17960 5568
rect 18012 5516 18018 5568
rect 18432 5565 18460 5596
rect 18417 5559 18475 5565
rect 18417 5525 18429 5559
rect 18463 5525 18475 5559
rect 18417 5519 18475 5525
rect 18877 5559 18935 5565
rect 18877 5525 18889 5559
rect 18923 5556 18935 5559
rect 19150 5556 19156 5568
rect 18923 5528 19156 5556
rect 18923 5525 18935 5528
rect 18877 5519 18935 5525
rect 19150 5516 19156 5528
rect 19208 5516 19214 5568
rect 20088 5556 20116 5596
rect 20898 5584 20904 5636
rect 20956 5584 20962 5636
rect 22646 5584 22652 5636
rect 22704 5584 22710 5636
rect 23658 5584 23664 5636
rect 23716 5584 23722 5636
rect 21082 5556 21088 5568
rect 20088 5528 21088 5556
rect 21082 5516 21088 5528
rect 21140 5556 21146 5568
rect 21358 5556 21364 5568
rect 21140 5528 21364 5556
rect 21140 5516 21146 5528
rect 21358 5516 21364 5528
rect 21416 5556 21422 5568
rect 24670 5556 24676 5568
rect 21416 5528 24676 5556
rect 21416 5516 21422 5528
rect 24670 5516 24676 5528
rect 24728 5516 24734 5568
rect 1104 5466 24840 5488
rect 1104 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 24214 5466
rect 24266 5414 24278 5466
rect 24330 5414 24342 5466
rect 24394 5414 24406 5466
rect 24458 5414 24470 5466
rect 24522 5414 24840 5466
rect 1104 5392 24840 5414
rect 2222 5312 2228 5364
rect 2280 5352 2286 5364
rect 4157 5355 4215 5361
rect 4157 5352 4169 5355
rect 2280 5324 4169 5352
rect 2280 5312 2286 5324
rect 4157 5321 4169 5324
rect 4203 5321 4215 5355
rect 4157 5315 4215 5321
rect 1670 5244 1676 5296
rect 1728 5244 1734 5296
rect 4172 5284 4200 5315
rect 7282 5312 7288 5364
rect 7340 5312 7346 5364
rect 7374 5312 7380 5364
rect 7432 5352 7438 5364
rect 7926 5352 7932 5364
rect 7432 5324 7932 5352
rect 7432 5312 7438 5324
rect 7926 5312 7932 5324
rect 7984 5312 7990 5364
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5321 8815 5355
rect 8757 5315 8815 5321
rect 5534 5284 5540 5296
rect 4172 5256 5028 5284
rect 2406 5176 2412 5228
rect 2464 5216 2470 5228
rect 2593 5219 2651 5225
rect 2593 5216 2605 5219
rect 2464 5188 2605 5216
rect 2464 5176 2470 5188
rect 2593 5185 2605 5188
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 3050 5176 3056 5228
rect 3108 5176 3114 5228
rect 3605 5219 3663 5225
rect 3605 5185 3617 5219
rect 3651 5185 3663 5219
rect 3605 5179 3663 5185
rect 3620 5148 3648 5179
rect 3970 5176 3976 5228
rect 4028 5216 4034 5228
rect 4065 5219 4123 5225
rect 4065 5216 4077 5219
rect 4028 5188 4077 5216
rect 4028 5176 4034 5188
rect 4065 5185 4077 5188
rect 4111 5185 4123 5219
rect 4065 5179 4123 5185
rect 4341 5219 4399 5225
rect 4341 5185 4353 5219
rect 4387 5216 4399 5219
rect 4890 5216 4896 5228
rect 4387 5188 4896 5216
rect 4387 5185 4399 5188
rect 4341 5179 4399 5185
rect 4890 5176 4896 5188
rect 4948 5176 4954 5228
rect 4614 5148 4620 5160
rect 3620 5120 4620 5148
rect 4614 5108 4620 5120
rect 4672 5108 4678 5160
rect 4798 5108 4804 5160
rect 4856 5108 4862 5160
rect 5000 5148 5028 5256
rect 5184 5256 5540 5284
rect 5184 5225 5212 5256
rect 5534 5244 5540 5256
rect 5592 5284 5598 5296
rect 6454 5284 6460 5296
rect 5592 5256 6460 5284
rect 5592 5244 5598 5256
rect 6454 5244 6460 5256
rect 6512 5244 6518 5296
rect 8772 5284 8800 5315
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 12345 5355 12403 5361
rect 10376 5324 10916 5352
rect 10376 5312 10382 5324
rect 9490 5284 9496 5296
rect 8772 5256 9496 5284
rect 9490 5244 9496 5256
rect 9548 5284 9554 5296
rect 9548 5256 10732 5284
rect 9548 5244 9554 5256
rect 10704 5228 10732 5256
rect 5169 5219 5227 5225
rect 5169 5185 5181 5219
rect 5215 5185 5227 5219
rect 5721 5219 5779 5225
rect 5721 5216 5733 5219
rect 5169 5179 5227 5185
rect 5276 5188 5733 5216
rect 5276 5148 5304 5188
rect 5721 5185 5733 5188
rect 5767 5216 5779 5219
rect 6270 5216 6276 5228
rect 5767 5188 6276 5216
rect 5767 5185 5779 5188
rect 5721 5179 5779 5185
rect 6270 5176 6276 5188
rect 6328 5176 6334 5228
rect 7006 5176 7012 5228
rect 7064 5176 7070 5228
rect 7101 5219 7159 5225
rect 7101 5185 7113 5219
rect 7147 5216 7159 5219
rect 7558 5216 7564 5228
rect 7147 5188 7564 5216
rect 7147 5185 7159 5188
rect 7101 5179 7159 5185
rect 7558 5176 7564 5188
rect 7616 5176 7622 5228
rect 7834 5176 7840 5228
rect 7892 5176 7898 5228
rect 8205 5219 8263 5225
rect 8205 5185 8217 5219
rect 8251 5185 8263 5219
rect 8205 5179 8263 5185
rect 5000 5120 5304 5148
rect 5537 5151 5595 5157
rect 5537 5117 5549 5151
rect 5583 5148 5595 5151
rect 6178 5148 6184 5160
rect 5583 5120 6184 5148
rect 5583 5117 5595 5120
rect 5537 5111 5595 5117
rect 6178 5108 6184 5120
rect 6236 5108 6242 5160
rect 7469 5151 7527 5157
rect 7469 5117 7481 5151
rect 7515 5148 7527 5151
rect 8110 5148 8116 5160
rect 7515 5120 8116 5148
rect 7515 5117 7527 5120
rect 7469 5111 7527 5117
rect 2038 5040 2044 5092
rect 2096 5040 2102 5092
rect 2314 5040 2320 5092
rect 2372 5080 2378 5092
rect 6089 5083 6147 5089
rect 2372 5052 3556 5080
rect 2372 5040 2378 5052
rect 3528 5024 3556 5052
rect 6089 5049 6101 5083
rect 6135 5080 6147 5083
rect 7484 5080 7512 5111
rect 8110 5108 8116 5120
rect 8168 5148 8174 5160
rect 8220 5148 8248 5179
rect 8662 5176 8668 5228
rect 8720 5176 8726 5228
rect 10226 5176 10232 5228
rect 10284 5176 10290 5228
rect 10410 5176 10416 5228
rect 10468 5176 10474 5228
rect 10686 5176 10692 5228
rect 10744 5176 10750 5228
rect 10888 5225 10916 5324
rect 12345 5321 12357 5355
rect 12391 5352 12403 5355
rect 12618 5352 12624 5364
rect 12391 5324 12624 5352
rect 12391 5321 12403 5324
rect 12345 5315 12403 5321
rect 12618 5312 12624 5324
rect 12676 5312 12682 5364
rect 12710 5312 12716 5364
rect 12768 5352 12774 5364
rect 15102 5352 15108 5364
rect 12768 5324 15108 5352
rect 12768 5312 12774 5324
rect 15102 5312 15108 5324
rect 15160 5312 15166 5364
rect 15381 5355 15439 5361
rect 15381 5321 15393 5355
rect 15427 5352 15439 5355
rect 15562 5352 15568 5364
rect 15427 5324 15568 5352
rect 15427 5321 15439 5324
rect 15381 5315 15439 5321
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 15856 5324 18644 5352
rect 11606 5244 11612 5296
rect 11664 5284 11670 5296
rect 14277 5287 14335 5293
rect 11664 5256 12112 5284
rect 11664 5244 11670 5256
rect 10873 5219 10931 5225
rect 10873 5185 10885 5219
rect 10919 5185 10931 5219
rect 11974 5216 11980 5228
rect 11935 5188 11980 5216
rect 10873 5179 10931 5185
rect 11974 5176 11980 5188
rect 12032 5176 12038 5228
rect 12084 5225 12112 5256
rect 12406 5256 13952 5284
rect 12069 5219 12127 5225
rect 12069 5185 12081 5219
rect 12115 5185 12127 5219
rect 12069 5179 12127 5185
rect 8168 5120 8248 5148
rect 8168 5108 8174 5120
rect 9122 5108 9128 5160
rect 9180 5148 9186 5160
rect 9674 5148 9680 5160
rect 9180 5120 9680 5148
rect 9180 5108 9186 5120
rect 9674 5108 9680 5120
rect 9732 5108 9738 5160
rect 10597 5151 10655 5157
rect 10597 5117 10609 5151
rect 10643 5148 10655 5151
rect 12406 5148 12434 5256
rect 12544 5225 12572 5256
rect 12529 5219 12587 5225
rect 12529 5185 12541 5219
rect 12575 5185 12587 5219
rect 12529 5179 12587 5185
rect 13538 5176 13544 5228
rect 13596 5176 13602 5228
rect 13725 5219 13783 5225
rect 13725 5185 13737 5219
rect 13771 5185 13783 5219
rect 13725 5179 13783 5185
rect 10643 5120 12434 5148
rect 12621 5151 12679 5157
rect 10643 5117 10655 5120
rect 10597 5111 10655 5117
rect 12621 5117 12633 5151
rect 12667 5117 12679 5151
rect 12621 5111 12679 5117
rect 6135 5052 7512 5080
rect 11701 5083 11759 5089
rect 6135 5049 6147 5052
rect 6089 5043 6147 5049
rect 11701 5049 11713 5083
rect 11747 5049 11759 5083
rect 11701 5043 11759 5049
rect 2133 5015 2191 5021
rect 2133 4981 2145 5015
rect 2179 5012 2191 5015
rect 3326 5012 3332 5024
rect 2179 4984 3332 5012
rect 2179 4981 2191 4984
rect 2133 4975 2191 4981
rect 3326 4972 3332 4984
rect 3384 4972 3390 5024
rect 3510 4972 3516 5024
rect 3568 4972 3574 5024
rect 4341 5015 4399 5021
rect 4341 4981 4353 5015
rect 4387 5012 4399 5015
rect 5258 5012 5264 5024
rect 4387 4984 5264 5012
rect 4387 4981 4399 4984
rect 4341 4975 4399 4981
rect 5258 4972 5264 4984
rect 5316 4972 5322 5024
rect 6454 4972 6460 5024
rect 6512 4972 6518 5024
rect 6825 5015 6883 5021
rect 6825 4981 6837 5015
rect 6871 5012 6883 5015
rect 7006 5012 7012 5024
rect 6871 4984 7012 5012
rect 6871 4981 6883 4984
rect 6825 4975 6883 4981
rect 7006 4972 7012 4984
rect 7064 4972 7070 5024
rect 7374 4972 7380 5024
rect 7432 5012 7438 5024
rect 9217 5015 9275 5021
rect 9217 5012 9229 5015
rect 7432 4984 9229 5012
rect 7432 4972 7438 4984
rect 9217 4981 9229 4984
rect 9263 4981 9275 5015
rect 11716 5012 11744 5043
rect 11882 5040 11888 5092
rect 11940 5080 11946 5092
rect 12636 5080 12664 5111
rect 12710 5108 12716 5160
rect 12768 5108 12774 5160
rect 12802 5108 12808 5160
rect 12860 5108 12866 5160
rect 13446 5108 13452 5160
rect 13504 5148 13510 5160
rect 13740 5148 13768 5179
rect 13814 5176 13820 5228
rect 13872 5176 13878 5228
rect 13924 5216 13952 5256
rect 14277 5253 14289 5287
rect 14323 5284 14335 5287
rect 14366 5284 14372 5296
rect 14323 5256 14372 5284
rect 14323 5253 14335 5256
rect 14277 5247 14335 5253
rect 14366 5244 14372 5256
rect 14424 5244 14430 5296
rect 14461 5287 14519 5293
rect 14461 5253 14473 5287
rect 14507 5284 14519 5287
rect 14826 5284 14832 5296
rect 14507 5256 14832 5284
rect 14507 5253 14519 5256
rect 14461 5247 14519 5253
rect 14826 5244 14832 5256
rect 14884 5244 14890 5296
rect 14553 5219 14611 5225
rect 13924 5188 14504 5216
rect 13504 5120 14412 5148
rect 13504 5108 13510 5120
rect 13725 5083 13783 5089
rect 13725 5080 13737 5083
rect 11940 5052 13737 5080
rect 11940 5040 11946 5052
rect 13725 5049 13737 5052
rect 13771 5080 13783 5083
rect 13906 5080 13912 5092
rect 13771 5052 13912 5080
rect 13771 5049 13783 5052
rect 13725 5043 13783 5049
rect 13906 5040 13912 5052
rect 13964 5040 13970 5092
rect 14384 5089 14412 5120
rect 14369 5083 14427 5089
rect 14369 5049 14381 5083
rect 14415 5049 14427 5083
rect 14476 5080 14504 5188
rect 14553 5185 14565 5219
rect 14599 5216 14611 5219
rect 14599 5188 14688 5216
rect 14599 5185 14611 5188
rect 14553 5179 14611 5185
rect 14660 5148 14688 5188
rect 15010 5176 15016 5228
rect 15068 5216 15074 5228
rect 15856 5225 15884 5324
rect 17954 5244 17960 5296
rect 18012 5244 18018 5296
rect 18616 5284 18644 5324
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 19058 5352 19064 5364
rect 18748 5324 19064 5352
rect 18748 5312 18754 5324
rect 19058 5312 19064 5324
rect 19116 5312 19122 5364
rect 19168 5324 20668 5352
rect 19168 5284 19196 5324
rect 18616 5256 19196 5284
rect 19245 5287 19303 5293
rect 19245 5253 19257 5287
rect 19291 5284 19303 5287
rect 19518 5284 19524 5296
rect 19291 5256 19524 5284
rect 19291 5253 19303 5256
rect 19245 5247 19303 5253
rect 19518 5244 19524 5256
rect 19576 5244 19582 5296
rect 19702 5244 19708 5296
rect 19760 5244 19766 5296
rect 15381 5219 15439 5225
rect 15381 5216 15393 5219
rect 15068 5188 15393 5216
rect 15068 5176 15074 5188
rect 15381 5185 15393 5188
rect 15427 5185 15439 5219
rect 15381 5179 15439 5185
rect 15841 5219 15899 5225
rect 15841 5185 15853 5219
rect 15887 5185 15899 5219
rect 15841 5179 15899 5185
rect 15933 5219 15991 5225
rect 15933 5185 15945 5219
rect 15979 5216 15991 5219
rect 16850 5216 16856 5228
rect 15979 5188 16856 5216
rect 15979 5185 15991 5188
rect 15933 5179 15991 5185
rect 16850 5176 16856 5188
rect 16908 5176 16914 5228
rect 14734 5148 14740 5160
rect 14660 5120 14740 5148
rect 14734 5108 14740 5120
rect 14792 5148 14798 5160
rect 15473 5151 15531 5157
rect 15473 5148 15485 5151
rect 14792 5120 15485 5148
rect 14792 5108 14798 5120
rect 15473 5117 15485 5120
rect 15519 5148 15531 5151
rect 15746 5148 15752 5160
rect 15519 5120 15752 5148
rect 15519 5117 15531 5120
rect 15473 5111 15531 5117
rect 15746 5108 15752 5120
rect 15804 5108 15810 5160
rect 16114 5108 16120 5160
rect 16172 5108 16178 5160
rect 16758 5108 16764 5160
rect 16816 5148 16822 5160
rect 16945 5151 17003 5157
rect 16945 5148 16957 5151
rect 16816 5120 16957 5148
rect 16816 5108 16822 5120
rect 16945 5117 16957 5120
rect 16991 5117 17003 5151
rect 16945 5111 17003 5117
rect 17221 5151 17279 5157
rect 17221 5117 17233 5151
rect 17267 5148 17279 5151
rect 17310 5148 17316 5160
rect 17267 5120 17316 5148
rect 17267 5117 17279 5120
rect 17221 5111 17279 5117
rect 15378 5080 15384 5092
rect 14476 5052 15384 5080
rect 14369 5043 14427 5049
rect 15378 5040 15384 5052
rect 15436 5040 15442 5092
rect 16574 5080 16580 5092
rect 15488 5052 16580 5080
rect 11974 5012 11980 5024
rect 11716 4984 11980 5012
rect 9217 4975 9275 4981
rect 11974 4972 11980 4984
rect 12032 4972 12038 5024
rect 12802 4972 12808 5024
rect 12860 5012 12866 5024
rect 15488 5012 15516 5052
rect 16574 5040 16580 5052
rect 16632 5040 16638 5092
rect 12860 4984 15516 5012
rect 16025 5015 16083 5021
rect 12860 4972 12866 4984
rect 16025 4981 16037 5015
rect 16071 5012 16083 5015
rect 16666 5012 16672 5024
rect 16071 4984 16672 5012
rect 16071 4981 16083 4984
rect 16025 4975 16083 4981
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 16960 5012 16988 5111
rect 17310 5108 17316 5120
rect 17368 5108 17374 5160
rect 18969 5151 19027 5157
rect 18969 5117 18981 5151
rect 19015 5148 19027 5151
rect 19978 5148 19984 5160
rect 19015 5120 19984 5148
rect 19015 5117 19027 5120
rect 18969 5111 19027 5117
rect 18984 5012 19012 5111
rect 19978 5108 19984 5120
rect 20036 5108 20042 5160
rect 20640 5148 20668 5324
rect 20714 5312 20720 5364
rect 20772 5312 20778 5364
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 20993 5355 21051 5361
rect 20993 5352 21005 5355
rect 20956 5324 21005 5352
rect 20956 5312 20962 5324
rect 20993 5321 21005 5324
rect 21039 5321 21051 5355
rect 20993 5315 21051 5321
rect 21161 5355 21219 5361
rect 21161 5321 21173 5355
rect 21207 5352 21219 5355
rect 21542 5352 21548 5364
rect 21207 5324 21548 5352
rect 21207 5321 21219 5324
rect 21161 5315 21219 5321
rect 21542 5312 21548 5324
rect 21600 5352 21606 5364
rect 21600 5324 22416 5352
rect 21600 5312 21606 5324
rect 20732 5284 20760 5312
rect 20732 5256 21036 5284
rect 21008 5228 21036 5256
rect 21358 5244 21364 5296
rect 21416 5284 21422 5296
rect 22388 5293 22416 5324
rect 22646 5312 22652 5364
rect 22704 5352 22710 5364
rect 22833 5355 22891 5361
rect 22833 5352 22845 5355
rect 22704 5324 22845 5352
rect 22704 5312 22710 5324
rect 22833 5321 22845 5324
rect 22879 5321 22891 5355
rect 22833 5315 22891 5321
rect 23014 5312 23020 5364
rect 23072 5352 23078 5364
rect 23201 5355 23259 5361
rect 23201 5352 23213 5355
rect 23072 5324 23213 5352
rect 23072 5312 23078 5324
rect 23201 5321 23213 5324
rect 23247 5321 23259 5355
rect 23201 5315 23259 5321
rect 23290 5312 23296 5364
rect 23348 5312 23354 5364
rect 23934 5312 23940 5364
rect 23992 5352 23998 5364
rect 24029 5355 24087 5361
rect 24029 5352 24041 5355
rect 23992 5324 24041 5352
rect 23992 5312 23998 5324
rect 24029 5321 24041 5324
rect 24075 5321 24087 5355
rect 24029 5315 24087 5321
rect 22189 5287 22247 5293
rect 22189 5284 22201 5287
rect 21416 5256 22201 5284
rect 21416 5244 21422 5256
rect 22189 5253 22201 5256
rect 22235 5253 22247 5287
rect 22388 5287 22463 5293
rect 22388 5256 22417 5287
rect 22189 5247 22247 5253
rect 22405 5253 22417 5256
rect 22451 5284 22463 5287
rect 24181 5287 24239 5293
rect 24181 5284 24193 5287
rect 22451 5256 24193 5284
rect 22451 5253 22463 5256
rect 22405 5247 22463 5253
rect 24181 5253 24193 5256
rect 24227 5253 24239 5287
rect 24181 5247 24239 5253
rect 24397 5287 24455 5293
rect 24397 5253 24409 5287
rect 24443 5253 24455 5287
rect 24397 5247 24455 5253
rect 20990 5176 20996 5228
rect 21048 5176 21054 5228
rect 21726 5176 21732 5228
rect 21784 5216 21790 5228
rect 24412 5216 24440 5247
rect 21784 5188 22094 5216
rect 21784 5176 21790 5188
rect 21358 5148 21364 5160
rect 20640 5120 21364 5148
rect 21358 5108 21364 5120
rect 21416 5108 21422 5160
rect 22066 5148 22094 5188
rect 23308 5188 24440 5216
rect 23308 5148 23336 5188
rect 22066 5120 23336 5148
rect 23382 5108 23388 5160
rect 23440 5108 23446 5160
rect 22388 5052 24256 5080
rect 16960 4984 19012 5012
rect 20714 4972 20720 5024
rect 20772 5012 20778 5024
rect 21174 5012 21180 5024
rect 20772 4984 21180 5012
rect 20772 4972 20778 4984
rect 21174 4972 21180 4984
rect 21232 5012 21238 5024
rect 22388 5021 22416 5052
rect 22373 5015 22431 5021
rect 22373 5012 22385 5015
rect 21232 4984 22385 5012
rect 21232 4972 21238 4984
rect 22373 4981 22385 4984
rect 22419 4981 22431 5015
rect 22373 4975 22431 4981
rect 22557 5015 22615 5021
rect 22557 4981 22569 5015
rect 22603 5012 22615 5015
rect 22738 5012 22744 5024
rect 22603 4984 22744 5012
rect 22603 4981 22615 4984
rect 22557 4975 22615 4981
rect 22738 4972 22744 4984
rect 22796 4972 22802 5024
rect 24228 5021 24256 5052
rect 24213 5015 24271 5021
rect 24213 4981 24225 5015
rect 24259 4981 24271 5015
rect 24213 4975 24271 4981
rect 1104 4922 24840 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 20214 4922
rect 20266 4870 20278 4922
rect 20330 4870 20342 4922
rect 20394 4870 20406 4922
rect 20458 4870 20470 4922
rect 20522 4870 24840 4922
rect 1104 4848 24840 4870
rect 1394 4768 1400 4820
rect 1452 4808 1458 4820
rect 1489 4811 1547 4817
rect 1489 4808 1501 4811
rect 1452 4780 1501 4808
rect 1452 4768 1458 4780
rect 1489 4777 1501 4780
rect 1535 4777 1547 4811
rect 1489 4771 1547 4777
rect 2038 4768 2044 4820
rect 2096 4808 2102 4820
rect 2593 4811 2651 4817
rect 2593 4808 2605 4811
rect 2096 4780 2605 4808
rect 2096 4768 2102 4780
rect 2593 4777 2605 4780
rect 2639 4777 2651 4811
rect 2593 4771 2651 4777
rect 2682 4768 2688 4820
rect 2740 4808 2746 4820
rect 2740 4780 2901 4808
rect 2740 4768 2746 4780
rect 1854 4700 1860 4752
rect 1912 4700 1918 4752
rect 2774 4740 2780 4752
rect 2056 4712 2780 4740
rect 2056 4613 2084 4712
rect 2774 4700 2780 4712
rect 2832 4700 2838 4752
rect 2873 4681 2901 4780
rect 4890 4768 4896 4820
rect 4948 4808 4954 4820
rect 5169 4811 5227 4817
rect 5169 4808 5181 4811
rect 4948 4780 5181 4808
rect 4948 4768 4954 4780
rect 5169 4777 5181 4780
rect 5215 4777 5227 4811
rect 5169 4771 5227 4777
rect 5184 4740 5212 4771
rect 7282 4768 7288 4820
rect 7340 4808 7346 4820
rect 8754 4808 8760 4820
rect 7340 4780 8760 4808
rect 7340 4768 7346 4780
rect 8754 4768 8760 4780
rect 8812 4768 8818 4820
rect 9861 4811 9919 4817
rect 9861 4808 9873 4811
rect 9232 4780 9873 4808
rect 5184 4712 6132 4740
rect 2869 4675 2927 4681
rect 2869 4641 2881 4675
rect 2915 4641 2927 4675
rect 2869 4635 2927 4641
rect 2958 4632 2964 4684
rect 3016 4632 3022 4684
rect 3053 4675 3111 4681
rect 3053 4641 3065 4675
rect 3099 4672 3111 4675
rect 4062 4672 4068 4684
rect 3099 4644 4068 4672
rect 3099 4641 3111 4644
rect 3053 4635 3111 4641
rect 4062 4632 4068 4644
rect 4120 4632 4126 4684
rect 5353 4675 5411 4681
rect 5353 4641 5365 4675
rect 5399 4672 5411 4675
rect 5534 4672 5540 4684
rect 5399 4644 5540 4672
rect 5399 4641 5411 4644
rect 5353 4635 5411 4641
rect 5534 4632 5540 4644
rect 5592 4632 5598 4684
rect 6104 4681 6132 4712
rect 6089 4675 6147 4681
rect 6089 4641 6101 4675
rect 6135 4641 6147 4675
rect 6089 4635 6147 4641
rect 6178 4632 6184 4684
rect 6236 4632 6242 4684
rect 6270 4632 6276 4684
rect 6328 4632 6334 4684
rect 6917 4675 6975 4681
rect 6917 4641 6929 4675
rect 6963 4672 6975 4675
rect 7190 4672 7196 4684
rect 6963 4644 7196 4672
rect 6963 4641 6975 4644
rect 6917 4635 6975 4641
rect 7190 4632 7196 4644
rect 7248 4632 7254 4684
rect 7374 4632 7380 4684
rect 7432 4632 7438 4684
rect 8389 4675 8447 4681
rect 8389 4641 8401 4675
rect 8435 4672 8447 4675
rect 9122 4672 9128 4684
rect 8435 4644 9128 4672
rect 8435 4641 8447 4644
rect 8389 4635 8447 4641
rect 9122 4632 9128 4644
rect 9180 4632 9186 4684
rect 2041 4607 2099 4613
rect 2041 4573 2053 4607
rect 2087 4573 2099 4607
rect 2041 4567 2099 4573
rect 2314 4564 2320 4616
rect 2372 4564 2378 4616
rect 2777 4607 2835 4613
rect 2777 4573 2789 4607
rect 2823 4604 2835 4607
rect 3234 4604 3240 4616
rect 2823 4576 3240 4604
rect 2823 4573 2835 4576
rect 2777 4567 2835 4573
rect 2222 4428 2228 4480
rect 2280 4428 2286 4480
rect 2498 4428 2504 4480
rect 2556 4468 2562 4480
rect 2792 4468 2820 4567
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3510 4564 3516 4616
rect 3568 4604 3574 4616
rect 3881 4607 3939 4613
rect 3881 4604 3893 4607
rect 3568 4576 3893 4604
rect 3568 4564 3574 4576
rect 3881 4573 3893 4576
rect 3927 4573 3939 4607
rect 3881 4567 3939 4573
rect 3970 4564 3976 4616
rect 4028 4604 4034 4616
rect 4249 4607 4307 4613
rect 4249 4604 4261 4607
rect 4028 4576 4261 4604
rect 4028 4564 4034 4576
rect 4249 4573 4261 4576
rect 4295 4573 4307 4607
rect 4249 4567 4307 4573
rect 4264 4536 4292 4567
rect 4614 4564 4620 4616
rect 4672 4564 4678 4616
rect 4798 4564 4804 4616
rect 4856 4604 4862 4616
rect 5442 4604 5448 4616
rect 4856 4576 5448 4604
rect 4856 4564 4862 4576
rect 5442 4564 5448 4576
rect 5500 4564 5506 4616
rect 6196 4536 6224 4632
rect 6365 4607 6423 4613
rect 6365 4573 6377 4607
rect 6411 4573 6423 4607
rect 6365 4567 6423 4573
rect 4264 4508 6224 4536
rect 6380 4536 6408 4567
rect 7006 4564 7012 4616
rect 7064 4564 7070 4616
rect 7098 4564 7104 4616
rect 7156 4604 7162 4616
rect 7285 4607 7343 4613
rect 7285 4604 7297 4607
rect 7156 4576 7297 4604
rect 7156 4564 7162 4576
rect 7285 4573 7297 4576
rect 7331 4604 7343 4607
rect 7650 4604 7656 4616
rect 7331 4576 7656 4604
rect 7331 4573 7343 4576
rect 7285 4567 7343 4573
rect 7650 4564 7656 4576
rect 7708 4564 7714 4616
rect 8662 4564 8668 4616
rect 8720 4564 8726 4616
rect 9232 4613 9260 4780
rect 9861 4777 9873 4780
rect 9907 4808 9919 4811
rect 10870 4808 10876 4820
rect 9907 4780 10876 4808
rect 9907 4777 9919 4780
rect 9861 4771 9919 4777
rect 10870 4768 10876 4780
rect 10928 4768 10934 4820
rect 12710 4768 12716 4820
rect 12768 4808 12774 4820
rect 13081 4811 13139 4817
rect 13081 4808 13093 4811
rect 12768 4780 13093 4808
rect 12768 4768 12774 4780
rect 13081 4777 13093 4780
rect 13127 4777 13139 4811
rect 13081 4771 13139 4777
rect 13814 4768 13820 4820
rect 13872 4808 13878 4820
rect 15473 4811 15531 4817
rect 15473 4808 15485 4811
rect 13872 4780 15485 4808
rect 13872 4768 13878 4780
rect 15473 4777 15485 4780
rect 15519 4777 15531 4811
rect 15473 4771 15531 4777
rect 17310 4768 17316 4820
rect 17368 4768 17374 4820
rect 19521 4811 19579 4817
rect 19521 4777 19533 4811
rect 19567 4777 19579 4811
rect 19521 4771 19579 4777
rect 11698 4740 11704 4752
rect 9784 4712 11704 4740
rect 9033 4607 9091 4613
rect 9033 4573 9045 4607
rect 9079 4573 9091 4607
rect 9033 4567 9091 4573
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4573 9275 4607
rect 9674 4604 9680 4616
rect 9217 4567 9275 4573
rect 9508 4576 9680 4604
rect 7116 4536 7144 4564
rect 6380 4508 7144 4536
rect 9048 4536 9076 4567
rect 9508 4536 9536 4576
rect 9674 4564 9680 4576
rect 9732 4564 9738 4616
rect 9784 4613 9812 4712
rect 11698 4700 11704 4712
rect 11756 4700 11762 4752
rect 12618 4700 12624 4752
rect 12676 4700 12682 4752
rect 14274 4700 14280 4752
rect 14332 4740 14338 4752
rect 15010 4740 15016 4752
rect 14332 4712 15016 4740
rect 14332 4700 14338 4712
rect 15010 4700 15016 4712
rect 15068 4700 15074 4752
rect 15102 4700 15108 4752
rect 15160 4740 15166 4752
rect 15197 4743 15255 4749
rect 15197 4740 15209 4743
rect 15160 4712 15209 4740
rect 15160 4700 15166 4712
rect 15197 4709 15209 4712
rect 15243 4709 15255 4743
rect 18417 4743 18475 4749
rect 18417 4740 18429 4743
rect 15197 4703 15255 4709
rect 16776 4712 18429 4740
rect 11974 4672 11980 4684
rect 9876 4644 11980 4672
rect 9876 4613 9904 4644
rect 9769 4607 9827 4613
rect 9769 4573 9781 4607
rect 9815 4573 9827 4607
rect 9769 4567 9827 4573
rect 9861 4607 9919 4613
rect 9861 4573 9873 4607
rect 9907 4573 9919 4607
rect 9861 4567 9919 4573
rect 10229 4607 10287 4613
rect 10229 4573 10241 4607
rect 10275 4604 10287 4607
rect 10318 4604 10324 4616
rect 10275 4576 10324 4604
rect 10275 4573 10287 4576
rect 10229 4567 10287 4573
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 10505 4607 10563 4613
rect 10505 4573 10517 4607
rect 10551 4604 10563 4607
rect 10686 4604 10692 4616
rect 10551 4576 10692 4604
rect 10551 4573 10563 4576
rect 10505 4567 10563 4573
rect 10686 4564 10692 4576
rect 10744 4564 10750 4616
rect 10781 4607 10839 4613
rect 10781 4573 10793 4607
rect 10827 4573 10839 4607
rect 10781 4567 10839 4573
rect 9048 4508 9536 4536
rect 9585 4539 9643 4545
rect 9585 4505 9597 4539
rect 9631 4536 9643 4539
rect 9950 4536 9956 4548
rect 9631 4508 9956 4536
rect 9631 4505 9643 4508
rect 9585 4499 9643 4505
rect 9950 4496 9956 4508
rect 10008 4496 10014 4548
rect 10042 4496 10048 4548
rect 10100 4536 10106 4548
rect 10100 4508 10732 4536
rect 10100 4496 10106 4508
rect 10704 4480 10732 4508
rect 2556 4440 2820 4468
rect 2556 4428 2562 4440
rect 2866 4428 2872 4480
rect 2924 4468 2930 4480
rect 3421 4471 3479 4477
rect 3421 4468 3433 4471
rect 2924 4440 3433 4468
rect 2924 4428 2930 4440
rect 3421 4437 3433 4440
rect 3467 4437 3479 4471
rect 3421 4431 3479 4437
rect 5350 4428 5356 4480
rect 5408 4468 5414 4480
rect 5905 4471 5963 4477
rect 5905 4468 5917 4471
rect 5408 4440 5917 4468
rect 5408 4428 5414 4440
rect 5905 4437 5917 4440
rect 5951 4437 5963 4471
rect 5905 4431 5963 4437
rect 6733 4471 6791 4477
rect 6733 4437 6745 4471
rect 6779 4468 6791 4471
rect 6822 4468 6828 4480
rect 6779 4440 6828 4468
rect 6779 4437 6791 4440
rect 6733 4431 6791 4437
rect 6822 4428 6828 4440
rect 6880 4428 6886 4480
rect 9217 4471 9275 4477
rect 9217 4437 9229 4471
rect 9263 4468 9275 4471
rect 10410 4468 10416 4480
rect 9263 4440 10416 4468
rect 9263 4437 9275 4440
rect 9217 4431 9275 4437
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10686 4428 10692 4480
rect 10744 4428 10750 4480
rect 10796 4468 10824 4567
rect 10962 4564 10968 4616
rect 11020 4564 11026 4616
rect 11422 4564 11428 4616
rect 11480 4564 11486 4616
rect 11624 4613 11652 4644
rect 11974 4632 11980 4644
rect 12032 4672 12038 4684
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 12032 4644 13303 4672
rect 12032 4632 12038 4644
rect 11609 4607 11667 4613
rect 11609 4573 11621 4607
rect 11655 4573 11667 4607
rect 11609 4567 11667 4573
rect 11698 4564 11704 4616
rect 11756 4564 11762 4616
rect 12529 4607 12587 4613
rect 12529 4573 12541 4607
rect 12575 4604 12587 4607
rect 12713 4607 12771 4613
rect 12575 4576 12664 4604
rect 12575 4573 12587 4576
rect 12529 4567 12587 4573
rect 10870 4496 10876 4548
rect 10928 4496 10934 4548
rect 11882 4536 11888 4548
rect 10980 4508 11888 4536
rect 10980 4468 11008 4508
rect 11882 4496 11888 4508
rect 11940 4496 11946 4548
rect 12636 4536 12664 4576
rect 12713 4573 12725 4607
rect 12759 4604 12771 4607
rect 12802 4604 12808 4616
rect 12759 4576 12808 4604
rect 12759 4573 12771 4576
rect 12713 4567 12771 4573
rect 12802 4564 12808 4576
rect 12860 4564 12866 4616
rect 13275 4613 13303 4644
rect 13592 4644 14197 4672
rect 13592 4616 13620 4644
rect 14185 4641 14197 4644
rect 14231 4641 14243 4675
rect 14185 4635 14243 4641
rect 14458 4632 14464 4684
rect 14516 4672 14522 4684
rect 14516 4644 15608 4672
rect 14516 4632 14522 4644
rect 13260 4607 13318 4613
rect 13260 4573 13272 4607
rect 13306 4573 13318 4607
rect 13260 4567 13318 4573
rect 12894 4536 12900 4548
rect 12636 4508 12900 4536
rect 12894 4496 12900 4508
rect 12952 4496 12958 4548
rect 13275 4536 13303 4567
rect 13354 4564 13360 4616
rect 13412 4564 13418 4616
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 13538 4564 13544 4616
rect 13596 4613 13620 4616
rect 13596 4607 13635 4613
rect 13623 4573 13635 4607
rect 13596 4567 13635 4573
rect 13596 4564 13602 4567
rect 13722 4564 13728 4616
rect 13780 4604 13786 4616
rect 14274 4604 14280 4616
rect 13780 4576 14280 4604
rect 13780 4564 13786 4576
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14366 4564 14372 4616
rect 14424 4564 14430 4616
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14645 4607 14703 4613
rect 14645 4573 14657 4607
rect 14691 4604 14703 4607
rect 14826 4604 14832 4616
rect 14691 4576 14832 4604
rect 14691 4573 14703 4576
rect 14645 4567 14703 4573
rect 14826 4564 14832 4576
rect 14884 4564 14890 4616
rect 14918 4564 14924 4616
rect 14976 4564 14982 4616
rect 15010 4564 15016 4616
rect 15068 4604 15074 4616
rect 15473 4607 15531 4613
rect 15473 4604 15485 4607
rect 15068 4576 15485 4604
rect 15068 4564 15074 4576
rect 15473 4573 15485 4576
rect 15519 4573 15531 4607
rect 15580 4604 15608 4644
rect 15654 4632 15660 4684
rect 15712 4672 15718 4684
rect 16776 4681 16804 4712
rect 18417 4709 18429 4712
rect 18463 4709 18475 4743
rect 19536 4740 19564 4771
rect 19702 4768 19708 4820
rect 19760 4768 19766 4820
rect 20714 4808 20720 4820
rect 19812 4780 20720 4808
rect 19812 4740 19840 4780
rect 20714 4768 20720 4780
rect 20772 4768 20778 4820
rect 22370 4768 22376 4820
rect 22428 4808 22434 4820
rect 23014 4808 23020 4820
rect 22428 4780 23020 4808
rect 22428 4768 22434 4780
rect 23014 4768 23020 4780
rect 23072 4808 23078 4820
rect 23750 4808 23756 4820
rect 23072 4780 23756 4808
rect 23072 4768 23078 4780
rect 23750 4768 23756 4780
rect 23808 4768 23814 4820
rect 24118 4768 24124 4820
rect 24176 4768 24182 4820
rect 19536 4712 19840 4740
rect 18417 4703 18475 4709
rect 16761 4675 16819 4681
rect 16761 4672 16773 4675
rect 15712 4644 16773 4672
rect 15712 4632 15718 4644
rect 16761 4641 16773 4644
rect 16807 4641 16819 4675
rect 16761 4635 16819 4641
rect 17494 4632 17500 4684
rect 17552 4672 17558 4684
rect 17865 4675 17923 4681
rect 17865 4672 17877 4675
rect 17552 4644 17877 4672
rect 17552 4632 17558 4644
rect 17865 4641 17877 4644
rect 17911 4672 17923 4675
rect 19610 4672 19616 4684
rect 17911 4644 19616 4672
rect 17911 4641 17923 4644
rect 17865 4635 17923 4641
rect 19610 4632 19616 4644
rect 19668 4632 19674 4684
rect 19812 4616 19840 4712
rect 21542 4672 21548 4684
rect 19904 4644 21548 4672
rect 15749 4607 15807 4613
rect 15749 4604 15761 4607
rect 15580 4576 15761 4604
rect 15473 4567 15531 4573
rect 15749 4573 15761 4576
rect 15795 4573 15807 4607
rect 15749 4567 15807 4573
rect 17681 4607 17739 4613
rect 17681 4573 17693 4607
rect 17727 4604 17739 4607
rect 18690 4604 18696 4616
rect 17727 4576 18696 4604
rect 17727 4573 17739 4576
rect 17681 4567 17739 4573
rect 15197 4539 15255 4545
rect 13275 4508 15148 4536
rect 10796 4440 11008 4468
rect 11238 4428 11244 4480
rect 11296 4428 11302 4480
rect 11698 4428 11704 4480
rect 11756 4468 11762 4480
rect 11977 4471 12035 4477
rect 11977 4468 11989 4471
rect 11756 4440 11989 4468
rect 11756 4428 11762 4440
rect 11977 4437 11989 4440
rect 12023 4437 12035 4471
rect 11977 4431 12035 4437
rect 13814 4428 13820 4480
rect 13872 4468 13878 4480
rect 15013 4471 15071 4477
rect 15013 4468 15025 4471
rect 13872 4440 15025 4468
rect 13872 4428 13878 4440
rect 15013 4437 15025 4440
rect 15059 4437 15071 4471
rect 15120 4468 15148 4508
rect 15197 4505 15209 4539
rect 15243 4536 15255 4539
rect 15378 4536 15384 4548
rect 15243 4508 15384 4536
rect 15243 4505 15255 4508
rect 15197 4499 15255 4505
rect 15378 4496 15384 4508
rect 15436 4496 15442 4548
rect 15764 4536 15792 4567
rect 18690 4564 18696 4576
rect 18748 4564 18754 4616
rect 18874 4564 18880 4616
rect 18932 4564 18938 4616
rect 19794 4564 19800 4616
rect 19852 4564 19858 4616
rect 17773 4539 17831 4545
rect 17773 4536 17785 4539
rect 15764 4508 17785 4536
rect 17773 4505 17785 4508
rect 17819 4505 17831 4539
rect 19334 4536 19340 4548
rect 17773 4499 17831 4505
rect 19306 4496 19340 4536
rect 19392 4496 19398 4548
rect 19610 4545 19616 4548
rect 19553 4539 19616 4545
rect 19553 4505 19565 4539
rect 19599 4505 19616 4539
rect 19553 4499 19616 4505
rect 19610 4496 19616 4499
rect 19668 4536 19674 4548
rect 19904 4536 19932 4644
rect 21542 4632 21548 4644
rect 21600 4632 21606 4684
rect 23198 4632 23204 4684
rect 23256 4632 23262 4684
rect 19978 4564 19984 4616
rect 20036 4564 20042 4616
rect 20257 4539 20315 4545
rect 20257 4536 20269 4539
rect 19668 4508 19932 4536
rect 20088 4508 20269 4536
rect 19668 4496 19674 4508
rect 15657 4471 15715 4477
rect 15657 4468 15669 4471
rect 15120 4440 15669 4468
rect 15013 4431 15071 4437
rect 15657 4437 15669 4440
rect 15703 4437 15715 4471
rect 15657 4431 15715 4437
rect 15838 4428 15844 4480
rect 15896 4468 15902 4480
rect 16301 4471 16359 4477
rect 16301 4468 16313 4471
rect 15896 4440 16313 4468
rect 15896 4428 15902 4440
rect 16301 4437 16313 4440
rect 16347 4437 16359 4471
rect 16301 4431 16359 4437
rect 17586 4428 17592 4480
rect 17644 4468 17650 4480
rect 19306 4468 19334 4496
rect 20088 4480 20116 4508
rect 20257 4505 20269 4508
rect 20303 4505 20315 4539
rect 20257 4499 20315 4505
rect 20714 4496 20720 4548
rect 20772 4496 20778 4548
rect 22094 4496 22100 4548
rect 22152 4496 22158 4548
rect 17644 4440 19334 4468
rect 17644 4428 17650 4440
rect 20070 4428 20076 4480
rect 20128 4428 20134 4480
rect 21726 4428 21732 4480
rect 21784 4428 21790 4480
rect 23290 4428 23296 4480
rect 23348 4428 23354 4480
rect 23382 4428 23388 4480
rect 23440 4428 23446 4480
rect 23753 4471 23811 4477
rect 23753 4437 23765 4471
rect 23799 4468 23811 4471
rect 23934 4468 23940 4480
rect 23799 4440 23940 4468
rect 23799 4437 23811 4440
rect 23753 4431 23811 4437
rect 23934 4428 23940 4440
rect 23992 4428 23998 4480
rect 1104 4378 24840 4400
rect 1104 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 24214 4378
rect 24266 4326 24278 4378
rect 24330 4326 24342 4378
rect 24394 4326 24406 4378
rect 24458 4326 24470 4378
rect 24522 4326 24840 4378
rect 1104 4304 24840 4326
rect 2774 4224 2780 4276
rect 2832 4264 2838 4276
rect 4157 4267 4215 4273
rect 4157 4264 4169 4267
rect 2832 4236 4169 4264
rect 2832 4224 2838 4236
rect 4157 4233 4169 4236
rect 4203 4264 4215 4267
rect 4614 4264 4620 4276
rect 4203 4236 4620 4264
rect 4203 4233 4215 4236
rect 4157 4227 4215 4233
rect 4614 4224 4620 4236
rect 4672 4224 4678 4276
rect 7098 4264 7104 4276
rect 5644 4236 7104 4264
rect 1949 4199 2007 4205
rect 1949 4165 1961 4199
rect 1995 4196 2007 4199
rect 2038 4196 2044 4208
rect 1995 4168 2044 4196
rect 1995 4165 2007 4168
rect 1949 4159 2007 4165
rect 2038 4156 2044 4168
rect 2096 4156 2102 4208
rect 2406 4156 2412 4208
rect 2464 4156 2470 4208
rect 5644 4205 5672 4236
rect 7098 4224 7104 4236
rect 7156 4224 7162 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 10594 4264 10600 4276
rect 9732 4236 10600 4264
rect 9732 4224 9738 4236
rect 10594 4224 10600 4236
rect 10652 4264 10658 4276
rect 11238 4264 11244 4276
rect 10652 4236 11244 4264
rect 10652 4224 10658 4236
rect 11238 4224 11244 4236
rect 11296 4224 11302 4276
rect 12529 4267 12587 4273
rect 12529 4233 12541 4267
rect 12575 4264 12587 4267
rect 13722 4264 13728 4276
rect 12575 4236 13728 4264
rect 12575 4233 12587 4236
rect 12529 4227 12587 4233
rect 13722 4224 13728 4236
rect 13780 4224 13786 4276
rect 13906 4264 13912 4276
rect 13832 4236 13912 4264
rect 5629 4199 5687 4205
rect 5629 4165 5641 4199
rect 5675 4165 5687 4199
rect 5629 4159 5687 4165
rect 3970 4088 3976 4140
rect 4028 4088 4034 4140
rect 4062 4088 4068 4140
rect 4120 4128 4126 4140
rect 4433 4131 4491 4137
rect 4433 4128 4445 4131
rect 4120 4100 4445 4128
rect 4120 4088 4126 4100
rect 4433 4097 4445 4100
rect 4479 4097 4491 4131
rect 4433 4091 4491 4097
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4128 4675 4131
rect 4890 4128 4896 4140
rect 4663 4100 4896 4128
rect 4663 4097 4675 4100
rect 4617 4091 4675 4097
rect 4890 4088 4896 4100
rect 4948 4088 4954 4140
rect 5258 4088 5264 4140
rect 5316 4088 5322 4140
rect 5350 4088 5356 4140
rect 5408 4088 5414 4140
rect 1486 4020 1492 4072
rect 1544 4060 1550 4072
rect 1673 4063 1731 4069
rect 1673 4060 1685 4063
rect 1544 4032 1685 4060
rect 1544 4020 1550 4032
rect 1673 4029 1685 4032
rect 1719 4029 1731 4063
rect 1673 4023 1731 4029
rect 1688 3924 1716 4023
rect 3142 4020 3148 4072
rect 3200 4060 3206 4072
rect 3697 4063 3755 4069
rect 3697 4060 3709 4063
rect 3200 4032 3709 4060
rect 3200 4020 3206 4032
rect 3697 4029 3709 4032
rect 3743 4060 3755 4063
rect 4706 4060 4712 4072
rect 3743 4032 4712 4060
rect 3743 4029 3755 4032
rect 3697 4023 3755 4029
rect 4706 4020 4712 4032
rect 4764 4020 4770 4072
rect 4801 4063 4859 4069
rect 4801 4029 4813 4063
rect 4847 4060 4859 4063
rect 5644 4060 5672 4159
rect 6822 4156 6828 4208
rect 6880 4196 6886 4208
rect 6917 4199 6975 4205
rect 6917 4196 6929 4199
rect 6880 4168 6929 4196
rect 6880 4156 6886 4168
rect 6917 4165 6929 4168
rect 6963 4165 6975 4199
rect 6917 4159 6975 4165
rect 7374 4156 7380 4208
rect 7432 4156 7438 4208
rect 9582 4156 9588 4208
rect 9640 4196 9646 4208
rect 9640 4168 10180 4196
rect 9640 4156 9646 4168
rect 9217 4131 9275 4137
rect 9217 4097 9229 4131
rect 9263 4128 9275 4131
rect 9306 4128 9312 4140
rect 9263 4100 9312 4128
rect 9263 4097 9275 4100
rect 9217 4091 9275 4097
rect 9306 4088 9312 4100
rect 9364 4088 9370 4140
rect 9401 4131 9459 4137
rect 9401 4097 9413 4131
rect 9447 4128 9459 4131
rect 9766 4128 9772 4140
rect 9447 4100 9772 4128
rect 9447 4097 9459 4100
rect 9401 4091 9459 4097
rect 9766 4088 9772 4100
rect 9824 4088 9830 4140
rect 9861 4131 9919 4137
rect 9861 4097 9873 4131
rect 9907 4097 9919 4131
rect 9861 4091 9919 4097
rect 4847 4032 5672 4060
rect 5721 4063 5779 4069
rect 4847 4029 4859 4032
rect 4801 4023 4859 4029
rect 5721 4029 5733 4063
rect 5767 4060 5779 4063
rect 5994 4060 6000 4072
rect 5767 4032 6000 4060
rect 5767 4029 5779 4032
rect 5721 4023 5779 4029
rect 5994 4020 6000 4032
rect 6052 4020 6058 4072
rect 6641 4063 6699 4069
rect 6641 4029 6653 4063
rect 6687 4029 6699 4063
rect 6641 4023 6699 4029
rect 3326 3952 3332 4004
rect 3384 3992 3390 4004
rect 3789 3995 3847 4001
rect 3789 3992 3801 3995
rect 3384 3964 3801 3992
rect 3384 3952 3390 3964
rect 3789 3961 3801 3964
rect 3835 3961 3847 3995
rect 3789 3955 3847 3961
rect 3234 3924 3240 3936
rect 1688 3896 3240 3924
rect 3234 3884 3240 3896
rect 3292 3884 3298 3936
rect 3421 3927 3479 3933
rect 3421 3893 3433 3927
rect 3467 3924 3479 3927
rect 4890 3924 4896 3936
rect 3467 3896 4896 3924
rect 3467 3893 3479 3896
rect 3421 3887 3479 3893
rect 4890 3884 4896 3896
rect 4948 3884 4954 3936
rect 5077 3927 5135 3933
rect 5077 3893 5089 3927
rect 5123 3924 5135 3927
rect 5166 3924 5172 3936
rect 5123 3896 5172 3924
rect 5123 3893 5135 3896
rect 5077 3887 5135 3893
rect 5166 3884 5172 3896
rect 5224 3884 5230 3936
rect 6089 3927 6147 3933
rect 6089 3893 6101 3927
rect 6135 3924 6147 3927
rect 6546 3924 6552 3936
rect 6135 3896 6552 3924
rect 6135 3893 6147 3896
rect 6089 3887 6147 3893
rect 6546 3884 6552 3896
rect 6604 3884 6610 3936
rect 6656 3924 6684 4023
rect 7006 4020 7012 4072
rect 7064 4060 7070 4072
rect 7466 4060 7472 4072
rect 7064 4032 7472 4060
rect 7064 4020 7070 4032
rect 7466 4020 7472 4032
rect 7524 4020 7530 4072
rect 7650 4020 7656 4072
rect 7708 4060 7714 4072
rect 9674 4060 9680 4072
rect 7708 4032 9680 4060
rect 7708 4020 7714 4032
rect 9674 4020 9680 4032
rect 9732 4060 9738 4072
rect 9876 4060 9904 4091
rect 9950 4088 9956 4140
rect 10008 4088 10014 4140
rect 10045 4131 10103 4137
rect 10045 4097 10057 4131
rect 10091 4097 10103 4131
rect 10152 4128 10180 4168
rect 10318 4156 10324 4208
rect 10376 4196 10382 4208
rect 10376 4168 10824 4196
rect 10376 4156 10382 4168
rect 10612 4140 10640 4168
rect 10229 4131 10287 4137
rect 10229 4128 10241 4131
rect 10152 4100 10241 4128
rect 10045 4091 10103 4097
rect 10229 4097 10241 4100
rect 10275 4097 10287 4131
rect 10229 4091 10287 4097
rect 9732 4032 9904 4060
rect 10060 4060 10088 4091
rect 10594 4088 10600 4140
rect 10652 4088 10658 4140
rect 10686 4088 10692 4140
rect 10744 4088 10750 4140
rect 10796 4128 10824 4168
rect 10870 4156 10876 4208
rect 10928 4196 10934 4208
rect 13832 4196 13860 4236
rect 13906 4224 13912 4236
rect 13964 4264 13970 4276
rect 14918 4264 14924 4276
rect 13964 4236 14924 4264
rect 13964 4224 13970 4236
rect 14918 4224 14924 4236
rect 14976 4224 14982 4276
rect 15930 4264 15936 4276
rect 15488 4236 15936 4264
rect 10928 4168 13308 4196
rect 10928 4156 10934 4168
rect 10965 4131 11023 4137
rect 10965 4128 10977 4131
rect 10796 4100 10977 4128
rect 10965 4097 10977 4100
rect 11011 4097 11023 4131
rect 10965 4091 11023 4097
rect 11609 4131 11667 4137
rect 11609 4097 11621 4131
rect 11655 4097 11667 4131
rect 11609 4091 11667 4097
rect 11793 4131 11851 4137
rect 11793 4097 11805 4131
rect 11839 4128 11851 4131
rect 11974 4128 11980 4140
rect 11839 4100 11980 4128
rect 11839 4097 11851 4100
rect 11793 4091 11851 4097
rect 10505 4063 10563 4069
rect 10505 4060 10517 4063
rect 10060 4032 10517 4060
rect 9732 4020 9738 4032
rect 10505 4029 10517 4032
rect 10551 4029 10563 4063
rect 10505 4023 10563 4029
rect 10778 4020 10784 4072
rect 10836 4060 10842 4072
rect 10873 4063 10931 4069
rect 10873 4060 10885 4063
rect 10836 4032 10885 4060
rect 10836 4020 10842 4032
rect 10873 4029 10885 4032
rect 10919 4029 10931 4063
rect 11624 4060 11652 4091
rect 11974 4088 11980 4100
rect 12032 4088 12038 4140
rect 12710 4088 12716 4140
rect 12768 4128 12774 4140
rect 13173 4131 13231 4137
rect 13173 4128 13185 4131
rect 12768 4100 13185 4128
rect 12768 4088 12774 4100
rect 13173 4097 13185 4100
rect 13219 4097 13231 4131
rect 13173 4091 13231 4097
rect 11882 4060 11888 4072
rect 11624 4032 11888 4060
rect 10873 4023 10931 4029
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 12066 4020 12072 4072
rect 12124 4020 12130 4072
rect 12802 4060 12808 4072
rect 12360 4032 12808 4060
rect 8754 3992 8760 4004
rect 7944 3964 8760 3992
rect 7098 3924 7104 3936
rect 6656 3896 7104 3924
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 7466 3884 7472 3936
rect 7524 3924 7530 3936
rect 7944 3924 7972 3964
rect 8754 3952 8760 3964
rect 8812 3952 8818 4004
rect 9309 3995 9367 4001
rect 9309 3961 9321 3995
rect 9355 3992 9367 3995
rect 12360 3992 12388 4032
rect 12802 4020 12808 4032
rect 12860 4020 12866 4072
rect 9355 3964 12388 3992
rect 12437 3995 12495 4001
rect 9355 3961 9367 3964
rect 9309 3955 9367 3961
rect 12437 3961 12449 3995
rect 12483 3992 12495 3995
rect 12710 3992 12716 4004
rect 12483 3964 12716 3992
rect 12483 3961 12495 3964
rect 12437 3955 12495 3961
rect 12710 3952 12716 3964
rect 12768 3952 12774 4004
rect 13188 3992 13216 4091
rect 13280 4060 13308 4168
rect 13464 4168 13860 4196
rect 14476 4168 14688 4196
rect 13357 4131 13415 4137
rect 13357 4097 13369 4131
rect 13403 4128 13415 4131
rect 13464 4128 13492 4168
rect 13403 4100 13492 4128
rect 13403 4097 13415 4100
rect 13357 4091 13415 4097
rect 13538 4088 13544 4140
rect 13596 4128 13602 4140
rect 14476 4137 14504 4168
rect 13817 4131 13875 4137
rect 13817 4128 13829 4131
rect 13596 4100 13829 4128
rect 13596 4088 13602 4100
rect 13817 4097 13829 4100
rect 13863 4097 13875 4131
rect 13817 4091 13875 4097
rect 14461 4131 14519 4137
rect 14461 4097 14473 4131
rect 14507 4097 14519 4131
rect 14461 4091 14519 4097
rect 14553 4131 14611 4137
rect 14553 4097 14565 4131
rect 14599 4097 14611 4131
rect 14553 4091 14611 4097
rect 14568 4060 14596 4091
rect 13280 4032 14596 4060
rect 14660 4060 14688 4168
rect 15010 4088 15016 4140
rect 15068 4128 15074 4140
rect 15488 4128 15516 4236
rect 15930 4224 15936 4236
rect 15988 4224 15994 4276
rect 16114 4224 16120 4276
rect 16172 4224 16178 4276
rect 17678 4224 17684 4276
rect 17736 4264 17742 4276
rect 19219 4267 19277 4273
rect 19219 4264 19231 4267
rect 17736 4236 19231 4264
rect 17736 4224 17742 4236
rect 15562 4156 15568 4208
rect 15620 4196 15626 4208
rect 15620 4168 16344 4196
rect 15620 4156 15626 4168
rect 15068 4100 15516 4128
rect 15068 4088 15074 4100
rect 15654 4088 15660 4140
rect 15712 4088 15718 4140
rect 16316 4137 16344 4168
rect 17034 4156 17040 4208
rect 17092 4196 17098 4208
rect 18785 4199 18843 4205
rect 17092 4168 17526 4196
rect 17092 4156 17098 4168
rect 18785 4165 18797 4199
rect 18831 4196 18843 4199
rect 18874 4196 18880 4208
rect 18831 4168 18880 4196
rect 18831 4165 18843 4168
rect 18785 4159 18843 4165
rect 16301 4131 16359 4137
rect 16301 4097 16313 4131
rect 16347 4097 16359 4131
rect 16301 4091 16359 4097
rect 16393 4131 16451 4137
rect 16393 4097 16405 4131
rect 16439 4097 16451 4131
rect 16393 4091 16451 4097
rect 15289 4063 15347 4069
rect 15289 4060 15301 4063
rect 14660 4032 15301 4060
rect 15289 4029 15301 4032
rect 15335 4060 15347 4063
rect 15470 4060 15476 4072
rect 15335 4032 15476 4060
rect 15335 4029 15347 4032
rect 15289 4023 15347 4029
rect 15470 4020 15476 4032
rect 15528 4020 15534 4072
rect 15562 4020 15568 4072
rect 15620 4020 15626 4072
rect 16117 4063 16175 4069
rect 16117 4060 16129 4063
rect 15764 4032 16129 4060
rect 13630 3992 13636 4004
rect 13188 3964 13636 3992
rect 13630 3952 13636 3964
rect 13688 3952 13694 4004
rect 15194 3992 15200 4004
rect 13832 3964 15200 3992
rect 7524 3896 7972 3924
rect 8389 3927 8447 3933
rect 7524 3884 7530 3896
rect 8389 3893 8401 3927
rect 8435 3924 8447 3927
rect 8662 3924 8668 3936
rect 8435 3896 8668 3924
rect 8435 3893 8447 3896
rect 8389 3887 8447 3893
rect 8662 3884 8668 3896
rect 8720 3884 8726 3936
rect 9674 3884 9680 3936
rect 9732 3884 9738 3936
rect 11701 3927 11759 3933
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 11882 3924 11888 3936
rect 11747 3896 11888 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12897 3927 12955 3933
rect 12897 3893 12909 3927
rect 12943 3924 12955 3927
rect 13446 3924 13452 3936
rect 12943 3896 13452 3924
rect 12943 3893 12955 3896
rect 12897 3887 12955 3893
rect 13446 3884 13452 3896
rect 13504 3884 13510 3936
rect 13541 3927 13599 3933
rect 13541 3893 13553 3927
rect 13587 3924 13599 3927
rect 13832 3924 13860 3964
rect 15194 3952 15200 3964
rect 15252 3952 15258 4004
rect 15764 3936 15792 4032
rect 16117 4029 16129 4032
rect 16163 4029 16175 4063
rect 16117 4023 16175 4029
rect 13587 3896 13860 3924
rect 13909 3927 13967 3933
rect 13587 3893 13599 3896
rect 13541 3887 13599 3893
rect 13909 3893 13921 3927
rect 13955 3924 13967 3927
rect 14182 3924 14188 3936
rect 13955 3896 14188 3924
rect 13955 3893 13967 3896
rect 13909 3887 13967 3893
rect 14182 3884 14188 3896
rect 14240 3924 14246 3936
rect 15746 3924 15752 3936
rect 14240 3896 15752 3924
rect 14240 3884 14246 3896
rect 15746 3884 15752 3896
rect 15804 3884 15810 3936
rect 16114 3884 16120 3936
rect 16172 3924 16178 3936
rect 16408 3924 16436 4091
rect 16758 4020 16764 4072
rect 16816 4020 16822 4072
rect 17034 4020 17040 4072
rect 17092 4020 17098 4072
rect 18800 4060 18828 4159
rect 18874 4156 18880 4168
rect 18932 4156 18938 4208
rect 18064 4032 18828 4060
rect 18064 3924 18092 4032
rect 18874 4020 18880 4072
rect 18932 4060 18938 4072
rect 18968 4060 18996 4236
rect 19219 4233 19231 4236
rect 19265 4264 19277 4267
rect 19610 4264 19616 4276
rect 19265 4236 19616 4264
rect 19265 4233 19277 4236
rect 19219 4227 19277 4233
rect 19610 4224 19616 4236
rect 19668 4264 19674 4276
rect 19905 4267 19963 4273
rect 19905 4264 19917 4267
rect 19668 4236 19917 4264
rect 19668 4224 19674 4236
rect 19905 4233 19917 4236
rect 19951 4233 19963 4267
rect 19905 4227 19963 4233
rect 20070 4224 20076 4276
rect 20128 4264 20134 4276
rect 20349 4267 20407 4273
rect 20349 4264 20361 4267
rect 20128 4236 20361 4264
rect 20128 4224 20134 4236
rect 20349 4233 20361 4236
rect 20395 4233 20407 4267
rect 20349 4227 20407 4233
rect 20809 4267 20867 4273
rect 20809 4233 20821 4267
rect 20855 4264 20867 4267
rect 20990 4264 20996 4276
rect 20855 4236 20996 4264
rect 20855 4233 20867 4236
rect 20809 4227 20867 4233
rect 20990 4224 20996 4236
rect 21048 4224 21054 4276
rect 21542 4224 21548 4276
rect 21600 4224 21606 4276
rect 23474 4264 23480 4276
rect 22204 4236 23480 4264
rect 19334 4156 19340 4208
rect 19392 4196 19398 4208
rect 19429 4199 19487 4205
rect 19429 4196 19441 4199
rect 19392 4168 19441 4196
rect 19392 4156 19398 4168
rect 19429 4165 19441 4168
rect 19475 4196 19487 4199
rect 19705 4199 19763 4205
rect 19705 4196 19717 4199
rect 19475 4168 19717 4196
rect 19475 4165 19487 4168
rect 19429 4159 19487 4165
rect 19705 4165 19717 4168
rect 19751 4165 19763 4199
rect 19705 4159 19763 4165
rect 20717 4199 20775 4205
rect 20717 4165 20729 4199
rect 20763 4196 20775 4199
rect 21726 4196 21732 4208
rect 20763 4168 21732 4196
rect 20763 4165 20775 4168
rect 20717 4159 20775 4165
rect 19720 4128 19748 4159
rect 21726 4156 21732 4168
rect 21784 4156 21790 4208
rect 20806 4128 20812 4140
rect 19720 4100 20812 4128
rect 20806 4088 20812 4100
rect 20864 4128 20870 4140
rect 21082 4128 21088 4140
rect 20864 4100 21088 4128
rect 20864 4088 20870 4100
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 21361 4131 21419 4137
rect 21361 4097 21373 4131
rect 21407 4128 21419 4131
rect 22204 4128 22232 4236
rect 23474 4224 23480 4236
rect 23532 4224 23538 4276
rect 24118 4196 24124 4208
rect 23690 4168 24124 4196
rect 24118 4156 24124 4168
rect 24176 4156 24182 4208
rect 21407 4100 22232 4128
rect 24397 4131 24455 4137
rect 21407 4097 21419 4100
rect 21361 4091 21419 4097
rect 24397 4097 24409 4131
rect 24443 4128 24455 4131
rect 24578 4128 24584 4140
rect 24443 4100 24584 4128
rect 24443 4097 24455 4100
rect 24397 4091 24455 4097
rect 24578 4088 24584 4100
rect 24636 4088 24642 4140
rect 18932 4032 18996 4060
rect 20993 4063 21051 4069
rect 18932 4020 18938 4032
rect 20993 4029 21005 4063
rect 21039 4060 21051 4063
rect 21174 4060 21180 4072
rect 21039 4032 21180 4060
rect 21039 4029 21051 4032
rect 20993 4023 21051 4029
rect 21174 4020 21180 4032
rect 21232 4060 21238 4072
rect 22002 4060 22008 4072
rect 21232 4032 22008 4060
rect 21232 4020 21238 4032
rect 22002 4020 22008 4032
rect 22060 4020 22066 4072
rect 22189 4063 22247 4069
rect 22189 4029 22201 4063
rect 22235 4029 22247 4063
rect 22189 4023 22247 4029
rect 22465 4063 22523 4069
rect 22465 4029 22477 4063
rect 22511 4060 22523 4063
rect 22554 4060 22560 4072
rect 22511 4032 22560 4060
rect 22511 4029 22523 4032
rect 22465 4023 22523 4029
rect 18966 3952 18972 4004
rect 19024 3992 19030 4004
rect 19024 3964 19288 3992
rect 19024 3952 19030 3964
rect 16172 3896 18092 3924
rect 16172 3884 16178 3896
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 19260 3933 19288 3964
rect 19978 3952 19984 4004
rect 20036 3992 20042 4004
rect 21910 3992 21916 4004
rect 20036 3964 21916 3992
rect 20036 3952 20042 3964
rect 21910 3952 21916 3964
rect 21968 3992 21974 4004
rect 22204 3992 22232 4023
rect 22554 4020 22560 4032
rect 22612 4020 22618 4072
rect 23198 4020 23204 4072
rect 23256 4060 23262 4072
rect 23937 4063 23995 4069
rect 23937 4060 23949 4063
rect 23256 4032 23949 4060
rect 23256 4020 23262 4032
rect 23937 4029 23949 4032
rect 23983 4029 23995 4063
rect 23937 4023 23995 4029
rect 21968 3964 22232 3992
rect 21968 3952 21974 3964
rect 19061 3927 19119 3933
rect 19061 3924 19073 3927
rect 18288 3896 19073 3924
rect 18288 3884 18294 3896
rect 19061 3893 19073 3896
rect 19107 3893 19119 3927
rect 19061 3887 19119 3893
rect 19245 3927 19303 3933
rect 19245 3893 19257 3927
rect 19291 3924 19303 3927
rect 19794 3924 19800 3936
rect 19291 3896 19800 3924
rect 19291 3893 19303 3896
rect 19245 3887 19303 3893
rect 19794 3884 19800 3896
rect 19852 3924 19858 3936
rect 19889 3927 19947 3933
rect 19889 3924 19901 3927
rect 19852 3896 19901 3924
rect 19852 3884 19858 3896
rect 19889 3893 19901 3896
rect 19935 3893 19947 3927
rect 19889 3887 19947 3893
rect 20073 3927 20131 3933
rect 20073 3893 20085 3927
rect 20119 3924 20131 3927
rect 20714 3924 20720 3936
rect 20119 3896 20720 3924
rect 20119 3893 20131 3896
rect 20073 3887 20131 3893
rect 20714 3884 20720 3896
rect 20772 3884 20778 3936
rect 22204 3924 22232 3964
rect 23842 3952 23848 4004
rect 23900 3992 23906 4004
rect 24213 3995 24271 4001
rect 24213 3992 24225 3995
rect 23900 3964 24225 3992
rect 23900 3952 23906 3964
rect 24213 3961 24225 3964
rect 24259 3961 24271 3995
rect 24213 3955 24271 3961
rect 23750 3924 23756 3936
rect 22204 3896 23756 3924
rect 23750 3884 23756 3896
rect 23808 3884 23814 3936
rect 1104 3834 24840 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 20214 3834
rect 20266 3782 20278 3834
rect 20330 3782 20342 3834
rect 20394 3782 20406 3834
rect 20458 3782 20470 3834
rect 20522 3782 24840 3834
rect 1104 3760 24840 3782
rect 2038 3680 2044 3732
rect 2096 3720 2102 3732
rect 2133 3723 2191 3729
rect 2133 3720 2145 3723
rect 2096 3692 2145 3720
rect 2096 3680 2102 3692
rect 2133 3689 2145 3692
rect 2179 3689 2191 3723
rect 2133 3683 2191 3689
rect 2317 3723 2375 3729
rect 2317 3689 2329 3723
rect 2363 3720 2375 3723
rect 2406 3720 2412 3732
rect 2363 3692 2412 3720
rect 2363 3689 2375 3692
rect 2317 3683 2375 3689
rect 2406 3680 2412 3692
rect 2464 3680 2470 3732
rect 2516 3692 6316 3720
rect 1673 3655 1731 3661
rect 1673 3621 1685 3655
rect 1719 3652 1731 3655
rect 2516 3652 2544 3692
rect 1719 3624 2544 3652
rect 1719 3621 1731 3624
rect 1673 3615 1731 3621
rect 2590 3612 2596 3664
rect 2648 3612 2654 3664
rect 3970 3652 3976 3664
rect 2884 3624 3976 3652
rect 2314 3544 2320 3596
rect 2372 3584 2378 3596
rect 2884 3593 2912 3624
rect 3970 3612 3976 3624
rect 4028 3612 4034 3664
rect 6288 3652 6316 3692
rect 6362 3680 6368 3732
rect 6420 3720 6426 3732
rect 7006 3720 7012 3732
rect 6420 3692 7012 3720
rect 6420 3680 6426 3692
rect 7006 3680 7012 3692
rect 7064 3720 7070 3732
rect 7193 3723 7251 3729
rect 7193 3720 7205 3723
rect 7064 3692 7205 3720
rect 7064 3680 7070 3692
rect 7193 3689 7205 3692
rect 7239 3689 7251 3723
rect 7193 3683 7251 3689
rect 7374 3680 7380 3732
rect 7432 3680 7438 3732
rect 9858 3720 9864 3732
rect 7484 3692 9864 3720
rect 7484 3652 7512 3692
rect 9858 3680 9864 3692
rect 9916 3680 9922 3732
rect 9950 3680 9956 3732
rect 10008 3720 10014 3732
rect 10410 3720 10416 3732
rect 10008 3692 10416 3720
rect 10008 3680 10014 3692
rect 10410 3680 10416 3692
rect 10468 3720 10474 3732
rect 10781 3723 10839 3729
rect 10781 3720 10793 3723
rect 10468 3692 10793 3720
rect 10468 3680 10474 3692
rect 10781 3689 10793 3692
rect 10827 3720 10839 3723
rect 11606 3720 11612 3732
rect 10827 3692 11612 3720
rect 10827 3689 10839 3692
rect 10781 3683 10839 3689
rect 11606 3680 11612 3692
rect 11664 3720 11670 3732
rect 12710 3720 12716 3732
rect 11664 3692 12716 3720
rect 11664 3680 11670 3692
rect 12710 3680 12716 3692
rect 12768 3680 12774 3732
rect 15390 3723 15448 3729
rect 15390 3689 15402 3723
rect 15436 3689 15448 3723
rect 15390 3683 15448 3689
rect 16393 3723 16451 3729
rect 16393 3689 16405 3723
rect 16439 3720 16451 3723
rect 17034 3720 17040 3732
rect 16439 3692 17040 3720
rect 16439 3689 16451 3692
rect 16393 3683 16451 3689
rect 6288 3624 7512 3652
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 7708 3624 8432 3652
rect 7708 3612 7714 3624
rect 2777 3587 2835 3593
rect 2777 3584 2789 3587
rect 2372 3556 2789 3584
rect 2372 3544 2378 3556
rect 2777 3553 2789 3556
rect 2823 3553 2835 3587
rect 2777 3547 2835 3553
rect 2869 3587 2927 3593
rect 2869 3553 2881 3587
rect 2915 3553 2927 3587
rect 2869 3547 2927 3553
rect 1394 3476 1400 3528
rect 1452 3516 1458 3528
rect 1489 3519 1547 3525
rect 1489 3516 1501 3519
rect 1452 3488 1501 3516
rect 1452 3476 1458 3488
rect 1489 3485 1501 3488
rect 1535 3485 1547 3519
rect 1489 3479 1547 3485
rect 2222 3476 2228 3528
rect 2280 3516 2286 3528
rect 2685 3519 2743 3525
rect 2685 3516 2697 3519
rect 2280 3488 2697 3516
rect 2280 3476 2286 3488
rect 2685 3485 2697 3488
rect 2731 3485 2743 3519
rect 2685 3479 2743 3485
rect 1949 3451 2007 3457
rect 1949 3417 1961 3451
rect 1995 3448 2007 3451
rect 1995 3420 2360 3448
rect 1995 3417 2007 3420
rect 1949 3411 2007 3417
rect 2130 3340 2136 3392
rect 2188 3389 2194 3392
rect 2188 3383 2207 3389
rect 2195 3349 2207 3383
rect 2332 3380 2360 3420
rect 2406 3408 2412 3460
rect 2464 3448 2470 3460
rect 2884 3448 2912 3547
rect 3142 3544 3148 3596
rect 3200 3544 3206 3596
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 4893 3587 4951 3593
rect 4893 3584 4905 3587
rect 3292 3556 4905 3584
rect 3292 3544 3298 3556
rect 4893 3553 4905 3556
rect 4939 3584 4951 3587
rect 7098 3584 7104 3596
rect 4939 3556 7104 3584
rect 4939 3553 4951 3556
rect 4893 3547 4951 3553
rect 7098 3544 7104 3556
rect 7156 3544 7162 3596
rect 7190 3544 7196 3596
rect 7248 3584 7254 3596
rect 7837 3587 7895 3593
rect 7837 3584 7849 3587
rect 7248 3556 7849 3584
rect 7248 3544 7254 3556
rect 7837 3553 7849 3556
rect 7883 3553 7895 3587
rect 7837 3547 7895 3553
rect 2961 3519 3019 3525
rect 2961 3485 2973 3519
rect 3007 3516 3019 3519
rect 3326 3516 3332 3528
rect 3007 3488 3332 3516
rect 3007 3485 3019 3488
rect 2961 3479 3019 3485
rect 3326 3476 3332 3488
rect 3384 3476 3390 3528
rect 3513 3519 3571 3525
rect 3513 3485 3525 3519
rect 3559 3516 3571 3519
rect 4617 3519 4675 3525
rect 4617 3516 4629 3519
rect 3559 3488 4629 3516
rect 3559 3485 3571 3488
rect 3513 3479 3571 3485
rect 4617 3485 4629 3488
rect 4663 3516 4675 3519
rect 4663 3488 4936 3516
rect 4663 3485 4675 3488
rect 4617 3479 4675 3485
rect 2464 3420 2912 3448
rect 2464 3408 2470 3420
rect 3050 3408 3056 3460
rect 3108 3448 3114 3460
rect 4065 3451 4123 3457
rect 4065 3448 4077 3451
rect 3108 3420 4077 3448
rect 3108 3408 3114 3420
rect 4065 3417 4077 3420
rect 4111 3448 4123 3451
rect 4798 3448 4804 3460
rect 4111 3420 4804 3448
rect 4111 3417 4123 3420
rect 4065 3411 4123 3417
rect 4798 3408 4804 3420
rect 4856 3408 4862 3460
rect 3694 3380 3700 3392
rect 2332 3352 3700 3380
rect 2188 3343 2207 3349
rect 2188 3340 2194 3343
rect 3694 3340 3700 3352
rect 3752 3340 3758 3392
rect 3786 3340 3792 3392
rect 3844 3380 3850 3392
rect 3973 3383 4031 3389
rect 3973 3380 3985 3383
rect 3844 3352 3985 3380
rect 3844 3340 3850 3352
rect 3973 3349 3985 3352
rect 4019 3349 4031 3383
rect 3973 3343 4031 3349
rect 4433 3383 4491 3389
rect 4433 3349 4445 3383
rect 4479 3380 4491 3383
rect 4706 3380 4712 3392
rect 4479 3352 4712 3380
rect 4479 3349 4491 3352
rect 4433 3343 4491 3349
rect 4706 3340 4712 3352
rect 4764 3340 4770 3392
rect 4908 3380 4936 3488
rect 7282 3476 7288 3528
rect 7340 3516 7346 3528
rect 7709 3519 7767 3525
rect 7709 3516 7721 3519
rect 7340 3488 7721 3516
rect 7340 3476 7346 3488
rect 7709 3485 7721 3488
rect 7755 3485 7767 3519
rect 7709 3479 7767 3485
rect 7926 3476 7932 3528
rect 7984 3476 7990 3528
rect 8110 3476 8116 3528
rect 8168 3476 8174 3528
rect 8404 3525 8432 3624
rect 10686 3612 10692 3664
rect 10744 3652 10750 3664
rect 11149 3655 11207 3661
rect 11149 3652 11161 3655
rect 10744 3624 11161 3652
rect 10744 3612 10750 3624
rect 11149 3621 11161 3624
rect 11195 3621 11207 3655
rect 15396 3652 15424 3683
rect 17034 3680 17040 3692
rect 17092 3680 17098 3732
rect 18506 3680 18512 3732
rect 18564 3720 18570 3732
rect 19797 3723 19855 3729
rect 19797 3720 19809 3723
rect 18564 3692 19809 3720
rect 18564 3680 18570 3692
rect 19797 3689 19809 3692
rect 19843 3689 19855 3723
rect 19797 3683 19855 3689
rect 19886 3680 19892 3732
rect 19944 3720 19950 3732
rect 20165 3723 20223 3729
rect 20165 3720 20177 3723
rect 19944 3692 20177 3720
rect 19944 3680 19950 3692
rect 20165 3689 20177 3692
rect 20211 3689 20223 3723
rect 20165 3683 20223 3689
rect 21358 3680 21364 3732
rect 21416 3720 21422 3732
rect 21910 3720 21916 3732
rect 21416 3692 21916 3720
rect 21416 3680 21422 3692
rect 21910 3680 21916 3692
rect 21968 3680 21974 3732
rect 22554 3680 22560 3732
rect 22612 3680 22618 3732
rect 23937 3723 23995 3729
rect 23937 3689 23949 3723
rect 23983 3720 23995 3723
rect 24026 3720 24032 3732
rect 23983 3692 24032 3720
rect 23983 3689 23995 3692
rect 23937 3683 23995 3689
rect 24026 3680 24032 3692
rect 24084 3680 24090 3732
rect 15396 3624 15470 3652
rect 11149 3615 11207 3621
rect 9309 3587 9367 3593
rect 9309 3553 9321 3587
rect 9355 3584 9367 3587
rect 9674 3584 9680 3596
rect 9355 3556 9680 3584
rect 9355 3553 9367 3556
rect 9309 3547 9367 3553
rect 9674 3544 9680 3556
rect 9732 3544 9738 3596
rect 11054 3544 11060 3596
rect 11112 3584 11118 3596
rect 11112 3556 11928 3584
rect 11112 3544 11118 3556
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3485 8447 3519
rect 8389 3479 8447 3485
rect 9033 3519 9091 3525
rect 9033 3485 9045 3519
rect 9079 3485 9091 3519
rect 9033 3479 9091 3485
rect 5166 3408 5172 3460
rect 5224 3408 5230 3460
rect 6178 3408 6184 3460
rect 6236 3408 6242 3460
rect 6730 3408 6736 3460
rect 6788 3448 6794 3460
rect 7009 3451 7067 3457
rect 7009 3448 7021 3451
rect 6788 3420 7021 3448
rect 6788 3408 6794 3420
rect 7009 3417 7021 3420
rect 7055 3448 7067 3451
rect 7055 3420 7328 3448
rect 7055 3417 7067 3420
rect 7009 3411 7067 3417
rect 5534 3380 5540 3392
rect 4908 3352 5540 3380
rect 5534 3340 5540 3352
rect 5592 3340 5598 3392
rect 5994 3340 6000 3392
rect 6052 3380 6058 3392
rect 6641 3383 6699 3389
rect 6641 3380 6653 3383
rect 6052 3352 6653 3380
rect 6052 3340 6058 3352
rect 6641 3349 6653 3352
rect 6687 3349 6699 3383
rect 6641 3343 6699 3349
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7209 3383 7267 3389
rect 7209 3380 7221 3383
rect 6972 3352 7221 3380
rect 6972 3340 6978 3352
rect 7209 3349 7221 3352
rect 7255 3349 7267 3383
rect 7300 3380 7328 3420
rect 7558 3408 7564 3460
rect 7616 3448 7622 3460
rect 7837 3451 7895 3457
rect 7837 3448 7849 3451
rect 7616 3420 7849 3448
rect 7616 3408 7622 3420
rect 7837 3417 7849 3420
rect 7883 3417 7895 3451
rect 9048 3448 9076 3479
rect 10870 3476 10876 3528
rect 10928 3516 10934 3528
rect 11793 3519 11851 3525
rect 11793 3516 11805 3519
rect 10928 3488 11805 3516
rect 10928 3476 10934 3488
rect 11793 3485 11805 3488
rect 11839 3485 11851 3519
rect 11900 3516 11928 3556
rect 13538 3544 13544 3596
rect 13596 3544 13602 3596
rect 13630 3544 13636 3596
rect 13688 3584 13694 3596
rect 13814 3584 13820 3596
rect 13688 3556 13820 3584
rect 13688 3544 13694 3556
rect 13814 3544 13820 3556
rect 13872 3544 13878 3596
rect 15442 3584 15470 3624
rect 15838 3612 15844 3664
rect 15896 3612 15902 3664
rect 19058 3612 19064 3664
rect 19116 3652 19122 3664
rect 19116 3624 20484 3652
rect 19116 3612 19122 3624
rect 14292 3556 15470 3584
rect 15856 3584 15884 3612
rect 18969 3587 19027 3593
rect 15856 3556 16160 3584
rect 14292 3528 14320 3556
rect 12069 3519 12127 3525
rect 12069 3516 12081 3519
rect 11900 3488 12081 3516
rect 11793 3479 11851 3485
rect 12069 3485 12081 3488
rect 12115 3485 12127 3519
rect 14090 3516 14096 3528
rect 12069 3479 12127 3485
rect 12820 3488 14096 3516
rect 9214 3448 9220 3460
rect 7837 3411 7895 3417
rect 7944 3420 8708 3448
rect 9048 3420 9220 3448
rect 7944 3380 7972 3420
rect 7300 3352 7972 3380
rect 7209 3343 7267 3349
rect 8018 3340 8024 3392
rect 8076 3380 8082 3392
rect 8573 3383 8631 3389
rect 8573 3380 8585 3383
rect 8076 3352 8585 3380
rect 8076 3340 8082 3352
rect 8573 3349 8585 3352
rect 8619 3349 8631 3383
rect 8680 3380 8708 3420
rect 9214 3408 9220 3420
rect 9272 3408 9278 3460
rect 10534 3420 11376 3448
rect 9398 3380 9404 3392
rect 8680 3352 9404 3380
rect 8573 3343 8631 3349
rect 9398 3340 9404 3352
rect 9456 3340 9462 3392
rect 11348 3380 11376 3420
rect 11422 3408 11428 3460
rect 11480 3408 11486 3460
rect 12820 3448 12848 3488
rect 14090 3476 14096 3488
rect 14148 3476 14154 3528
rect 14274 3476 14280 3528
rect 14332 3476 14338 3528
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3485 14611 3519
rect 14553 3479 14611 3485
rect 11992 3420 12848 3448
rect 11992 3380 12020 3420
rect 12894 3408 12900 3460
rect 12952 3448 12958 3460
rect 14568 3448 14596 3479
rect 14734 3476 14740 3528
rect 14792 3476 14798 3528
rect 15286 3476 15292 3528
rect 15344 3516 15350 3528
rect 15344 3488 15608 3516
rect 15344 3476 15350 3488
rect 15580 3457 15608 3488
rect 15746 3476 15752 3528
rect 15804 3516 15810 3528
rect 16132 3525 16160 3556
rect 18969 3553 18981 3587
rect 19015 3584 19027 3587
rect 19978 3584 19984 3596
rect 19015 3556 19984 3584
rect 19015 3553 19027 3556
rect 18969 3547 19027 3553
rect 19978 3544 19984 3556
rect 20036 3544 20042 3596
rect 15841 3519 15899 3525
rect 15841 3516 15853 3519
rect 15804 3488 15853 3516
rect 15804 3476 15810 3488
rect 15841 3485 15853 3488
rect 15887 3485 15899 3519
rect 15841 3479 15899 3485
rect 16117 3519 16175 3525
rect 16117 3485 16129 3519
rect 16163 3485 16175 3519
rect 16117 3479 16175 3485
rect 16209 3519 16267 3525
rect 16209 3485 16221 3519
rect 16255 3516 16267 3519
rect 16574 3516 16580 3528
rect 16255 3488 16580 3516
rect 16255 3485 16267 3488
rect 16209 3479 16267 3485
rect 16574 3476 16580 3488
rect 16632 3476 16638 3528
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3516 16727 3519
rect 16942 3516 16948 3528
rect 16715 3488 16948 3516
rect 16715 3485 16727 3488
rect 16669 3479 16727 3485
rect 16942 3476 16948 3488
rect 17000 3516 17006 3528
rect 17218 3516 17224 3528
rect 17000 3488 17224 3516
rect 17000 3476 17006 3488
rect 17218 3476 17224 3488
rect 17276 3476 17282 3528
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 19337 3519 19395 3525
rect 19337 3516 19349 3519
rect 19300 3488 19349 3516
rect 19300 3476 19306 3488
rect 19337 3485 19349 3488
rect 19383 3485 19395 3519
rect 19337 3479 19395 3485
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20070 3516 20076 3528
rect 19484 3488 20076 3516
rect 19484 3476 19490 3488
rect 20070 3476 20076 3488
rect 20128 3516 20134 3528
rect 20349 3519 20407 3525
rect 20349 3516 20361 3519
rect 20128 3488 20361 3516
rect 20128 3476 20134 3488
rect 20349 3485 20361 3488
rect 20395 3485 20407 3519
rect 20456 3516 20484 3624
rect 20714 3612 20720 3664
rect 20772 3652 20778 3664
rect 20772 3624 21404 3652
rect 20772 3612 20778 3624
rect 21376 3596 21404 3624
rect 21542 3612 21548 3664
rect 21600 3652 21606 3664
rect 23474 3652 23480 3664
rect 21600 3624 23480 3652
rect 21600 3612 21606 3624
rect 23474 3612 23480 3624
rect 23532 3612 23538 3664
rect 23753 3655 23811 3661
rect 23753 3621 23765 3655
rect 23799 3652 23811 3655
rect 24118 3652 24124 3664
rect 23799 3624 24124 3652
rect 23799 3621 23811 3624
rect 23753 3615 23811 3621
rect 24118 3612 24124 3624
rect 24176 3612 24182 3664
rect 21174 3544 21180 3596
rect 21232 3544 21238 3596
rect 21358 3544 21364 3596
rect 21416 3544 21422 3596
rect 21726 3544 21732 3596
rect 21784 3584 21790 3596
rect 23017 3587 23075 3593
rect 23017 3584 23029 3587
rect 21784 3556 23029 3584
rect 21784 3544 21790 3556
rect 23017 3553 23029 3556
rect 23063 3553 23075 3587
rect 23017 3547 23075 3553
rect 23106 3544 23112 3596
rect 23164 3544 23170 3596
rect 22094 3516 22100 3528
rect 20456 3488 22100 3516
rect 20349 3479 20407 3485
rect 22094 3476 22100 3488
rect 22152 3476 22158 3528
rect 22186 3476 22192 3528
rect 22244 3476 22250 3528
rect 22925 3519 22983 3525
rect 22925 3485 22937 3519
rect 22971 3516 22983 3519
rect 23290 3516 23296 3528
rect 22971 3488 23296 3516
rect 22971 3485 22983 3488
rect 22925 3479 22983 3485
rect 23290 3476 23296 3488
rect 23348 3476 23354 3528
rect 23566 3476 23572 3528
rect 23624 3516 23630 3528
rect 24578 3516 24584 3528
rect 23624 3488 24584 3516
rect 23624 3476 23630 3488
rect 24578 3476 24584 3488
rect 24636 3476 24642 3528
rect 15565 3451 15623 3457
rect 12952 3420 14596 3448
rect 15120 3420 15516 3448
rect 12952 3408 12958 3420
rect 11348 3352 12020 3380
rect 12066 3340 12072 3392
rect 12124 3380 12130 3392
rect 15120 3380 15148 3420
rect 12124 3352 15148 3380
rect 12124 3340 12130 3352
rect 15194 3340 15200 3392
rect 15252 3340 15258 3392
rect 15378 3389 15384 3392
rect 15365 3383 15384 3389
rect 15365 3349 15377 3383
rect 15365 3343 15384 3349
rect 15378 3340 15384 3343
rect 15436 3340 15442 3392
rect 15488 3380 15516 3420
rect 15565 3417 15577 3451
rect 15611 3417 15623 3451
rect 15565 3411 15623 3417
rect 16022 3408 16028 3460
rect 16080 3408 16086 3460
rect 16132 3420 17264 3448
rect 16132 3380 16160 3420
rect 15488 3352 16160 3380
rect 16850 3340 16856 3392
rect 16908 3340 16914 3392
rect 17236 3389 17264 3420
rect 18230 3408 18236 3460
rect 18288 3408 18294 3460
rect 18690 3408 18696 3460
rect 18748 3408 18754 3460
rect 18782 3408 18788 3460
rect 18840 3448 18846 3460
rect 18840 3420 21220 3448
rect 18840 3408 18846 3420
rect 17221 3383 17279 3389
rect 17221 3349 17233 3383
rect 17267 3380 17279 3383
rect 18598 3380 18604 3392
rect 17267 3352 18604 3380
rect 17267 3349 17279 3352
rect 17221 3343 17279 3349
rect 18598 3340 18604 3352
rect 18656 3340 18662 3392
rect 20622 3340 20628 3392
rect 20680 3340 20686 3392
rect 20990 3340 20996 3392
rect 21048 3340 21054 3392
rect 21082 3340 21088 3392
rect 21140 3340 21146 3392
rect 21192 3380 21220 3420
rect 21358 3408 21364 3460
rect 21416 3448 21422 3460
rect 21913 3451 21971 3457
rect 21913 3448 21925 3451
rect 21416 3420 21925 3448
rect 21416 3408 21422 3420
rect 21913 3417 21925 3420
rect 21959 3417 21971 3451
rect 21913 3411 21971 3417
rect 22370 3408 22376 3460
rect 22428 3448 22434 3460
rect 24121 3451 24179 3457
rect 24121 3448 24133 3451
rect 22428 3420 24133 3448
rect 22428 3408 22434 3420
rect 24121 3417 24133 3420
rect 24167 3448 24179 3451
rect 24670 3448 24676 3460
rect 24167 3420 24676 3448
rect 24167 3417 24179 3420
rect 24121 3411 24179 3417
rect 24670 3408 24676 3420
rect 24728 3408 24734 3460
rect 23566 3380 23572 3392
rect 21192 3352 23572 3380
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 23921 3383 23979 3389
rect 23921 3349 23933 3383
rect 23967 3380 23979 3383
rect 24762 3380 24768 3392
rect 23967 3352 24768 3380
rect 23967 3349 23979 3352
rect 23921 3343 23979 3349
rect 24762 3340 24768 3352
rect 24820 3340 24826 3392
rect 1104 3290 24840 3312
rect 1104 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 24214 3290
rect 24266 3238 24278 3290
rect 24330 3238 24342 3290
rect 24394 3238 24406 3290
rect 24458 3238 24470 3290
rect 24522 3238 24840 3290
rect 1104 3216 24840 3238
rect 2038 3136 2044 3188
rect 2096 3176 2102 3188
rect 2222 3176 2228 3188
rect 2096 3148 2228 3176
rect 2096 3136 2102 3148
rect 2222 3136 2228 3148
rect 2280 3136 2286 3188
rect 3697 3179 3755 3185
rect 3697 3145 3709 3179
rect 3743 3176 3755 3179
rect 5718 3176 5724 3188
rect 3743 3148 5724 3176
rect 3743 3145 3755 3148
rect 3697 3139 3755 3145
rect 5718 3136 5724 3148
rect 5776 3136 5782 3188
rect 5810 3136 5816 3188
rect 5868 3185 5874 3188
rect 5868 3179 5887 3185
rect 5875 3145 5887 3179
rect 5868 3139 5887 3145
rect 5997 3179 6055 3185
rect 5997 3145 6009 3179
rect 6043 3176 6055 3179
rect 6178 3176 6184 3188
rect 6043 3148 6184 3176
rect 6043 3145 6055 3148
rect 5997 3139 6055 3145
rect 5868 3136 5874 3139
rect 6178 3136 6184 3148
rect 6236 3136 6242 3188
rect 6546 3136 6552 3188
rect 6604 3176 6610 3188
rect 8297 3179 8355 3185
rect 6604 3148 8156 3176
rect 6604 3136 6610 3148
rect 2406 3108 2412 3120
rect 1780 3080 2412 3108
rect 1578 3000 1584 3052
rect 1636 3040 1642 3052
rect 1780 3049 1808 3080
rect 2406 3068 2412 3080
rect 2464 3068 2470 3120
rect 3050 3108 3056 3120
rect 2746 3080 3056 3108
rect 1765 3043 1823 3049
rect 1765 3040 1777 3043
rect 1636 3012 1777 3040
rect 1636 3000 1642 3012
rect 1765 3009 1777 3012
rect 1811 3009 1823 3043
rect 1765 3003 1823 3009
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2746 3040 2774 3080
rect 3050 3068 3056 3080
rect 3108 3068 3114 3120
rect 4157 3111 4215 3117
rect 4157 3077 4169 3111
rect 4203 3108 4215 3111
rect 4203 3080 4568 3108
rect 4203 3077 4215 3080
rect 4157 3071 4215 3077
rect 2271 3012 2774 3040
rect 2961 3043 3019 3049
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2961 3009 2973 3043
rect 3007 3040 3019 3043
rect 3142 3040 3148 3052
rect 3007 3012 3148 3040
rect 3007 3009 3019 3012
rect 2961 3003 3019 3009
rect 3142 3000 3148 3012
rect 3200 3000 3206 3052
rect 3510 3000 3516 3052
rect 3568 3040 3574 3052
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3568 3012 3617 3040
rect 3568 3000 3574 3012
rect 3605 3009 3617 3012
rect 3651 3009 3663 3043
rect 3605 3003 3663 3009
rect 3789 3043 3847 3049
rect 3789 3009 3801 3043
rect 3835 3040 3847 3043
rect 3970 3040 3976 3052
rect 3835 3012 3976 3040
rect 3835 3009 3847 3012
rect 3789 3003 3847 3009
rect 3970 3000 3976 3012
rect 4028 3000 4034 3052
rect 4540 3049 4568 3080
rect 4798 3068 4804 3120
rect 4856 3108 4862 3120
rect 4856 3080 5120 3108
rect 4856 3068 4862 3080
rect 4065 3043 4123 3049
rect 4065 3009 4077 3043
rect 4111 3009 4123 3043
rect 4065 3003 4123 3009
rect 4249 3043 4307 3049
rect 4249 3009 4261 3043
rect 4295 3009 4307 3043
rect 4249 3003 4307 3009
rect 4525 3043 4583 3049
rect 4525 3009 4537 3043
rect 4571 3009 4583 3043
rect 4525 3003 4583 3009
rect 4709 3043 4767 3049
rect 4709 3009 4721 3043
rect 4755 3009 4767 3043
rect 4709 3003 4767 3009
rect 2498 2932 2504 2984
rect 2556 2972 2562 2984
rect 2685 2975 2743 2981
rect 2685 2972 2697 2975
rect 2556 2944 2697 2972
rect 2556 2932 2562 2944
rect 2685 2941 2697 2944
rect 2731 2941 2743 2975
rect 2685 2935 2743 2941
rect 2869 2975 2927 2981
rect 2869 2941 2881 2975
rect 2915 2972 2927 2975
rect 3326 2972 3332 2984
rect 2915 2944 3332 2972
rect 2915 2941 2927 2944
rect 2869 2935 2927 2941
rect 3326 2932 3332 2944
rect 3384 2932 3390 2984
rect 4080 2972 4108 3003
rect 4264 2972 4292 3003
rect 4614 2972 4620 2984
rect 4080 2944 4200 2972
rect 4264 2944 4620 2972
rect 2409 2907 2467 2913
rect 2409 2873 2421 2907
rect 2455 2904 2467 2907
rect 4062 2904 4068 2916
rect 2455 2876 4068 2904
rect 2455 2873 2467 2876
rect 2409 2867 2467 2873
rect 4062 2864 4068 2876
rect 4120 2864 4126 2916
rect 4172 2904 4200 2944
rect 4614 2932 4620 2944
rect 4672 2932 4678 2984
rect 4724 2972 4752 3003
rect 4890 3000 4896 3052
rect 4948 3040 4954 3052
rect 5092 3049 5120 3080
rect 5442 3068 5448 3120
rect 5500 3108 5506 3120
rect 5629 3111 5687 3117
rect 5629 3108 5641 3111
rect 5500 3080 5641 3108
rect 5500 3068 5506 3080
rect 5629 3077 5641 3080
rect 5675 3108 5687 3111
rect 6270 3108 6276 3120
rect 5675 3080 6276 3108
rect 5675 3077 5687 3080
rect 5629 3071 5687 3077
rect 6270 3068 6276 3080
rect 6328 3068 6334 3120
rect 4985 3043 5043 3049
rect 4985 3040 4997 3043
rect 4948 3012 4997 3040
rect 4948 3000 4954 3012
rect 4985 3009 4997 3012
rect 5031 3009 5043 3043
rect 4985 3003 5043 3009
rect 5078 3043 5136 3049
rect 5078 3009 5090 3043
rect 5124 3009 5136 3043
rect 5078 3003 5136 3009
rect 5276 3012 6684 3040
rect 4798 2972 4804 2984
rect 4724 2944 4804 2972
rect 4798 2932 4804 2944
rect 4856 2932 4862 2984
rect 5276 2904 5304 3012
rect 6546 2932 6552 2984
rect 6604 2932 6610 2984
rect 6656 2972 6684 3012
rect 6730 3000 6736 3052
rect 6788 3000 6794 3052
rect 7282 3000 7288 3052
rect 7340 3000 7346 3052
rect 7837 3043 7895 3049
rect 7837 3009 7849 3043
rect 7883 3040 7895 3043
rect 8018 3040 8024 3052
rect 7883 3012 8024 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 8018 3000 8024 3012
rect 8076 3000 8082 3052
rect 8128 3049 8156 3148
rect 8297 3145 8309 3179
rect 8343 3145 8355 3179
rect 8297 3139 8355 3145
rect 8312 3108 8340 3139
rect 10594 3136 10600 3188
rect 10652 3176 10658 3188
rect 12805 3179 12863 3185
rect 10652 3148 12020 3176
rect 10652 3136 10658 3148
rect 11992 3117 12020 3148
rect 12805 3145 12817 3179
rect 12851 3176 12863 3179
rect 13354 3176 13360 3188
rect 12851 3148 13360 3176
rect 12851 3145 12863 3148
rect 12805 3139 12863 3145
rect 13354 3136 13360 3148
rect 13412 3136 13418 3188
rect 16022 3136 16028 3188
rect 16080 3136 16086 3188
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 17678 3176 17684 3188
rect 16908 3148 17684 3176
rect 16908 3136 16914 3148
rect 17678 3136 17684 3148
rect 17736 3176 17742 3188
rect 17789 3179 17847 3185
rect 17789 3176 17801 3179
rect 17736 3148 17801 3176
rect 17736 3136 17742 3148
rect 17789 3145 17801 3148
rect 17835 3145 17847 3179
rect 17789 3139 17847 3145
rect 17957 3179 18015 3185
rect 17957 3145 17969 3179
rect 18003 3176 18015 3179
rect 18233 3179 18291 3185
rect 18003 3148 18200 3176
rect 18003 3145 18015 3148
rect 17957 3139 18015 3145
rect 11977 3111 12035 3117
rect 8312 3080 11928 3108
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 9674 3040 9680 3052
rect 8159 3012 9680 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 9674 3000 9680 3012
rect 9732 3000 9738 3052
rect 9784 3049 9812 3080
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3009 9827 3043
rect 9769 3003 9827 3009
rect 10410 3000 10416 3052
rect 10468 3000 10474 3052
rect 10870 3000 10876 3052
rect 10928 3000 10934 3052
rect 11146 3000 11152 3052
rect 11204 3040 11210 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11204 3012 11621 3040
rect 11204 3000 11210 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11609 3003 11667 3009
rect 11793 3043 11851 3049
rect 11793 3009 11805 3043
rect 11839 3009 11851 3043
rect 11900 3040 11928 3080
rect 11977 3077 11989 3111
rect 12023 3077 12035 3111
rect 11977 3071 12035 3077
rect 12710 3068 12716 3120
rect 12768 3108 12774 3120
rect 13446 3108 13452 3120
rect 12768 3080 13452 3108
rect 12768 3068 12774 3080
rect 13446 3068 13452 3080
rect 13504 3068 13510 3120
rect 14737 3111 14795 3117
rect 14737 3108 14749 3111
rect 13556 3080 14749 3108
rect 11900 3012 12434 3040
rect 11793 3003 11851 3009
rect 8570 2972 8576 2984
rect 6656 2944 8576 2972
rect 8570 2932 8576 2944
rect 8628 2972 8634 2984
rect 9217 2975 9275 2981
rect 8628 2944 8800 2972
rect 8628 2932 8634 2944
rect 4172 2876 5304 2904
rect 5350 2864 5356 2916
rect 5408 2864 5414 2916
rect 5736 2876 6592 2904
rect 1857 2839 1915 2845
rect 1857 2805 1869 2839
rect 1903 2836 1915 2839
rect 2314 2836 2320 2848
rect 1903 2808 2320 2836
rect 1903 2805 1915 2808
rect 1857 2799 1915 2805
rect 2314 2796 2320 2808
rect 2372 2796 2378 2848
rect 2774 2796 2780 2848
rect 2832 2796 2838 2848
rect 4617 2839 4675 2845
rect 4617 2805 4629 2839
rect 4663 2836 4675 2839
rect 5736 2836 5764 2876
rect 4663 2808 5764 2836
rect 5813 2839 5871 2845
rect 4663 2805 4675 2808
rect 4617 2799 4675 2805
rect 5813 2805 5825 2839
rect 5859 2836 5871 2839
rect 6362 2836 6368 2848
rect 5859 2808 6368 2836
rect 5859 2805 5871 2808
rect 5813 2799 5871 2805
rect 6362 2796 6368 2808
rect 6420 2796 6426 2848
rect 6564 2836 6592 2876
rect 7466 2864 7472 2916
rect 7524 2864 7530 2916
rect 8772 2913 8800 2944
rect 9217 2941 9229 2975
rect 9263 2972 9275 2975
rect 9582 2972 9588 2984
rect 9263 2944 9588 2972
rect 9263 2941 9275 2944
rect 9217 2935 9275 2941
rect 9582 2932 9588 2944
rect 9640 2932 9646 2984
rect 10778 2932 10784 2984
rect 10836 2932 10842 2984
rect 11808 2972 11836 3003
rect 10980 2944 11836 2972
rect 10980 2916 11008 2944
rect 11882 2932 11888 2984
rect 11940 2972 11946 2984
rect 12253 2975 12311 2981
rect 12253 2972 12265 2975
rect 11940 2944 12265 2972
rect 11940 2932 11946 2944
rect 12253 2941 12265 2944
rect 12299 2941 12311 2975
rect 12406 2972 12434 3012
rect 12802 3000 12808 3052
rect 12860 3000 12866 3052
rect 13556 3049 13584 3080
rect 14737 3077 14749 3080
rect 14783 3077 14795 3111
rect 14737 3071 14795 3077
rect 17586 3068 17592 3120
rect 17644 3068 17650 3120
rect 18172 3108 18200 3148
rect 18233 3145 18245 3179
rect 18279 3176 18291 3179
rect 18690 3176 18696 3188
rect 18279 3148 18696 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18690 3136 18696 3148
rect 18748 3136 18754 3188
rect 18966 3136 18972 3188
rect 19024 3176 19030 3188
rect 19429 3179 19487 3185
rect 19429 3176 19441 3179
rect 19024 3148 19441 3176
rect 19024 3136 19030 3148
rect 19429 3145 19441 3148
rect 19475 3145 19487 3179
rect 20990 3176 20996 3188
rect 19429 3139 19487 3145
rect 19720 3148 20996 3176
rect 18506 3108 18512 3120
rect 18172 3080 18512 3108
rect 18506 3068 18512 3080
rect 18564 3068 18570 3120
rect 18598 3068 18604 3120
rect 18656 3068 18662 3120
rect 19720 3108 19748 3148
rect 20990 3136 20996 3148
rect 21048 3176 21054 3188
rect 21545 3179 21603 3185
rect 21545 3176 21557 3179
rect 21048 3148 21557 3176
rect 21048 3136 21054 3148
rect 21545 3145 21557 3148
rect 21591 3145 21603 3179
rect 21545 3139 21603 3145
rect 21913 3179 21971 3185
rect 21913 3145 21925 3179
rect 21959 3145 21971 3179
rect 21913 3139 21971 3145
rect 19978 3108 19984 3120
rect 18708 3080 19748 3108
rect 19812 3080 19984 3108
rect 13541 3043 13599 3049
rect 13541 3009 13553 3043
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 13998 3000 14004 3052
rect 14056 3000 14062 3052
rect 14182 3000 14188 3052
rect 14240 3000 14246 3052
rect 14645 3043 14703 3049
rect 14645 3009 14657 3043
rect 14691 3009 14703 3043
rect 14645 3003 14703 3009
rect 15013 3043 15071 3049
rect 15013 3009 15025 3043
rect 15059 3040 15071 3043
rect 15102 3040 15108 3052
rect 15059 3012 15108 3040
rect 15059 3009 15071 3012
rect 15013 3003 15071 3009
rect 12710 2972 12716 2984
rect 12406 2944 12716 2972
rect 12253 2935 12311 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 12894 2932 12900 2984
rect 12952 2932 12958 2984
rect 13262 2932 13268 2984
rect 13320 2932 13326 2984
rect 14660 2972 14688 3003
rect 15102 3000 15108 3012
rect 15160 3000 15166 3052
rect 15194 3000 15200 3052
rect 15252 3000 15258 3052
rect 15470 3000 15476 3052
rect 15528 3040 15534 3052
rect 15565 3043 15623 3049
rect 15565 3040 15577 3043
rect 15528 3012 15577 3040
rect 15528 3000 15534 3012
rect 15565 3009 15577 3012
rect 15611 3009 15623 3043
rect 15565 3003 15623 3009
rect 15841 3043 15899 3049
rect 15841 3009 15853 3043
rect 15887 3040 15899 3043
rect 16850 3040 16856 3052
rect 15887 3012 16856 3040
rect 15887 3009 15899 3012
rect 15841 3003 15899 3009
rect 16850 3000 16856 3012
rect 16908 3040 16914 3052
rect 17310 3040 17316 3052
rect 16908 3012 17316 3040
rect 16908 3000 16914 3012
rect 17310 3000 17316 3012
rect 17368 3040 17374 3052
rect 17494 3040 17500 3052
rect 17368 3012 17500 3040
rect 17368 3000 17374 3012
rect 17494 3000 17500 3012
rect 17552 3000 17558 3052
rect 18708 3049 18736 3080
rect 19812 3052 19840 3080
rect 19978 3068 19984 3080
rect 20036 3068 20042 3120
rect 21928 3108 21956 3139
rect 22554 3136 22560 3188
rect 22612 3176 22618 3188
rect 23382 3176 23388 3188
rect 22612 3148 23388 3176
rect 22612 3136 22618 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 22094 3117 22100 3120
rect 21298 3080 21956 3108
rect 22081 3111 22100 3117
rect 22081 3077 22093 3111
rect 22081 3071 22100 3077
rect 22094 3068 22100 3071
rect 22152 3068 22158 3120
rect 22281 3111 22339 3117
rect 22281 3077 22293 3111
rect 22327 3108 22339 3111
rect 22370 3108 22376 3120
rect 22327 3080 22376 3108
rect 22327 3077 22339 3080
rect 22281 3071 22339 3077
rect 22370 3068 22376 3080
rect 22428 3068 22434 3120
rect 23750 3068 23756 3120
rect 23808 3108 23814 3120
rect 23808 3080 24348 3108
rect 23808 3068 23814 3080
rect 18693 3043 18751 3049
rect 18693 3009 18705 3043
rect 18739 3009 18751 3043
rect 18693 3003 18751 3009
rect 19245 3043 19303 3049
rect 19245 3009 19257 3043
rect 19291 3040 19303 3043
rect 19334 3040 19340 3052
rect 19291 3012 19340 3040
rect 19291 3009 19303 3012
rect 19245 3003 19303 3009
rect 19334 3000 19340 3012
rect 19392 3000 19398 3052
rect 19794 3000 19800 3052
rect 19852 3000 19858 3052
rect 21634 3000 21640 3052
rect 21692 3040 21698 3052
rect 24320 3049 24348 3080
rect 24305 3043 24363 3049
rect 21692 3012 22954 3040
rect 21692 3000 21698 3012
rect 24305 3009 24317 3043
rect 24351 3009 24363 3043
rect 24305 3003 24363 3009
rect 14918 2972 14924 2984
rect 14660 2944 14924 2972
rect 14918 2932 14924 2944
rect 14976 2932 14982 2984
rect 15746 2932 15752 2984
rect 15804 2972 15810 2984
rect 16114 2972 16120 2984
rect 15804 2944 16120 2972
rect 15804 2932 15810 2944
rect 16114 2932 16120 2944
rect 16172 2972 16178 2984
rect 16761 2975 16819 2981
rect 16761 2972 16773 2975
rect 16172 2944 16773 2972
rect 16172 2932 16178 2944
rect 16761 2941 16773 2944
rect 16807 2972 16819 2975
rect 17218 2972 17224 2984
rect 16807 2944 17224 2972
rect 16807 2941 16819 2944
rect 16761 2935 16819 2941
rect 17218 2932 17224 2944
rect 17276 2932 17282 2984
rect 18877 2975 18935 2981
rect 18877 2941 18889 2975
rect 18923 2972 18935 2975
rect 20073 2975 20131 2981
rect 18923 2944 19748 2972
rect 18923 2941 18935 2944
rect 18877 2935 18935 2941
rect 8757 2907 8815 2913
rect 8757 2873 8769 2907
rect 8803 2873 8815 2907
rect 8757 2867 8815 2873
rect 9306 2864 9312 2916
rect 9364 2904 9370 2916
rect 9364 2876 10088 2904
rect 9364 2864 9370 2876
rect 7558 2836 7564 2848
rect 6564 2808 7564 2836
rect 7558 2796 7564 2808
rect 7616 2796 7622 2848
rect 7742 2796 7748 2848
rect 7800 2836 7806 2848
rect 9030 2836 9036 2848
rect 7800 2808 9036 2836
rect 7800 2796 7806 2808
rect 9030 2796 9036 2808
rect 9088 2796 9094 2848
rect 9950 2796 9956 2848
rect 10008 2796 10014 2848
rect 10060 2836 10088 2876
rect 10962 2864 10968 2916
rect 11020 2864 11026 2916
rect 11241 2907 11299 2913
rect 11241 2873 11253 2907
rect 11287 2904 11299 2907
rect 11330 2904 11336 2916
rect 11287 2876 11336 2904
rect 11287 2873 11299 2876
rect 11241 2867 11299 2873
rect 11330 2864 11336 2876
rect 11388 2864 11394 2916
rect 11624 2876 12434 2904
rect 11624 2836 11652 2876
rect 10060 2808 11652 2836
rect 12406 2836 12434 2876
rect 14826 2864 14832 2916
rect 14884 2904 14890 2916
rect 15657 2907 15715 2913
rect 15657 2904 15669 2907
rect 14884 2876 15669 2904
rect 14884 2864 14890 2876
rect 15657 2873 15669 2876
rect 15703 2873 15715 2907
rect 15657 2867 15715 2873
rect 16393 2907 16451 2913
rect 16393 2873 16405 2907
rect 16439 2904 16451 2907
rect 19610 2904 19616 2916
rect 16439 2876 19616 2904
rect 16439 2873 16451 2876
rect 16393 2867 16451 2873
rect 19610 2864 19616 2876
rect 19668 2864 19674 2916
rect 13538 2836 13544 2848
rect 12406 2808 13544 2836
rect 13538 2796 13544 2808
rect 13596 2796 13602 2848
rect 15010 2796 15016 2848
rect 15068 2836 15074 2848
rect 15470 2836 15476 2848
rect 15068 2808 15476 2836
rect 15068 2796 15074 2808
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 17221 2839 17279 2845
rect 17221 2805 17233 2839
rect 17267 2836 17279 2839
rect 17678 2836 17684 2848
rect 17267 2808 17684 2836
rect 17267 2805 17279 2808
rect 17221 2799 17279 2805
rect 17678 2796 17684 2808
rect 17736 2796 17742 2848
rect 17773 2839 17831 2845
rect 17773 2805 17785 2839
rect 17819 2836 17831 2839
rect 18230 2836 18236 2848
rect 17819 2808 18236 2836
rect 17819 2805 17831 2808
rect 17773 2799 17831 2805
rect 18230 2796 18236 2808
rect 18288 2836 18294 2848
rect 18966 2836 18972 2848
rect 18288 2808 18972 2836
rect 18288 2796 18294 2808
rect 18966 2796 18972 2808
rect 19024 2796 19030 2848
rect 19518 2796 19524 2848
rect 19576 2836 19582 2848
rect 19720 2836 19748 2944
rect 20073 2941 20085 2975
rect 20119 2972 20131 2975
rect 20622 2972 20628 2984
rect 20119 2944 20628 2972
rect 20119 2941 20131 2944
rect 20073 2935 20131 2941
rect 20622 2932 20628 2944
rect 20680 2932 20686 2984
rect 20806 2932 20812 2984
rect 20864 2972 20870 2984
rect 21266 2972 21272 2984
rect 20864 2944 21272 2972
rect 20864 2932 20870 2944
rect 21266 2932 21272 2944
rect 21324 2972 21330 2984
rect 21324 2944 22140 2972
rect 21324 2932 21330 2944
rect 21174 2836 21180 2848
rect 19576 2808 21180 2836
rect 19576 2796 19582 2808
rect 21174 2796 21180 2808
rect 21232 2796 21238 2848
rect 22112 2845 22140 2944
rect 23934 2932 23940 2984
rect 23992 2972 23998 2984
rect 24029 2975 24087 2981
rect 24029 2972 24041 2975
rect 23992 2944 24041 2972
rect 23992 2932 23998 2944
rect 24029 2941 24041 2944
rect 24075 2941 24087 2975
rect 24029 2935 24087 2941
rect 22112 2839 22195 2845
rect 22112 2808 22149 2839
rect 22137 2805 22149 2808
rect 22183 2836 22195 2839
rect 24026 2836 24032 2848
rect 22183 2808 24032 2836
rect 22183 2805 22195 2808
rect 22137 2799 22195 2805
rect 24026 2796 24032 2808
rect 24084 2796 24090 2848
rect 1104 2746 24840 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 20214 2746
rect 20266 2694 20278 2746
rect 20330 2694 20342 2746
rect 20394 2694 20406 2746
rect 20458 2694 20470 2746
rect 20522 2694 24840 2746
rect 1104 2672 24840 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 3142 2632 3148 2644
rect 1903 2604 3148 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 3142 2592 3148 2604
rect 3200 2592 3206 2644
rect 6546 2632 6552 2644
rect 3436 2604 6552 2632
rect 2774 2564 2780 2576
rect 2424 2536 2780 2564
rect 2424 2505 2452 2536
rect 2774 2524 2780 2536
rect 2832 2524 2838 2576
rect 3436 2573 3464 2604
rect 6546 2592 6552 2604
rect 6604 2592 6610 2644
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 10686 2632 10692 2644
rect 7248 2604 8156 2632
rect 7248 2592 7254 2604
rect 3421 2567 3479 2573
rect 3421 2533 3433 2567
rect 3467 2533 3479 2567
rect 7742 2564 7748 2576
rect 3421 2527 3479 2533
rect 4540 2536 7748 2564
rect 2409 2499 2467 2505
rect 2409 2465 2421 2499
rect 2455 2465 2467 2499
rect 2409 2459 2467 2465
rect 2682 2456 2688 2508
rect 2740 2456 2746 2508
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2397 1731 2431
rect 1673 2391 1731 2397
rect 1302 2320 1308 2372
rect 1360 2360 1366 2372
rect 1688 2360 1716 2391
rect 2314 2388 2320 2440
rect 2372 2388 2378 2440
rect 2961 2431 3019 2437
rect 2961 2397 2973 2431
rect 3007 2428 3019 2431
rect 3050 2428 3056 2440
rect 3007 2400 3056 2428
rect 3007 2397 3019 2400
rect 2961 2391 3019 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 3145 2431 3203 2437
rect 3145 2397 3157 2431
rect 3191 2428 3203 2431
rect 3326 2428 3332 2440
rect 3191 2400 3332 2428
rect 3191 2397 3203 2400
rect 3145 2391 3203 2397
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 3513 2431 3571 2437
rect 3513 2397 3525 2431
rect 3559 2397 3571 2431
rect 3513 2391 3571 2397
rect 2866 2360 2872 2372
rect 1360 2332 2872 2360
rect 1360 2320 1366 2332
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 3528 2360 3556 2391
rect 3970 2388 3976 2440
rect 4028 2388 4034 2440
rect 4540 2437 4568 2536
rect 7742 2524 7748 2536
rect 7800 2524 7806 2576
rect 8128 2564 8156 2604
rect 8496 2604 10692 2632
rect 8496 2564 8524 2604
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 11425 2635 11483 2641
rect 11425 2601 11437 2635
rect 11471 2632 11483 2635
rect 11514 2632 11520 2644
rect 11471 2604 11520 2632
rect 11471 2601 11483 2604
rect 11425 2595 11483 2601
rect 11514 2592 11520 2604
rect 11572 2592 11578 2644
rect 17681 2635 17739 2641
rect 17681 2601 17693 2635
rect 17727 2632 17739 2635
rect 17770 2632 17776 2644
rect 17727 2604 17776 2632
rect 17727 2601 17739 2604
rect 17681 2595 17739 2601
rect 17770 2592 17776 2604
rect 17828 2592 17834 2644
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18141 2635 18199 2641
rect 18141 2632 18153 2635
rect 18012 2604 18153 2632
rect 18012 2592 18018 2604
rect 18141 2601 18153 2604
rect 18187 2601 18199 2635
rect 18141 2595 18199 2601
rect 18509 2635 18567 2641
rect 18509 2601 18521 2635
rect 18555 2632 18567 2635
rect 18782 2632 18788 2644
rect 18555 2604 18788 2632
rect 18555 2601 18567 2604
rect 18509 2595 18567 2601
rect 18782 2592 18788 2604
rect 18840 2592 18846 2644
rect 20070 2592 20076 2644
rect 20128 2632 20134 2644
rect 22462 2632 22468 2644
rect 20128 2604 22468 2632
rect 20128 2592 20134 2604
rect 22462 2592 22468 2604
rect 22520 2592 22526 2644
rect 8128 2536 8524 2564
rect 4632 2468 4844 2496
rect 4525 2431 4583 2437
rect 4525 2397 4537 2431
rect 4571 2397 4583 2431
rect 4525 2391 4583 2397
rect 4632 2360 4660 2468
rect 4816 2440 4844 2468
rect 5350 2456 5356 2508
rect 5408 2496 5414 2508
rect 5408 2468 6316 2496
rect 5408 2456 5414 2468
rect 4709 2431 4767 2437
rect 4709 2397 4721 2431
rect 4755 2397 4767 2431
rect 4709 2391 4767 2397
rect 3528 2332 4660 2360
rect 4724 2292 4752 2391
rect 4798 2388 4804 2440
rect 4856 2428 4862 2440
rect 5537 2431 5595 2437
rect 5537 2428 5549 2431
rect 4856 2400 5549 2428
rect 4856 2388 4862 2400
rect 5537 2397 5549 2400
rect 5583 2397 5595 2431
rect 5537 2391 5595 2397
rect 5718 2388 5724 2440
rect 5776 2428 5782 2440
rect 6288 2437 6316 2468
rect 6730 2456 6736 2508
rect 6788 2456 6794 2508
rect 7834 2456 7840 2508
rect 7892 2456 7898 2508
rect 8110 2456 8116 2508
rect 8168 2496 8174 2508
rect 8205 2499 8263 2505
rect 8205 2496 8217 2499
rect 8168 2468 8217 2496
rect 8168 2456 8174 2468
rect 8205 2465 8217 2468
rect 8251 2465 8263 2499
rect 8205 2459 8263 2465
rect 8496 2447 8524 2536
rect 9030 2524 9036 2576
rect 9088 2564 9094 2576
rect 9585 2567 9643 2573
rect 9585 2564 9597 2567
rect 9088 2536 9597 2564
rect 9088 2524 9094 2536
rect 9585 2533 9597 2536
rect 9631 2533 9643 2567
rect 12618 2564 12624 2576
rect 9585 2527 9643 2533
rect 11532 2536 12624 2564
rect 8846 2456 8852 2508
rect 8904 2496 8910 2508
rect 9858 2496 9864 2508
rect 8904 2468 9864 2496
rect 8904 2456 8910 2468
rect 9858 2456 9864 2468
rect 9916 2456 9922 2508
rect 11241 2499 11299 2505
rect 11241 2465 11253 2499
rect 11287 2496 11299 2499
rect 11532 2496 11560 2536
rect 12618 2524 12624 2536
rect 12676 2524 12682 2576
rect 13170 2524 13176 2576
rect 13228 2564 13234 2576
rect 13541 2567 13599 2573
rect 13541 2564 13553 2567
rect 13228 2536 13553 2564
rect 13228 2524 13234 2536
rect 13541 2533 13553 2536
rect 13587 2533 13599 2567
rect 13541 2527 13599 2533
rect 13998 2524 14004 2576
rect 14056 2564 14062 2576
rect 14056 2536 15884 2564
rect 14056 2524 14062 2536
rect 14185 2499 14243 2505
rect 14185 2496 14197 2499
rect 11287 2468 11560 2496
rect 11623 2468 12480 2496
rect 11287 2465 11299 2468
rect 11241 2459 11299 2465
rect 8481 2441 8539 2447
rect 5813 2431 5871 2437
rect 5813 2428 5825 2431
rect 5776 2400 5825 2428
rect 5776 2388 5782 2400
rect 5813 2397 5825 2400
rect 5859 2397 5871 2431
rect 5813 2391 5871 2397
rect 6273 2431 6331 2437
rect 6273 2397 6285 2431
rect 6319 2397 6331 2431
rect 6273 2391 6331 2397
rect 6822 2388 6828 2440
rect 6880 2388 6886 2440
rect 7006 2388 7012 2440
rect 7064 2428 7070 2440
rect 7469 2431 7527 2437
rect 7469 2428 7481 2431
rect 7064 2400 7481 2428
rect 7064 2388 7070 2400
rect 7469 2397 7481 2400
rect 7515 2428 7527 2431
rect 7650 2428 7656 2440
rect 7515 2400 7656 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 7745 2431 7803 2437
rect 7745 2397 7757 2431
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 5077 2363 5135 2369
rect 5077 2329 5089 2363
rect 5123 2360 5135 2363
rect 7760 2360 7788 2391
rect 7926 2388 7932 2440
rect 7984 2388 7990 2440
rect 8018 2388 8024 2440
rect 8076 2428 8082 2440
rect 8076 2422 8340 2428
rect 8377 2425 8435 2431
rect 8377 2422 8389 2425
rect 8076 2400 8389 2422
rect 8076 2388 8082 2400
rect 8312 2394 8389 2400
rect 8377 2391 8389 2394
rect 8423 2391 8435 2425
rect 8481 2407 8493 2441
rect 8527 2407 8539 2441
rect 8481 2401 8539 2407
rect 8377 2385 8435 2391
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 9033 2431 9091 2437
rect 9033 2397 9045 2431
rect 9079 2430 9091 2431
rect 10045 2431 10103 2437
rect 9079 2402 9168 2430
rect 9079 2397 9091 2402
rect 9033 2391 9091 2397
rect 8110 2360 8116 2372
rect 5123 2332 7696 2360
rect 7760 2332 8116 2360
rect 5123 2329 5135 2332
rect 5077 2323 5135 2329
rect 6638 2292 6644 2304
rect 4724 2264 6644 2292
rect 6638 2252 6644 2264
rect 6696 2252 6702 2304
rect 7668 2292 7696 2332
rect 8110 2320 8116 2332
rect 8168 2320 8174 2372
rect 9140 2360 9168 2402
rect 10045 2397 10057 2431
rect 10091 2428 10103 2431
rect 10597 2431 10655 2437
rect 10091 2400 10548 2428
rect 10091 2397 10103 2400
rect 10045 2391 10103 2397
rect 9140 2332 9904 2360
rect 9030 2292 9036 2304
rect 7668 2264 9036 2292
rect 9030 2252 9036 2264
rect 9088 2252 9094 2304
rect 9217 2295 9275 2301
rect 9217 2261 9229 2295
rect 9263 2292 9275 2295
rect 9674 2292 9680 2304
rect 9263 2264 9680 2292
rect 9263 2261 9275 2264
rect 9217 2255 9275 2261
rect 9674 2252 9680 2264
rect 9732 2252 9738 2304
rect 9876 2292 9904 2332
rect 10410 2292 10416 2304
rect 9876 2264 10416 2292
rect 10410 2252 10416 2264
rect 10468 2252 10474 2304
rect 10520 2292 10548 2400
rect 10597 2397 10609 2431
rect 10643 2428 10655 2431
rect 10686 2428 10692 2440
rect 10643 2400 10692 2428
rect 10643 2397 10655 2400
rect 10597 2391 10655 2397
rect 10686 2388 10692 2400
rect 10744 2388 10750 2440
rect 11146 2388 11152 2440
rect 11204 2388 11210 2440
rect 11330 2320 11336 2372
rect 11388 2360 11394 2372
rect 11623 2360 11651 2468
rect 12452 2437 12480 2468
rect 13188 2468 14197 2496
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12345 2431 12403 2437
rect 12345 2397 12357 2431
rect 12391 2397 12403 2431
rect 12345 2391 12403 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2397 12495 2431
rect 12437 2391 12495 2397
rect 11388 2332 11651 2360
rect 11388 2320 11394 2332
rect 11992 2304 12020 2391
rect 12360 2360 12388 2391
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 12986 2428 12992 2440
rect 12676 2400 12992 2428
rect 12676 2388 12682 2400
rect 12986 2388 12992 2400
rect 13044 2388 13050 2440
rect 13188 2437 13216 2468
rect 14185 2465 14197 2468
rect 14231 2465 14243 2499
rect 14185 2459 14243 2465
rect 14734 2456 14740 2508
rect 14792 2456 14798 2508
rect 15378 2456 15384 2508
rect 15436 2496 15442 2508
rect 15856 2505 15884 2536
rect 18690 2524 18696 2576
rect 18748 2524 18754 2576
rect 20898 2564 20904 2576
rect 19444 2536 20904 2564
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 15436 2468 15577 2496
rect 15436 2456 15442 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 15841 2499 15899 2505
rect 15841 2465 15853 2499
rect 15887 2496 15899 2499
rect 15930 2496 15936 2508
rect 15887 2468 15936 2496
rect 15887 2465 15899 2468
rect 15841 2459 15899 2465
rect 15930 2456 15936 2468
rect 15988 2456 15994 2508
rect 16117 2499 16175 2505
rect 16117 2465 16129 2499
rect 16163 2496 16175 2499
rect 16577 2499 16635 2505
rect 16577 2496 16589 2499
rect 16163 2468 16589 2496
rect 16163 2465 16175 2468
rect 16117 2459 16175 2465
rect 16577 2465 16589 2468
rect 16623 2465 16635 2499
rect 16577 2459 16635 2465
rect 16666 2456 16672 2508
rect 16724 2456 16730 2508
rect 16761 2499 16819 2505
rect 16761 2465 16773 2499
rect 16807 2496 16819 2499
rect 16850 2496 16856 2508
rect 16807 2468 16856 2496
rect 16807 2465 16819 2468
rect 16761 2459 16819 2465
rect 16850 2456 16856 2468
rect 16908 2456 16914 2508
rect 16945 2499 17003 2505
rect 16945 2465 16957 2499
rect 16991 2496 17003 2499
rect 17034 2496 17040 2508
rect 16991 2468 17040 2496
rect 16991 2465 17003 2468
rect 16945 2459 17003 2465
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 17218 2456 17224 2508
rect 17276 2456 17282 2508
rect 17586 2456 17592 2508
rect 17644 2496 17650 2508
rect 17770 2496 17776 2508
rect 17644 2468 17776 2496
rect 17644 2456 17650 2468
rect 17770 2456 17776 2468
rect 17828 2456 17834 2508
rect 13173 2431 13231 2437
rect 13173 2397 13185 2431
rect 13219 2397 13231 2431
rect 13173 2391 13231 2397
rect 13354 2388 13360 2440
rect 13412 2388 13418 2440
rect 15013 2431 15071 2437
rect 15013 2397 15025 2431
rect 15059 2428 15071 2431
rect 15746 2428 15752 2440
rect 15059 2400 15752 2428
rect 15059 2397 15071 2400
rect 15013 2391 15071 2397
rect 15746 2388 15752 2400
rect 15804 2388 15810 2440
rect 16022 2388 16028 2440
rect 16080 2388 16086 2440
rect 16485 2431 16543 2437
rect 16485 2397 16497 2431
rect 16531 2397 16543 2431
rect 16485 2391 16543 2397
rect 12802 2360 12808 2372
rect 12360 2332 12808 2360
rect 12802 2320 12808 2332
rect 12860 2320 12866 2372
rect 15930 2320 15936 2372
rect 15988 2320 15994 2372
rect 16500 2360 16528 2391
rect 17678 2388 17684 2440
rect 17736 2428 17742 2440
rect 18049 2431 18107 2437
rect 18049 2428 18061 2431
rect 17736 2400 18061 2428
rect 17736 2388 17742 2400
rect 18049 2397 18061 2400
rect 18095 2397 18107 2431
rect 18049 2391 18107 2397
rect 18138 2388 18144 2440
rect 18196 2428 18202 2440
rect 18233 2431 18291 2437
rect 18233 2428 18245 2431
rect 18196 2400 18245 2428
rect 18196 2388 18202 2400
rect 18233 2397 18245 2400
rect 18279 2428 18291 2431
rect 19242 2428 19248 2440
rect 18279 2400 19248 2428
rect 18279 2397 18291 2400
rect 18233 2391 18291 2397
rect 19242 2388 19248 2400
rect 19300 2388 19306 2440
rect 17586 2360 17592 2372
rect 16500 2332 17592 2360
rect 17586 2320 17592 2332
rect 17644 2320 17650 2372
rect 18966 2320 18972 2372
rect 19024 2320 19030 2372
rect 11422 2292 11428 2304
rect 10520 2264 11428 2292
rect 11422 2252 11428 2264
rect 11480 2252 11486 2304
rect 11974 2252 11980 2304
rect 12032 2252 12038 2304
rect 15470 2252 15476 2304
rect 15528 2292 15534 2304
rect 19444 2292 19472 2536
rect 20898 2524 20904 2536
rect 20956 2564 20962 2576
rect 22373 2567 22431 2573
rect 22373 2564 22385 2567
rect 20956 2536 22385 2564
rect 20956 2524 20962 2536
rect 22373 2533 22385 2536
rect 22419 2533 22431 2567
rect 22373 2527 22431 2533
rect 19518 2456 19524 2508
rect 19576 2456 19582 2508
rect 19705 2499 19763 2505
rect 19705 2465 19717 2499
rect 19751 2496 19763 2499
rect 22554 2496 22560 2508
rect 19751 2468 22560 2496
rect 19751 2465 19763 2468
rect 19705 2459 19763 2465
rect 22554 2456 22560 2468
rect 22612 2456 22618 2508
rect 23106 2456 23112 2508
rect 23164 2496 23170 2508
rect 23661 2499 23719 2505
rect 23661 2496 23673 2499
rect 23164 2468 23673 2496
rect 23164 2456 23170 2468
rect 23661 2465 23673 2468
rect 23707 2465 23719 2499
rect 23661 2459 23719 2465
rect 19610 2388 19616 2440
rect 19668 2428 19674 2440
rect 20622 2428 20628 2440
rect 19668 2400 20628 2428
rect 19668 2388 19674 2400
rect 20622 2388 20628 2400
rect 20680 2388 20686 2440
rect 21637 2431 21695 2437
rect 21637 2397 21649 2431
rect 21683 2428 21695 2431
rect 22186 2428 22192 2440
rect 21683 2400 22192 2428
rect 21683 2397 21695 2400
rect 21637 2391 21695 2397
rect 22186 2388 22192 2400
rect 22244 2428 22250 2440
rect 22281 2431 22339 2437
rect 22281 2428 22293 2431
rect 22244 2400 22293 2428
rect 22244 2388 22250 2400
rect 22281 2397 22293 2400
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 23014 2388 23020 2440
rect 23072 2428 23078 2440
rect 23477 2431 23535 2437
rect 23477 2428 23489 2431
rect 23072 2400 23489 2428
rect 23072 2388 23078 2400
rect 23477 2397 23489 2400
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 19797 2363 19855 2369
rect 19797 2329 19809 2363
rect 19843 2360 19855 2363
rect 21082 2360 21088 2372
rect 19843 2332 21088 2360
rect 19843 2329 19855 2332
rect 19797 2323 19855 2329
rect 21082 2320 21088 2332
rect 21140 2320 21146 2372
rect 15528 2264 19472 2292
rect 15528 2252 15534 2264
rect 20070 2252 20076 2304
rect 20128 2292 20134 2304
rect 20165 2295 20223 2301
rect 20165 2292 20177 2295
rect 20128 2264 20177 2292
rect 20128 2252 20134 2264
rect 20165 2261 20177 2264
rect 20211 2261 20223 2295
rect 20165 2255 20223 2261
rect 1104 2202 24840 2224
rect 1104 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 24214 2202
rect 24266 2150 24278 2202
rect 24330 2150 24342 2202
rect 24394 2150 24406 2202
rect 24458 2150 24470 2202
rect 24522 2150 24840 2202
rect 1104 2128 24840 2150
rect 1489 2091 1547 2097
rect 1489 2057 1501 2091
rect 1535 2088 1547 2091
rect 1578 2088 1584 2100
rect 1535 2060 1584 2088
rect 1535 2057 1547 2060
rect 1489 2051 1547 2057
rect 1578 2048 1584 2060
rect 1636 2048 1642 2100
rect 3970 2048 3976 2100
rect 4028 2048 4034 2100
rect 4249 2091 4307 2097
rect 4249 2057 4261 2091
rect 4295 2088 4307 2091
rect 4798 2088 4804 2100
rect 4295 2060 4804 2088
rect 4295 2057 4307 2060
rect 4249 2051 4307 2057
rect 4798 2048 4804 2060
rect 4856 2048 4862 2100
rect 5166 2048 5172 2100
rect 5224 2097 5230 2100
rect 5224 2091 5243 2097
rect 5231 2057 5243 2091
rect 5224 2051 5243 2057
rect 5353 2091 5411 2097
rect 5353 2057 5365 2091
rect 5399 2088 5411 2091
rect 5399 2060 8156 2088
rect 5399 2057 5411 2060
rect 5353 2051 5411 2057
rect 5224 2048 5230 2051
rect 1946 1980 1952 2032
rect 2004 1980 2010 2032
rect 2682 1980 2688 2032
rect 2740 2020 2746 2032
rect 2961 2023 3019 2029
rect 2961 2020 2973 2023
rect 2740 1992 2973 2020
rect 2740 1980 2746 1992
rect 2961 1989 2973 1992
rect 3007 1989 3019 2023
rect 2961 1983 3019 1989
rect 4985 2023 5043 2029
rect 4985 1989 4997 2023
rect 5031 2020 5043 2023
rect 5442 2020 5448 2032
rect 5031 1992 5448 2020
rect 5031 1989 5043 1992
rect 4985 1983 5043 1989
rect 5442 1980 5448 1992
rect 5500 1980 5506 2032
rect 6549 2023 6607 2029
rect 6549 2020 6561 2023
rect 5552 1992 6561 2020
rect 3234 1912 3240 1964
rect 3292 1912 3298 1964
rect 3326 1912 3332 1964
rect 3384 1952 3390 1964
rect 3789 1955 3847 1961
rect 3789 1952 3801 1955
rect 3384 1924 3801 1952
rect 3384 1912 3390 1924
rect 3789 1921 3801 1924
rect 3835 1921 3847 1955
rect 3789 1915 3847 1921
rect 4709 1955 4767 1961
rect 4709 1921 4721 1955
rect 4755 1952 4767 1955
rect 5074 1952 5080 1964
rect 4755 1924 5080 1952
rect 4755 1921 4767 1924
rect 4709 1915 4767 1921
rect 5074 1912 5080 1924
rect 5132 1912 5138 1964
rect 2314 1844 2320 1896
rect 2372 1884 2378 1896
rect 3513 1887 3571 1893
rect 3513 1884 3525 1887
rect 2372 1856 3525 1884
rect 2372 1844 2378 1856
rect 3513 1853 3525 1856
rect 3559 1884 3571 1887
rect 5552 1884 5580 1992
rect 6549 1989 6561 1992
rect 6595 1989 6607 2023
rect 6549 1983 6607 1989
rect 6730 1980 6736 2032
rect 6788 1980 6794 2032
rect 7558 1980 7564 2032
rect 7616 2020 7622 2032
rect 8021 2023 8079 2029
rect 8021 2020 8033 2023
rect 7616 1992 8033 2020
rect 7616 1980 7622 1992
rect 8021 1989 8033 1992
rect 8067 1989 8079 2023
rect 8128 2020 8156 2060
rect 9030 2048 9036 2100
rect 9088 2088 9094 2100
rect 10134 2088 10140 2100
rect 9088 2060 10140 2088
rect 9088 2048 9094 2060
rect 10134 2048 10140 2060
rect 10192 2048 10198 2100
rect 11149 2091 11207 2097
rect 11149 2057 11161 2091
rect 11195 2088 11207 2091
rect 11606 2088 11612 2100
rect 11195 2060 11612 2088
rect 11195 2057 11207 2060
rect 11149 2051 11207 2057
rect 11606 2048 11612 2060
rect 11664 2048 11670 2100
rect 11974 2048 11980 2100
rect 12032 2088 12038 2100
rect 12032 2060 12112 2088
rect 12032 2048 12038 2060
rect 8128 1992 8510 2020
rect 8021 1983 8079 1989
rect 9674 1980 9680 2032
rect 9732 2020 9738 2032
rect 12084 2020 12112 2060
rect 14090 2048 14096 2100
rect 14148 2088 14154 2100
rect 14829 2091 14887 2097
rect 14829 2088 14841 2091
rect 14148 2060 14841 2088
rect 14148 2048 14154 2060
rect 14829 2057 14841 2060
rect 14875 2057 14887 2091
rect 17862 2088 17868 2100
rect 14829 2051 14887 2057
rect 15120 2060 17868 2088
rect 12161 2023 12219 2029
rect 12161 2020 12173 2023
rect 9732 1992 12020 2020
rect 12084 1992 12173 2020
rect 9732 1980 9738 1992
rect 6457 1955 6515 1961
rect 6457 1952 6469 1955
rect 5736 1924 6469 1952
rect 3559 1856 5580 1884
rect 3559 1853 3571 1856
rect 3513 1847 3571 1853
rect 5626 1844 5632 1896
rect 5684 1844 5690 1896
rect 3878 1776 3884 1828
rect 3936 1816 3942 1828
rect 4341 1819 4399 1825
rect 4341 1816 4353 1819
rect 3936 1788 4353 1816
rect 3936 1776 3942 1788
rect 4341 1785 4353 1788
rect 4387 1785 4399 1819
rect 5736 1816 5764 1924
rect 6457 1921 6469 1924
rect 6503 1921 6515 1955
rect 6457 1915 6515 1921
rect 7374 1912 7380 1964
rect 7432 1912 7438 1964
rect 9582 1912 9588 1964
rect 9640 1952 9646 1964
rect 9769 1955 9827 1961
rect 9769 1952 9781 1955
rect 9640 1924 9781 1952
rect 9640 1912 9646 1924
rect 9769 1921 9781 1924
rect 9815 1921 9827 1955
rect 9769 1915 9827 1921
rect 6012 1856 6868 1884
rect 6012 1825 6040 1856
rect 4341 1779 4399 1785
rect 4448 1788 5764 1816
rect 5997 1819 6055 1825
rect 3142 1708 3148 1760
rect 3200 1748 3206 1760
rect 3602 1748 3608 1760
rect 3200 1720 3608 1748
rect 3200 1708 3206 1720
rect 3602 1708 3608 1720
rect 3660 1748 3666 1760
rect 4448 1748 4476 1788
rect 5997 1785 6009 1819
rect 6043 1785 6055 1819
rect 5997 1779 6055 1785
rect 6730 1776 6736 1828
rect 6788 1776 6794 1828
rect 6840 1816 6868 1856
rect 7098 1844 7104 1896
rect 7156 1884 7162 1896
rect 7745 1887 7803 1893
rect 7745 1884 7757 1887
rect 7156 1856 7757 1884
rect 7156 1844 7162 1856
rect 7745 1853 7757 1856
rect 7791 1853 7803 1887
rect 7745 1847 7803 1853
rect 8110 1844 8116 1896
rect 8168 1884 8174 1896
rect 9674 1884 9680 1896
rect 8168 1856 9680 1884
rect 8168 1844 8174 1856
rect 9674 1844 9680 1856
rect 9732 1844 9738 1896
rect 9784 1884 9812 1915
rect 10042 1912 10048 1964
rect 10100 1912 10106 1964
rect 10199 1955 10257 1961
rect 10199 1921 10211 1955
rect 10245 1952 10257 1955
rect 11054 1952 11060 1964
rect 10245 1924 11060 1952
rect 10245 1921 10257 1924
rect 10199 1915 10257 1921
rect 11054 1912 11060 1924
rect 11112 1912 11118 1964
rect 11146 1912 11152 1964
rect 11204 1952 11210 1964
rect 11992 1961 12020 1992
rect 12161 1989 12173 1992
rect 12207 2020 12219 2023
rect 14981 2023 15039 2029
rect 14981 2020 14993 2023
rect 12207 1992 12756 2020
rect 12207 1989 12219 1992
rect 12161 1983 12219 1989
rect 11977 1955 12035 1961
rect 11204 1924 11928 1952
rect 11204 1912 11210 1924
rect 10689 1887 10747 1893
rect 10689 1884 10701 1887
rect 9784 1856 10701 1884
rect 10689 1853 10701 1856
rect 10735 1853 10747 1887
rect 11900 1884 11928 1924
rect 11977 1921 11989 1955
rect 12023 1921 12035 1955
rect 11977 1915 12035 1921
rect 12066 1912 12072 1964
rect 12124 1952 12130 1964
rect 12728 1961 12756 1992
rect 13464 1992 14993 2020
rect 12345 1955 12403 1961
rect 12345 1952 12357 1955
rect 12124 1924 12357 1952
rect 12124 1912 12130 1924
rect 12345 1921 12357 1924
rect 12391 1921 12403 1955
rect 12345 1915 12403 1921
rect 12713 1955 12771 1961
rect 12713 1921 12725 1955
rect 12759 1921 12771 1955
rect 12713 1915 12771 1921
rect 12805 1887 12863 1893
rect 12805 1884 12817 1887
rect 11900 1856 12817 1884
rect 10689 1847 10747 1853
rect 12805 1853 12817 1856
rect 12851 1853 12863 1887
rect 12805 1847 12863 1853
rect 7466 1816 7472 1828
rect 6840 1788 7472 1816
rect 7466 1776 7472 1788
rect 7524 1776 7530 1828
rect 9048 1788 11928 1816
rect 3660 1720 4476 1748
rect 3660 1708 3666 1720
rect 5166 1708 5172 1760
rect 5224 1708 5230 1760
rect 6089 1751 6147 1757
rect 6089 1717 6101 1751
rect 6135 1748 6147 1751
rect 7006 1748 7012 1760
rect 6135 1720 7012 1748
rect 6135 1717 6147 1720
rect 6089 1711 6147 1717
rect 7006 1708 7012 1720
rect 7064 1708 7070 1760
rect 7098 1708 7104 1760
rect 7156 1748 7162 1760
rect 7285 1751 7343 1757
rect 7285 1748 7297 1751
rect 7156 1720 7297 1748
rect 7156 1708 7162 1720
rect 7285 1717 7297 1720
rect 7331 1748 7343 1751
rect 9048 1748 9076 1788
rect 7331 1720 9076 1748
rect 7331 1717 7343 1720
rect 7285 1711 7343 1717
rect 9674 1708 9680 1760
rect 9732 1748 9738 1760
rect 9950 1748 9956 1760
rect 9732 1720 9956 1748
rect 9732 1708 9738 1720
rect 9950 1708 9956 1720
rect 10008 1708 10014 1760
rect 10229 1751 10287 1757
rect 10229 1717 10241 1751
rect 10275 1748 10287 1751
rect 11790 1748 11796 1760
rect 10275 1720 11796 1748
rect 10275 1717 10287 1720
rect 10229 1711 10287 1717
rect 11790 1708 11796 1720
rect 11848 1708 11854 1760
rect 11900 1748 11928 1788
rect 12066 1776 12072 1828
rect 12124 1816 12130 1828
rect 13262 1816 13268 1828
rect 12124 1788 13268 1816
rect 12124 1776 12130 1788
rect 13262 1776 13268 1788
rect 13320 1776 13326 1828
rect 13464 1748 13492 1992
rect 14981 1989 14993 1992
rect 15027 1989 15039 2023
rect 14981 1983 15039 1989
rect 13538 1912 13544 1964
rect 13596 1912 13602 1964
rect 13630 1912 13636 1964
rect 13688 1912 13694 1964
rect 14185 1955 14243 1961
rect 14185 1921 14197 1955
rect 14231 1952 14243 1955
rect 14274 1952 14280 1964
rect 14231 1924 14280 1952
rect 14231 1921 14243 1924
rect 14185 1915 14243 1921
rect 14274 1912 14280 1924
rect 14332 1912 14338 1964
rect 14553 1955 14611 1961
rect 14553 1921 14565 1955
rect 14599 1952 14611 1955
rect 14734 1952 14740 1964
rect 14599 1924 14740 1952
rect 14599 1921 14611 1924
rect 14553 1915 14611 1921
rect 14734 1912 14740 1924
rect 14792 1912 14798 1964
rect 13556 1884 13584 1912
rect 15120 1884 15148 2060
rect 17862 2048 17868 2060
rect 17920 2048 17926 2100
rect 18690 2048 18696 2100
rect 18748 2088 18754 2100
rect 18877 2091 18935 2097
rect 18877 2088 18889 2091
rect 18748 2060 18889 2088
rect 18748 2048 18754 2060
rect 18877 2057 18889 2060
rect 18923 2057 18935 2091
rect 18877 2051 18935 2057
rect 19058 2048 19064 2100
rect 19116 2088 19122 2100
rect 21377 2091 21435 2097
rect 21377 2088 21389 2091
rect 19116 2060 21389 2088
rect 19116 2048 19122 2060
rect 21377 2057 21389 2060
rect 21423 2088 21435 2091
rect 21545 2091 21603 2097
rect 21423 2060 21496 2088
rect 21423 2057 21435 2060
rect 21377 2051 21435 2057
rect 15197 2023 15255 2029
rect 15197 1989 15209 2023
rect 15243 2020 15255 2023
rect 15470 2020 15476 2032
rect 15243 1992 15476 2020
rect 15243 1989 15255 1992
rect 15197 1983 15255 1989
rect 15470 1980 15476 1992
rect 15528 1980 15534 2032
rect 16025 2023 16083 2029
rect 16025 1989 16037 2023
rect 16071 2020 16083 2023
rect 16574 2020 16580 2032
rect 16071 1992 16580 2020
rect 16071 1989 16083 1992
rect 16025 1983 16083 1989
rect 16574 1980 16580 1992
rect 16632 1980 16638 2032
rect 17034 1980 17040 2032
rect 17092 1980 17098 2032
rect 17494 1980 17500 2032
rect 17552 1980 17558 2032
rect 18414 1980 18420 2032
rect 18472 2020 18478 2032
rect 18472 1992 19182 2020
rect 18472 1980 18478 1992
rect 20714 1980 20720 2032
rect 20772 2020 20778 2032
rect 21177 2023 21235 2029
rect 21177 2020 21189 2023
rect 20772 1992 21189 2020
rect 20772 1980 20778 1992
rect 21177 1989 21189 1992
rect 21223 1989 21235 2023
rect 21177 1983 21235 1989
rect 15562 1912 15568 1964
rect 15620 1952 15626 1964
rect 16301 1955 16359 1961
rect 16301 1952 16313 1955
rect 15620 1924 16313 1952
rect 15620 1912 15626 1924
rect 16301 1921 16313 1924
rect 16347 1921 16359 1955
rect 16301 1915 16359 1921
rect 13556 1856 15148 1884
rect 16316 1884 16344 1915
rect 16758 1912 16764 1964
rect 16816 1912 16822 1964
rect 18782 1884 18788 1896
rect 16316 1856 18788 1884
rect 18782 1844 18788 1856
rect 18840 1844 18846 1896
rect 19886 1884 19892 1896
rect 18892 1856 19892 1884
rect 13630 1776 13636 1828
rect 13688 1816 13694 1828
rect 15194 1816 15200 1828
rect 13688 1788 15200 1816
rect 13688 1776 13694 1788
rect 15194 1776 15200 1788
rect 15252 1776 15258 1828
rect 18138 1776 18144 1828
rect 18196 1816 18202 1828
rect 18509 1819 18567 1825
rect 18509 1816 18521 1819
rect 18196 1788 18521 1816
rect 18196 1776 18202 1788
rect 18509 1785 18521 1788
rect 18555 1785 18567 1819
rect 18509 1779 18567 1785
rect 11900 1720 13492 1748
rect 13814 1708 13820 1760
rect 13872 1748 13878 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 13872 1720 15025 1748
rect 13872 1708 13878 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15930 1708 15936 1760
rect 15988 1748 15994 1760
rect 18892 1748 18920 1856
rect 19886 1844 19892 1856
rect 19944 1844 19950 1896
rect 19978 1844 19984 1896
rect 20036 1884 20042 1896
rect 20349 1887 20407 1893
rect 20349 1884 20361 1887
rect 20036 1856 20361 1884
rect 20036 1844 20042 1856
rect 20349 1853 20361 1856
rect 20395 1853 20407 1887
rect 20349 1847 20407 1853
rect 20625 1887 20683 1893
rect 20625 1853 20637 1887
rect 20671 1853 20683 1887
rect 21468 1884 21496 2060
rect 21545 2057 21557 2091
rect 21591 2088 21603 2091
rect 21591 2060 22094 2088
rect 21591 2057 21603 2060
rect 21545 2051 21603 2057
rect 22066 2020 22094 2060
rect 23658 2048 23664 2100
rect 23716 2088 23722 2100
rect 24029 2091 24087 2097
rect 24029 2088 24041 2091
rect 23716 2060 24041 2088
rect 23716 2048 23722 2060
rect 24029 2057 24041 2060
rect 24075 2057 24087 2091
rect 24762 2088 24768 2100
rect 24029 2051 24087 2057
rect 24320 2060 24768 2088
rect 23477 2023 23535 2029
rect 22066 1992 22310 2020
rect 23477 1989 23489 2023
rect 23523 2020 23535 2023
rect 23842 2020 23848 2032
rect 23523 1992 23848 2020
rect 23523 1989 23535 1992
rect 23477 1983 23535 1989
rect 23842 1980 23848 1992
rect 23900 1980 23906 2032
rect 24192 2023 24250 2029
rect 24192 2020 24204 2023
rect 24136 1992 24204 2020
rect 23750 1912 23756 1964
rect 23808 1912 23814 1964
rect 22094 1884 22100 1896
rect 21468 1856 22100 1884
rect 20625 1847 20683 1853
rect 15988 1720 18920 1748
rect 15988 1708 15994 1720
rect 19794 1708 19800 1760
rect 19852 1748 19858 1760
rect 20640 1748 20668 1847
rect 22094 1844 22100 1856
rect 22152 1884 22158 1896
rect 24136 1884 24164 1992
rect 24192 1989 24204 1992
rect 24238 2020 24250 2023
rect 24320 2020 24348 2060
rect 24762 2048 24768 2060
rect 24820 2048 24826 2100
rect 24238 1992 24348 2020
rect 24397 2023 24455 2029
rect 24238 1989 24250 1992
rect 24192 1983 24250 1989
rect 24397 1989 24409 2023
rect 24443 2020 24455 2023
rect 24670 2020 24676 2032
rect 24443 1992 24676 2020
rect 24443 1989 24455 1992
rect 24397 1983 24455 1989
rect 24670 1980 24676 1992
rect 24728 1980 24734 2032
rect 22152 1856 24164 1884
rect 22152 1844 22158 1856
rect 19852 1720 20668 1748
rect 19852 1708 19858 1720
rect 20806 1708 20812 1760
rect 20864 1748 20870 1760
rect 21361 1751 21419 1757
rect 21361 1748 21373 1751
rect 20864 1720 21373 1748
rect 20864 1708 20870 1720
rect 21361 1717 21373 1720
rect 21407 1717 21419 1751
rect 21361 1711 21419 1717
rect 22002 1708 22008 1760
rect 22060 1708 22066 1760
rect 23934 1708 23940 1760
rect 23992 1748 23998 1760
rect 24213 1751 24271 1757
rect 24213 1748 24225 1751
rect 23992 1720 24225 1748
rect 23992 1708 23998 1720
rect 24213 1717 24225 1720
rect 24259 1717 24271 1751
rect 24213 1711 24271 1717
rect 1104 1658 24840 1680
rect 1104 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 20214 1658
rect 20266 1606 20278 1658
rect 20330 1606 20342 1658
rect 20394 1606 20406 1658
rect 20458 1606 20470 1658
rect 20522 1606 24840 1658
rect 1104 1584 24840 1606
rect 1946 1504 1952 1556
rect 2004 1504 2010 1556
rect 2133 1547 2191 1553
rect 2133 1513 2145 1547
rect 2179 1544 2191 1547
rect 2222 1544 2228 1556
rect 2179 1516 2228 1544
rect 2179 1513 2191 1516
rect 2133 1507 2191 1513
rect 2222 1504 2228 1516
rect 2280 1544 2286 1556
rect 5166 1544 5172 1556
rect 2280 1516 5172 1544
rect 2280 1504 2286 1516
rect 5166 1504 5172 1516
rect 5224 1504 5230 1556
rect 6089 1547 6147 1553
rect 6089 1513 6101 1547
rect 6135 1544 6147 1547
rect 7282 1544 7288 1556
rect 6135 1516 7288 1544
rect 6135 1513 6147 1516
rect 6089 1507 6147 1513
rect 7282 1504 7288 1516
rect 7340 1504 7346 1556
rect 7466 1504 7472 1556
rect 7524 1544 7530 1556
rect 7834 1544 7840 1556
rect 7524 1516 7840 1544
rect 7524 1504 7530 1516
rect 7834 1504 7840 1516
rect 7892 1544 7898 1556
rect 8662 1544 8668 1556
rect 7892 1516 8668 1544
rect 7892 1504 7898 1516
rect 8662 1504 8668 1516
rect 8720 1504 8726 1556
rect 9490 1504 9496 1556
rect 9548 1544 9554 1556
rect 10686 1544 10692 1556
rect 9548 1516 10692 1544
rect 9548 1504 9554 1516
rect 10686 1504 10692 1516
rect 10744 1504 10750 1556
rect 10778 1504 10784 1556
rect 10836 1504 10842 1556
rect 15930 1544 15936 1556
rect 10888 1516 15936 1544
rect 3050 1436 3056 1488
rect 3108 1436 3114 1488
rect 3326 1436 3332 1488
rect 3384 1476 3390 1488
rect 7190 1476 7196 1488
rect 3384 1448 3832 1476
rect 3384 1436 3390 1448
rect 1578 1368 1584 1420
rect 1636 1408 1642 1420
rect 1636 1380 3310 1408
rect 1636 1368 1642 1380
rect 1486 1300 1492 1352
rect 1544 1300 1550 1352
rect 1670 1300 1676 1352
rect 1728 1340 1734 1352
rect 3282 1349 3310 1380
rect 2777 1343 2835 1349
rect 1728 1312 2360 1340
rect 1728 1300 1734 1312
rect 2130 1281 2136 1284
rect 2117 1275 2136 1281
rect 2117 1241 2129 1275
rect 2117 1235 2136 1241
rect 2130 1232 2136 1235
rect 2188 1232 2194 1284
rect 2332 1281 2360 1312
rect 2777 1309 2789 1343
rect 2823 1309 2835 1343
rect 2777 1303 2835 1309
rect 3267 1343 3325 1349
rect 3267 1309 3279 1343
rect 3313 1309 3325 1343
rect 3267 1303 3325 1309
rect 3421 1343 3479 1349
rect 3421 1309 3433 1343
rect 3467 1340 3479 1343
rect 3602 1340 3608 1352
rect 3467 1312 3608 1340
rect 3467 1309 3479 1312
rect 3421 1303 3479 1309
rect 2317 1275 2375 1281
rect 2317 1241 2329 1275
rect 2363 1241 2375 1275
rect 2792 1272 2820 1303
rect 3602 1300 3608 1312
rect 3660 1300 3666 1352
rect 3804 1272 3832 1448
rect 5368 1448 7196 1476
rect 3878 1368 3884 1420
rect 3936 1408 3942 1420
rect 3936 1380 4292 1408
rect 3936 1368 3942 1380
rect 4062 1300 4068 1352
rect 4120 1349 4126 1352
rect 4264 1349 4292 1380
rect 4614 1368 4620 1420
rect 4672 1408 4678 1420
rect 4985 1411 5043 1417
rect 4985 1408 4997 1411
rect 4672 1380 4997 1408
rect 4672 1368 4678 1380
rect 4985 1377 4997 1380
rect 5031 1377 5043 1411
rect 4985 1371 5043 1377
rect 4120 1343 4169 1349
rect 4120 1309 4123 1343
rect 4157 1309 4169 1343
rect 4120 1303 4169 1309
rect 4249 1343 4307 1349
rect 4249 1309 4261 1343
rect 4295 1309 4307 1343
rect 4249 1303 4307 1309
rect 4525 1343 4583 1349
rect 4525 1309 4537 1343
rect 4571 1340 4583 1343
rect 4798 1340 4804 1352
rect 4571 1312 4804 1340
rect 4571 1309 4583 1312
rect 4525 1303 4583 1309
rect 4120 1300 4126 1303
rect 4798 1300 4804 1312
rect 4856 1300 4862 1352
rect 5166 1300 5172 1352
rect 5224 1300 5230 1352
rect 5368 1349 5396 1448
rect 7190 1436 7196 1448
rect 7248 1436 7254 1488
rect 7374 1436 7380 1488
rect 7432 1476 7438 1488
rect 10888 1476 10916 1516
rect 15930 1504 15936 1516
rect 15988 1504 15994 1556
rect 17037 1547 17095 1553
rect 17037 1513 17049 1547
rect 17083 1544 17095 1547
rect 17126 1544 17132 1556
rect 17083 1516 17132 1544
rect 17083 1513 17095 1516
rect 17037 1507 17095 1513
rect 17126 1504 17132 1516
rect 17184 1504 17190 1556
rect 17221 1547 17279 1553
rect 17221 1513 17233 1547
rect 17267 1544 17279 1547
rect 17402 1544 17408 1556
rect 17267 1516 17408 1544
rect 17267 1513 17279 1516
rect 17221 1507 17279 1513
rect 17402 1504 17408 1516
rect 17460 1504 17466 1556
rect 17497 1547 17555 1553
rect 17497 1513 17509 1547
rect 17543 1544 17555 1547
rect 17586 1544 17592 1556
rect 17543 1516 17592 1544
rect 17543 1513 17555 1516
rect 17497 1507 17555 1513
rect 17586 1504 17592 1516
rect 17644 1504 17650 1556
rect 18141 1547 18199 1553
rect 18141 1513 18153 1547
rect 18187 1544 18199 1547
rect 18230 1544 18236 1556
rect 18187 1516 18236 1544
rect 18187 1513 18199 1516
rect 18141 1507 18199 1513
rect 18230 1504 18236 1516
rect 18288 1504 18294 1556
rect 18782 1504 18788 1556
rect 18840 1504 18846 1556
rect 20070 1553 20076 1556
rect 20060 1547 20076 1553
rect 20060 1513 20072 1547
rect 20060 1507 20076 1513
rect 20070 1504 20076 1507
rect 20128 1504 20134 1556
rect 21082 1504 21088 1556
rect 21140 1544 21146 1556
rect 21545 1547 21603 1553
rect 21545 1544 21557 1547
rect 21140 1516 21557 1544
rect 21140 1504 21146 1516
rect 21545 1513 21557 1516
rect 21591 1513 21603 1547
rect 21545 1507 21603 1513
rect 21910 1504 21916 1556
rect 21968 1504 21974 1556
rect 22002 1504 22008 1556
rect 22060 1544 22066 1556
rect 23857 1547 23915 1553
rect 23857 1544 23869 1547
rect 22060 1516 23869 1544
rect 22060 1504 22066 1516
rect 23857 1513 23869 1516
rect 23903 1513 23915 1547
rect 23857 1507 23915 1513
rect 7432 1448 10916 1476
rect 11793 1479 11851 1485
rect 7432 1436 7438 1448
rect 11793 1445 11805 1479
rect 11839 1476 11851 1479
rect 11974 1476 11980 1488
rect 11839 1448 11980 1476
rect 11839 1445 11851 1448
rect 11793 1439 11851 1445
rect 11974 1436 11980 1448
rect 12032 1436 12038 1488
rect 12066 1436 12072 1488
rect 12124 1476 12130 1488
rect 12161 1479 12219 1485
rect 12161 1476 12173 1479
rect 12124 1448 12173 1476
rect 12124 1436 12130 1448
rect 12161 1445 12173 1448
rect 12207 1445 12219 1479
rect 12161 1439 12219 1445
rect 16022 1436 16028 1488
rect 16080 1476 16086 1488
rect 19429 1479 19487 1485
rect 19429 1476 19441 1479
rect 16080 1448 19441 1476
rect 16080 1436 16086 1448
rect 19429 1445 19441 1448
rect 19475 1445 19487 1479
rect 19429 1439 19487 1445
rect 19720 1448 19932 1476
rect 6822 1408 6828 1420
rect 5552 1380 5764 1408
rect 5353 1343 5411 1349
rect 5353 1309 5365 1343
rect 5399 1309 5411 1343
rect 5353 1303 5411 1309
rect 3881 1275 3939 1281
rect 3881 1272 3893 1275
rect 2792 1244 3740 1272
rect 3804 1244 3893 1272
rect 2317 1235 2375 1241
rect 1670 1164 1676 1216
rect 1728 1164 1734 1216
rect 2685 1207 2743 1213
rect 2685 1173 2697 1207
rect 2731 1204 2743 1207
rect 3602 1204 3608 1216
rect 2731 1176 3608 1204
rect 2731 1173 2743 1176
rect 2685 1167 2743 1173
rect 3602 1164 3608 1176
rect 3660 1164 3666 1216
rect 3712 1204 3740 1244
rect 3881 1241 3893 1244
rect 3927 1241 3939 1275
rect 3881 1235 3939 1241
rect 3970 1232 3976 1284
rect 4028 1272 4034 1284
rect 5552 1272 5580 1380
rect 5736 1349 5764 1380
rect 5920 1380 6828 1408
rect 5920 1349 5948 1380
rect 6822 1368 6828 1380
rect 6880 1408 6886 1420
rect 7101 1411 7159 1417
rect 7101 1408 7113 1411
rect 6880 1380 7113 1408
rect 6880 1368 6886 1380
rect 7101 1377 7113 1380
rect 7147 1377 7159 1411
rect 7101 1371 7159 1377
rect 7926 1368 7932 1420
rect 7984 1408 7990 1420
rect 10870 1408 10876 1420
rect 7984 1380 10876 1408
rect 7984 1368 7990 1380
rect 5629 1343 5687 1349
rect 5629 1309 5641 1343
rect 5675 1309 5687 1343
rect 5629 1303 5687 1309
rect 5721 1343 5779 1349
rect 5721 1309 5733 1343
rect 5767 1309 5779 1343
rect 5721 1303 5779 1309
rect 5905 1343 5963 1349
rect 5905 1309 5917 1343
rect 5951 1309 5963 1343
rect 5905 1303 5963 1309
rect 4028 1244 5580 1272
rect 5644 1272 5672 1303
rect 6086 1300 6092 1352
rect 6144 1340 6150 1352
rect 6362 1340 6368 1352
rect 6144 1312 6368 1340
rect 6144 1300 6150 1312
rect 6362 1300 6368 1312
rect 6420 1340 6426 1352
rect 6457 1343 6515 1349
rect 6457 1340 6469 1343
rect 6420 1312 6469 1340
rect 6420 1300 6426 1312
rect 6457 1309 6469 1312
rect 6503 1309 6515 1343
rect 6457 1303 6515 1309
rect 6917 1343 6975 1349
rect 6917 1309 6929 1343
rect 6963 1309 6975 1343
rect 6917 1303 6975 1309
rect 5994 1272 6000 1284
rect 5644 1244 6000 1272
rect 4028 1232 4034 1244
rect 5994 1232 6000 1244
rect 6052 1232 6058 1284
rect 6932 1272 6960 1303
rect 7834 1300 7840 1352
rect 7892 1300 7898 1352
rect 9401 1343 9459 1349
rect 9401 1309 9413 1343
rect 9447 1340 9459 1343
rect 9582 1340 9588 1352
rect 9447 1312 9588 1340
rect 9447 1309 9459 1312
rect 9401 1303 9459 1309
rect 9582 1300 9588 1312
rect 9640 1300 9646 1352
rect 9950 1300 9956 1352
rect 10008 1300 10014 1352
rect 10428 1349 10456 1380
rect 10870 1368 10876 1380
rect 10928 1368 10934 1420
rect 13170 1368 13176 1420
rect 13228 1368 13234 1420
rect 14461 1411 14519 1417
rect 14461 1377 14473 1411
rect 14507 1408 14519 1411
rect 14734 1408 14740 1420
rect 14507 1380 14740 1408
rect 14507 1377 14519 1380
rect 14461 1371 14519 1377
rect 14734 1368 14740 1380
rect 14792 1368 14798 1420
rect 15194 1368 15200 1420
rect 15252 1408 15258 1420
rect 17402 1408 17408 1420
rect 15252 1380 17408 1408
rect 15252 1368 15258 1380
rect 17402 1368 17408 1380
rect 17460 1368 17466 1420
rect 17604 1380 19472 1408
rect 10413 1343 10471 1349
rect 10413 1309 10425 1343
rect 10459 1309 10471 1343
rect 10413 1303 10471 1309
rect 11054 1300 11060 1352
rect 11112 1300 11118 1352
rect 11514 1300 11520 1352
rect 11572 1340 11578 1352
rect 11609 1343 11667 1349
rect 11609 1340 11621 1343
rect 11572 1312 11621 1340
rect 11572 1300 11578 1312
rect 11609 1309 11621 1312
rect 11655 1340 11667 1343
rect 11882 1340 11888 1352
rect 11655 1312 11888 1340
rect 11655 1309 11667 1312
rect 11609 1303 11667 1309
rect 11882 1300 11888 1312
rect 11940 1300 11946 1352
rect 11974 1300 11980 1352
rect 12032 1340 12038 1352
rect 12069 1343 12127 1349
rect 12069 1340 12081 1343
rect 12032 1312 12081 1340
rect 12032 1300 12038 1312
rect 12069 1309 12081 1312
rect 12115 1309 12127 1343
rect 12069 1303 12127 1309
rect 12529 1343 12587 1349
rect 12529 1309 12541 1343
rect 12575 1340 12587 1343
rect 12618 1340 12624 1352
rect 12575 1312 12624 1340
rect 12575 1309 12587 1312
rect 12529 1303 12587 1309
rect 12618 1300 12624 1312
rect 12676 1300 12682 1352
rect 12710 1300 12716 1352
rect 12768 1340 12774 1352
rect 12897 1343 12955 1349
rect 12897 1340 12909 1343
rect 12768 1312 12909 1340
rect 12768 1300 12774 1312
rect 12897 1309 12909 1312
rect 12943 1309 12955 1343
rect 12897 1303 12955 1309
rect 13446 1300 13452 1352
rect 13504 1340 13510 1352
rect 13541 1343 13599 1349
rect 13541 1340 13553 1343
rect 13504 1312 13553 1340
rect 13504 1300 13510 1312
rect 13541 1309 13553 1312
rect 13587 1309 13599 1343
rect 13541 1303 13599 1309
rect 13998 1300 14004 1352
rect 14056 1340 14062 1352
rect 14185 1343 14243 1349
rect 14185 1340 14197 1343
rect 14056 1312 14197 1340
rect 14056 1300 14062 1312
rect 14185 1309 14197 1312
rect 14231 1309 14243 1343
rect 14185 1303 14243 1309
rect 15746 1300 15752 1352
rect 15804 1300 15810 1352
rect 16025 1343 16083 1349
rect 16025 1309 16037 1343
rect 16071 1340 16083 1343
rect 16071 1312 17172 1340
rect 16071 1309 16083 1312
rect 16025 1303 16083 1309
rect 6104 1244 6960 1272
rect 4614 1204 4620 1216
rect 3712 1176 4620 1204
rect 4614 1164 4620 1176
rect 4672 1164 4678 1216
rect 4709 1207 4767 1213
rect 4709 1173 4721 1207
rect 4755 1204 4767 1207
rect 5626 1204 5632 1216
rect 4755 1176 5632 1204
rect 4755 1173 4767 1176
rect 4709 1167 4767 1173
rect 5626 1164 5632 1176
rect 5684 1204 5690 1216
rect 6104 1204 6132 1244
rect 8570 1232 8576 1284
rect 8628 1232 8634 1284
rect 8754 1232 8760 1284
rect 8812 1272 8818 1284
rect 13814 1272 13820 1284
rect 8812 1244 13820 1272
rect 8812 1232 8818 1244
rect 13814 1232 13820 1244
rect 13872 1232 13878 1284
rect 14274 1232 14280 1284
rect 14332 1272 14338 1284
rect 16040 1272 16068 1303
rect 14332 1244 16068 1272
rect 14332 1232 14338 1244
rect 16850 1232 16856 1284
rect 16908 1232 16914 1284
rect 16942 1232 16948 1284
rect 17000 1272 17006 1284
rect 17053 1275 17111 1281
rect 17053 1272 17065 1275
rect 17000 1244 17065 1272
rect 17000 1232 17006 1244
rect 17053 1241 17065 1244
rect 17099 1241 17111 1275
rect 17144 1272 17172 1312
rect 17310 1300 17316 1352
rect 17368 1340 17374 1352
rect 17497 1343 17555 1349
rect 17497 1340 17509 1343
rect 17368 1312 17509 1340
rect 17368 1300 17374 1312
rect 17497 1309 17509 1312
rect 17543 1309 17555 1343
rect 17497 1303 17555 1309
rect 17604 1272 17632 1380
rect 17678 1300 17684 1352
rect 17736 1349 17742 1352
rect 17736 1343 17751 1349
rect 17739 1309 17751 1343
rect 17736 1303 17751 1309
rect 17736 1300 17742 1303
rect 18690 1300 18696 1352
rect 18748 1340 18754 1352
rect 18815 1343 18873 1349
rect 18815 1340 18827 1343
rect 18748 1312 18827 1340
rect 18748 1300 18754 1312
rect 18815 1309 18827 1312
rect 18861 1309 18873 1343
rect 18815 1303 18873 1309
rect 18966 1300 18972 1352
rect 19024 1300 19030 1352
rect 19334 1300 19340 1352
rect 19392 1300 19398 1352
rect 19444 1340 19472 1380
rect 19521 1343 19579 1349
rect 19521 1340 19533 1343
rect 19444 1312 19533 1340
rect 19521 1309 19533 1312
rect 19567 1340 19579 1343
rect 19720 1340 19748 1448
rect 19794 1368 19800 1420
rect 19852 1368 19858 1420
rect 19904 1408 19932 1448
rect 19904 1380 21312 1408
rect 19567 1312 19748 1340
rect 21284 1340 21312 1380
rect 23750 1368 23756 1420
rect 23808 1408 23814 1420
rect 24121 1411 24179 1417
rect 24121 1408 24133 1411
rect 23808 1380 24133 1408
rect 23808 1368 23814 1380
rect 24121 1377 24133 1380
rect 24167 1377 24179 1411
rect 24121 1371 24179 1377
rect 21913 1343 21971 1349
rect 21913 1340 21925 1343
rect 21284 1312 21925 1340
rect 19567 1309 19579 1312
rect 19521 1303 19579 1309
rect 21913 1309 21925 1312
rect 21959 1309 21971 1343
rect 21913 1303 21971 1309
rect 22094 1300 22100 1352
rect 22152 1300 22158 1352
rect 22738 1300 22744 1352
rect 22796 1300 22802 1352
rect 17144 1244 17632 1272
rect 17053 1235 17111 1241
rect 17862 1232 17868 1284
rect 17920 1272 17926 1284
rect 17957 1275 18015 1281
rect 17957 1272 17969 1275
rect 17920 1244 17969 1272
rect 17920 1232 17926 1244
rect 17957 1241 17969 1244
rect 18003 1241 18015 1275
rect 17957 1235 18015 1241
rect 18173 1275 18231 1281
rect 18173 1241 18185 1275
rect 18219 1272 18231 1275
rect 18984 1272 19012 1300
rect 18219 1244 18536 1272
rect 18984 1244 20024 1272
rect 18219 1241 18231 1244
rect 18173 1235 18231 1241
rect 5684 1176 6132 1204
rect 5684 1164 5690 1176
rect 6638 1164 6644 1216
rect 6696 1164 6702 1216
rect 8481 1207 8539 1213
rect 8481 1173 8493 1207
rect 8527 1204 8539 1207
rect 8772 1204 8800 1232
rect 8527 1176 8800 1204
rect 9125 1207 9183 1213
rect 8527 1173 8539 1176
rect 8481 1167 8539 1173
rect 9125 1173 9137 1207
rect 9171 1204 9183 1207
rect 13998 1204 14004 1216
rect 9171 1176 14004 1204
rect 9171 1173 9183 1176
rect 9125 1167 9183 1173
rect 13998 1164 14004 1176
rect 14056 1164 14062 1216
rect 18325 1207 18383 1213
rect 18325 1173 18337 1207
rect 18371 1204 18383 1207
rect 18414 1204 18420 1216
rect 18371 1176 18420 1204
rect 18371 1173 18383 1176
rect 18325 1167 18383 1173
rect 18414 1164 18420 1176
rect 18472 1164 18478 1216
rect 18508 1204 18536 1244
rect 19996 1216 20024 1244
rect 20070 1232 20076 1284
rect 20128 1272 20134 1284
rect 20128 1244 20562 1272
rect 20128 1232 20134 1244
rect 19058 1204 19064 1216
rect 18508 1176 19064 1204
rect 19058 1164 19064 1176
rect 19116 1164 19122 1216
rect 19978 1164 19984 1216
rect 20036 1204 20042 1216
rect 22373 1207 22431 1213
rect 22373 1204 22385 1207
rect 20036 1176 22385 1204
rect 20036 1164 20042 1176
rect 22373 1173 22385 1176
rect 22419 1173 22431 1207
rect 22373 1167 22431 1173
rect 1104 1114 24840 1136
rect 1104 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 24214 1114
rect 24266 1062 24278 1114
rect 24330 1062 24342 1114
rect 24394 1062 24406 1114
rect 24458 1062 24470 1114
rect 24522 1062 24840 1114
rect 1104 1040 24840 1062
rect 1670 960 1676 1012
rect 1728 1000 1734 1012
rect 13078 1000 13084 1012
rect 1728 972 13084 1000
rect 1728 960 1734 972
rect 13078 960 13084 972
rect 13136 960 13142 1012
rect 18506 960 18512 1012
rect 18564 1000 18570 1012
rect 20070 1000 20076 1012
rect 18564 972 20076 1000
rect 18564 960 18570 972
rect 20070 960 20076 972
rect 20128 960 20134 1012
rect 6638 892 6644 944
rect 6696 932 6702 944
rect 13722 932 13728 944
rect 6696 904 13728 932
rect 6696 892 6702 904
rect 13722 892 13728 904
rect 13780 892 13786 944
rect 18230 892 18236 944
rect 18288 932 18294 944
rect 21450 932 21456 944
rect 18288 904 21456 932
rect 18288 892 18294 904
rect 21450 892 21456 904
rect 21508 892 21514 944
rect 22094 932 22100 944
rect 22066 892 22100 932
rect 22152 892 22158 944
rect 4798 824 4804 876
rect 4856 864 4862 876
rect 6454 864 6460 876
rect 4856 836 6460 864
rect 4856 824 4862 836
rect 6454 824 6460 836
rect 6512 864 6518 876
rect 7558 864 7564 876
rect 6512 836 7564 864
rect 6512 824 6518 836
rect 7558 824 7564 836
rect 7616 824 7622 876
rect 8570 824 8576 876
rect 8628 864 8634 876
rect 8628 836 16068 864
rect 8628 824 8634 836
rect 16040 796 16068 836
rect 19334 824 19340 876
rect 19392 864 19398 876
rect 22066 864 22094 892
rect 19392 836 22094 864
rect 19392 824 19398 836
rect 19702 796 19708 808
rect 16040 768 19708 796
rect 19702 756 19708 768
rect 19760 756 19766 808
rect 17678 688 17684 740
rect 17736 728 17742 740
rect 19334 728 19340 740
rect 17736 700 19340 728
rect 17736 688 17742 700
rect 19334 688 19340 700
rect 19392 688 19398 740
<< via1 >>
rect 13820 19252 13872 19304
rect 24400 19252 24452 19304
rect 13360 18640 13412 18692
rect 21456 18640 21508 18692
rect 13176 18572 13228 18624
rect 23480 18572 23532 18624
rect 8214 18470 8266 18522
rect 8278 18470 8330 18522
rect 8342 18470 8394 18522
rect 8406 18470 8458 18522
rect 8470 18470 8522 18522
rect 16214 18470 16266 18522
rect 16278 18470 16330 18522
rect 16342 18470 16394 18522
rect 16406 18470 16458 18522
rect 16470 18470 16522 18522
rect 24214 18470 24266 18522
rect 24278 18470 24330 18522
rect 24342 18470 24394 18522
rect 24406 18470 24458 18522
rect 24470 18470 24522 18522
rect 10876 18368 10928 18420
rect 13360 18411 13412 18420
rect 13360 18377 13369 18411
rect 13369 18377 13403 18411
rect 13403 18377 13412 18411
rect 13360 18368 13412 18377
rect 14188 18368 14240 18420
rect 20628 18368 20680 18420
rect 20904 18368 20956 18420
rect 1860 18300 1912 18352
rect 2412 18300 2464 18352
rect 1308 18232 1360 18284
rect 2964 18275 3016 18284
rect 2964 18241 2973 18275
rect 2973 18241 3007 18275
rect 3007 18241 3016 18275
rect 2964 18232 3016 18241
rect 3884 18232 3936 18284
rect 5264 18275 5316 18284
rect 5264 18241 5273 18275
rect 5273 18241 5307 18275
rect 5307 18241 5316 18275
rect 5264 18232 5316 18241
rect 6460 18232 6512 18284
rect 9680 18300 9732 18352
rect 16948 18343 17000 18352
rect 16948 18309 16957 18343
rect 16957 18309 16991 18343
rect 16991 18309 17000 18343
rect 16948 18300 17000 18309
rect 17500 18300 17552 18352
rect 8852 18232 8904 18284
rect 9036 18232 9088 18284
rect 5356 18207 5408 18216
rect 5356 18173 5365 18207
rect 5365 18173 5399 18207
rect 5399 18173 5408 18207
rect 5356 18164 5408 18173
rect 5448 18207 5500 18216
rect 5448 18173 5457 18207
rect 5457 18173 5491 18207
rect 5491 18173 5500 18207
rect 5448 18164 5500 18173
rect 11520 18164 11572 18216
rect 12716 18232 12768 18284
rect 13176 18275 13228 18284
rect 13176 18241 13185 18275
rect 13185 18241 13219 18275
rect 13219 18241 13228 18275
rect 13176 18232 13228 18241
rect 13820 18232 13872 18284
rect 5172 18096 5224 18148
rect 1676 18071 1728 18080
rect 1676 18037 1685 18071
rect 1685 18037 1719 18071
rect 1719 18037 1728 18071
rect 1676 18028 1728 18037
rect 2504 18071 2556 18080
rect 2504 18037 2513 18071
rect 2513 18037 2547 18071
rect 2547 18037 2556 18071
rect 2504 18028 2556 18037
rect 2596 18028 2648 18080
rect 4620 18028 4672 18080
rect 7932 18028 7984 18080
rect 8576 18028 8628 18080
rect 9312 18071 9364 18080
rect 9312 18037 9321 18071
rect 9321 18037 9355 18071
rect 9355 18037 9364 18071
rect 9312 18028 9364 18037
rect 11152 18071 11204 18080
rect 11152 18037 11161 18071
rect 11161 18037 11195 18071
rect 11195 18037 11204 18071
rect 11152 18028 11204 18037
rect 12072 18139 12124 18148
rect 12072 18105 12081 18139
rect 12081 18105 12115 18139
rect 12115 18105 12124 18139
rect 12072 18096 12124 18105
rect 13912 18096 13964 18148
rect 14280 18139 14332 18148
rect 14280 18105 14289 18139
rect 14289 18105 14323 18139
rect 14323 18105 14332 18139
rect 14280 18096 14332 18105
rect 17408 18275 17460 18284
rect 17408 18241 17417 18275
rect 17417 18241 17451 18275
rect 17451 18241 17460 18275
rect 17408 18232 17460 18241
rect 18696 18232 18748 18284
rect 19340 18300 19392 18352
rect 23664 18300 23716 18352
rect 20812 18232 20864 18284
rect 14556 18164 14608 18216
rect 16120 18164 16172 18216
rect 15292 18139 15344 18148
rect 15292 18105 15301 18139
rect 15301 18105 15335 18139
rect 15335 18105 15344 18139
rect 15292 18096 15344 18105
rect 17868 18207 17920 18216
rect 17868 18173 17877 18207
rect 17877 18173 17911 18207
rect 17911 18173 17920 18207
rect 17868 18164 17920 18173
rect 18420 18207 18472 18216
rect 18420 18173 18429 18207
rect 18429 18173 18463 18207
rect 18463 18173 18472 18207
rect 18420 18164 18472 18173
rect 20904 18207 20956 18216
rect 20904 18173 20913 18207
rect 20913 18173 20947 18207
rect 20947 18173 20956 18207
rect 20904 18164 20956 18173
rect 23480 18275 23532 18284
rect 23480 18241 23489 18275
rect 23489 18241 23523 18275
rect 23523 18241 23532 18275
rect 23480 18232 23532 18241
rect 24124 18275 24176 18284
rect 24124 18241 24133 18275
rect 24133 18241 24167 18275
rect 24167 18241 24176 18275
rect 24124 18232 24176 18241
rect 22468 18207 22520 18216
rect 22468 18173 22477 18207
rect 22477 18173 22511 18207
rect 22511 18173 22520 18207
rect 22468 18164 22520 18173
rect 18328 18096 18380 18148
rect 19984 18096 20036 18148
rect 21824 18096 21876 18148
rect 18788 18071 18840 18080
rect 18788 18037 18797 18071
rect 18797 18037 18831 18071
rect 18831 18037 18840 18071
rect 18788 18028 18840 18037
rect 19432 18028 19484 18080
rect 19800 18071 19852 18080
rect 19800 18037 19809 18071
rect 19809 18037 19843 18071
rect 19843 18037 19852 18071
rect 19800 18028 19852 18037
rect 21640 18028 21692 18080
rect 23204 18028 23256 18080
rect 23388 18071 23440 18080
rect 23388 18037 23397 18071
rect 23397 18037 23431 18071
rect 23431 18037 23440 18071
rect 23388 18028 23440 18037
rect 23756 18028 23808 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 12214 17926 12266 17978
rect 12278 17926 12330 17978
rect 12342 17926 12394 17978
rect 12406 17926 12458 17978
rect 12470 17926 12522 17978
rect 20214 17926 20266 17978
rect 20278 17926 20330 17978
rect 20342 17926 20394 17978
rect 20406 17926 20458 17978
rect 20470 17926 20522 17978
rect 1676 17824 1728 17876
rect 9128 17824 9180 17876
rect 22468 17824 22520 17876
rect 15292 17756 15344 17808
rect 16764 17756 16816 17808
rect 17500 17799 17552 17808
rect 17500 17765 17509 17799
rect 17509 17765 17543 17799
rect 17543 17765 17552 17799
rect 17500 17756 17552 17765
rect 20628 17799 20680 17808
rect 20628 17765 20637 17799
rect 20637 17765 20671 17799
rect 20671 17765 20680 17799
rect 20628 17756 20680 17765
rect 23204 17799 23256 17808
rect 23204 17765 23213 17799
rect 23213 17765 23247 17799
rect 23247 17765 23256 17799
rect 23204 17756 23256 17765
rect 4620 17731 4672 17740
rect 4620 17697 4629 17731
rect 4629 17697 4663 17731
rect 4663 17697 4672 17731
rect 4620 17688 4672 17697
rect 5264 17688 5316 17740
rect 8760 17688 8812 17740
rect 11612 17688 11664 17740
rect 4068 17620 4120 17672
rect 5724 17620 5776 17672
rect 1952 17552 2004 17604
rect 2596 17552 2648 17604
rect 7932 17552 7984 17604
rect 3332 17527 3384 17536
rect 3332 17493 3341 17527
rect 3341 17493 3375 17527
rect 3375 17493 3384 17527
rect 3332 17484 3384 17493
rect 7380 17484 7432 17536
rect 8116 17484 8168 17536
rect 10692 17620 10744 17672
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 14464 17663 14516 17672
rect 14464 17629 14473 17663
rect 14473 17629 14507 17663
rect 14507 17629 14516 17663
rect 14464 17620 14516 17629
rect 16120 17620 16172 17672
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 17408 17688 17460 17740
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 21640 17620 21692 17672
rect 21824 17620 21876 17672
rect 23296 17663 23348 17672
rect 23296 17629 23305 17663
rect 23305 17629 23339 17663
rect 23339 17629 23348 17663
rect 23296 17620 23348 17629
rect 12808 17595 12860 17604
rect 12808 17561 12817 17595
rect 12817 17561 12851 17595
rect 12851 17561 12860 17595
rect 12808 17552 12860 17561
rect 13544 17552 13596 17604
rect 20076 17484 20128 17536
rect 23940 17527 23992 17536
rect 23940 17493 23949 17527
rect 23949 17493 23983 17527
rect 23983 17493 23992 17527
rect 23940 17484 23992 17493
rect 8214 17382 8266 17434
rect 8278 17382 8330 17434
rect 8342 17382 8394 17434
rect 8406 17382 8458 17434
rect 8470 17382 8522 17434
rect 16214 17382 16266 17434
rect 16278 17382 16330 17434
rect 16342 17382 16394 17434
rect 16406 17382 16458 17434
rect 16470 17382 16522 17434
rect 24214 17382 24266 17434
rect 24278 17382 24330 17434
rect 24342 17382 24394 17434
rect 24406 17382 24458 17434
rect 24470 17382 24522 17434
rect 1952 17280 2004 17332
rect 2872 17323 2924 17332
rect 2872 17289 2881 17323
rect 2881 17289 2915 17323
rect 2915 17289 2924 17323
rect 2872 17280 2924 17289
rect 3332 17280 3384 17332
rect 1860 17255 1912 17264
rect 1860 17221 1869 17255
rect 1869 17221 1903 17255
rect 1903 17221 1912 17255
rect 1860 17212 1912 17221
rect 2412 17212 2464 17264
rect 5264 17280 5316 17332
rect 8116 17280 8168 17332
rect 8760 17280 8812 17332
rect 9956 17280 10008 17332
rect 4804 17212 4856 17264
rect 6828 17144 6880 17196
rect 10600 17212 10652 17264
rect 11152 17212 11204 17264
rect 12072 17212 12124 17264
rect 12716 17212 12768 17264
rect 14372 17212 14424 17264
rect 2780 17008 2832 17060
rect 1952 16940 2004 16992
rect 2504 16940 2556 16992
rect 3976 17119 4028 17128
rect 3976 17085 3985 17119
rect 3985 17085 4019 17119
rect 4019 17085 4028 17119
rect 3976 17076 4028 17085
rect 4712 17076 4764 17128
rect 7932 17119 7984 17128
rect 7932 17085 7941 17119
rect 7941 17085 7975 17119
rect 7975 17085 7984 17119
rect 7932 17076 7984 17085
rect 5356 17008 5408 17060
rect 4988 16940 5040 16992
rect 6736 16940 6788 16992
rect 7380 16940 7432 16992
rect 9312 17144 9364 17196
rect 10232 17187 10284 17196
rect 10232 17153 10241 17187
rect 10241 17153 10275 17187
rect 10275 17153 10284 17187
rect 10232 17144 10284 17153
rect 11612 17187 11664 17196
rect 11612 17153 11621 17187
rect 11621 17153 11655 17187
rect 11655 17153 11664 17187
rect 11612 17144 11664 17153
rect 13084 17144 13136 17196
rect 14280 17187 14332 17196
rect 14280 17153 14289 17187
rect 14289 17153 14323 17187
rect 14323 17153 14332 17187
rect 14648 17187 14700 17196
rect 14280 17144 14332 17153
rect 14648 17153 14657 17187
rect 14657 17153 14691 17187
rect 14691 17153 14700 17187
rect 14648 17144 14700 17153
rect 15568 17187 15620 17196
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 18328 17280 18380 17332
rect 24124 17280 24176 17332
rect 24584 17280 24636 17332
rect 18696 17255 18748 17264
rect 18696 17221 18705 17255
rect 18705 17221 18739 17255
rect 18739 17221 18748 17255
rect 18696 17212 18748 17221
rect 20076 17212 20128 17264
rect 8944 17119 8996 17128
rect 8944 17085 8953 17119
rect 8953 17085 8987 17119
rect 8987 17085 8996 17119
rect 8944 17076 8996 17085
rect 9036 17119 9088 17128
rect 9036 17085 9045 17119
rect 9045 17085 9079 17119
rect 9079 17085 9088 17119
rect 9036 17076 9088 17085
rect 10692 17119 10744 17128
rect 10692 17085 10701 17119
rect 10701 17085 10735 17119
rect 10735 17085 10744 17119
rect 10692 17076 10744 17085
rect 12716 17076 12768 17128
rect 13360 17076 13412 17128
rect 11612 17008 11664 17060
rect 13360 16940 13412 16992
rect 13544 17008 13596 17060
rect 15200 17076 15252 17128
rect 18236 17187 18288 17196
rect 18236 17153 18245 17187
rect 18245 17153 18279 17187
rect 18279 17153 18288 17187
rect 18236 17144 18288 17153
rect 20812 17144 20864 17196
rect 21364 17076 21416 17128
rect 19616 17008 19668 17060
rect 23388 17212 23440 17264
rect 22192 17144 22244 17196
rect 23940 17187 23992 17196
rect 23940 17153 23949 17187
rect 23949 17153 23983 17187
rect 23983 17153 23992 17187
rect 23940 17144 23992 17153
rect 22468 17076 22520 17128
rect 22928 17076 22980 17128
rect 22284 17008 22336 17060
rect 23296 17008 23348 17060
rect 20904 16940 20956 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 12214 16838 12266 16890
rect 12278 16838 12330 16890
rect 12342 16838 12394 16890
rect 12406 16838 12458 16890
rect 12470 16838 12522 16890
rect 20214 16838 20266 16890
rect 20278 16838 20330 16890
rect 20342 16838 20394 16890
rect 20406 16838 20458 16890
rect 20470 16838 20522 16890
rect 4068 16600 4120 16652
rect 4712 16779 4764 16788
rect 4712 16745 4721 16779
rect 4721 16745 4755 16779
rect 4755 16745 4764 16779
rect 4712 16736 4764 16745
rect 5724 16779 5776 16788
rect 5724 16745 5733 16779
rect 5733 16745 5767 16779
rect 5767 16745 5776 16779
rect 5724 16736 5776 16745
rect 5908 16779 5960 16788
rect 5908 16745 5917 16779
rect 5917 16745 5951 16779
rect 5951 16745 5960 16779
rect 5908 16736 5960 16745
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7932 16736 7984 16788
rect 4804 16668 4856 16720
rect 8576 16736 8628 16788
rect 11060 16668 11112 16720
rect 4988 16600 5040 16652
rect 5448 16600 5500 16652
rect 7196 16643 7248 16652
rect 7196 16609 7205 16643
rect 7205 16609 7239 16643
rect 7239 16609 7248 16643
rect 7196 16600 7248 16609
rect 7380 16643 7432 16652
rect 7380 16609 7389 16643
rect 7389 16609 7423 16643
rect 7423 16609 7432 16643
rect 7380 16600 7432 16609
rect 13544 16711 13596 16720
rect 13544 16677 13553 16711
rect 13553 16677 13587 16711
rect 13587 16677 13596 16711
rect 13544 16668 13596 16677
rect 15568 16736 15620 16788
rect 16120 16736 16172 16788
rect 17684 16736 17736 16788
rect 18420 16736 18472 16788
rect 18696 16736 18748 16788
rect 19340 16736 19392 16788
rect 20904 16779 20956 16788
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 5356 16532 5408 16584
rect 6736 16532 6788 16584
rect 1768 16507 1820 16516
rect 1768 16473 1777 16507
rect 1777 16473 1811 16507
rect 1811 16473 1820 16507
rect 1768 16464 1820 16473
rect 2780 16464 2832 16516
rect 3056 16464 3108 16516
rect 5724 16464 5776 16516
rect 8024 16464 8076 16516
rect 2688 16396 2740 16448
rect 5080 16396 5132 16448
rect 5356 16396 5408 16448
rect 6000 16396 6052 16448
rect 7104 16396 7156 16448
rect 8852 16464 8904 16516
rect 11060 16532 11112 16584
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 12808 16532 12860 16584
rect 14372 16575 14424 16584
rect 14372 16541 14381 16575
rect 14381 16541 14415 16575
rect 14415 16541 14424 16575
rect 14372 16532 14424 16541
rect 14648 16575 14700 16584
rect 14648 16541 14657 16575
rect 14657 16541 14691 16575
rect 14691 16541 14700 16575
rect 14648 16532 14700 16541
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 15844 16532 15896 16584
rect 16028 16575 16080 16584
rect 16028 16541 16037 16575
rect 16037 16541 16071 16575
rect 16071 16541 16080 16575
rect 16028 16532 16080 16541
rect 16120 16532 16172 16584
rect 17960 16600 18012 16652
rect 8576 16396 8628 16448
rect 12624 16507 12676 16516
rect 12624 16473 12633 16507
rect 12633 16473 12667 16507
rect 12667 16473 12676 16507
rect 12624 16464 12676 16473
rect 15200 16464 15252 16516
rect 15660 16464 15712 16516
rect 17684 16575 17736 16584
rect 17684 16541 17693 16575
rect 17693 16541 17727 16575
rect 17727 16541 17736 16575
rect 17684 16532 17736 16541
rect 18236 16532 18288 16584
rect 23296 16668 23348 16720
rect 18696 16532 18748 16584
rect 19984 16532 20036 16584
rect 18328 16507 18380 16516
rect 18328 16473 18337 16507
rect 18337 16473 18371 16507
rect 18371 16473 18380 16507
rect 18328 16464 18380 16473
rect 19524 16507 19576 16516
rect 19524 16473 19533 16507
rect 19533 16473 19567 16507
rect 19567 16473 19576 16507
rect 19524 16464 19576 16473
rect 16028 16396 16080 16448
rect 17868 16396 17920 16448
rect 17960 16396 18012 16448
rect 19432 16396 19484 16448
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 21088 16575 21140 16584
rect 21088 16541 21097 16575
rect 21097 16541 21131 16575
rect 21131 16541 21140 16575
rect 21088 16532 21140 16541
rect 21180 16575 21232 16584
rect 21180 16541 21189 16575
rect 21189 16541 21223 16575
rect 21223 16541 21232 16575
rect 21180 16532 21232 16541
rect 21548 16532 21600 16584
rect 22376 16532 22428 16584
rect 22468 16575 22520 16584
rect 22468 16541 22477 16575
rect 22477 16541 22511 16575
rect 22511 16541 22520 16575
rect 22468 16532 22520 16541
rect 21272 16507 21324 16516
rect 21272 16473 21281 16507
rect 21281 16473 21315 16507
rect 21315 16473 21324 16507
rect 21272 16464 21324 16473
rect 21732 16464 21784 16516
rect 23572 16464 23624 16516
rect 21180 16396 21232 16448
rect 8214 16294 8266 16346
rect 8278 16294 8330 16346
rect 8342 16294 8394 16346
rect 8406 16294 8458 16346
rect 8470 16294 8522 16346
rect 16214 16294 16266 16346
rect 16278 16294 16330 16346
rect 16342 16294 16394 16346
rect 16406 16294 16458 16346
rect 16470 16294 16522 16346
rect 24214 16294 24266 16346
rect 24278 16294 24330 16346
rect 24342 16294 24394 16346
rect 24406 16294 24458 16346
rect 24470 16294 24522 16346
rect 1768 16192 1820 16244
rect 2688 16235 2740 16244
rect 2688 16201 2697 16235
rect 2697 16201 2731 16235
rect 2731 16201 2740 16235
rect 2688 16192 2740 16201
rect 2872 16192 2924 16244
rect 2136 16124 2188 16176
rect 1492 16099 1544 16108
rect 1492 16065 1501 16099
rect 1501 16065 1535 16099
rect 1535 16065 1544 16099
rect 1492 16056 1544 16065
rect 2872 16056 2924 16108
rect 4988 16192 5040 16244
rect 5080 16192 5132 16244
rect 7104 16192 7156 16244
rect 4068 16124 4120 16176
rect 5264 16056 5316 16108
rect 7104 16056 7156 16108
rect 8116 16192 8168 16244
rect 8944 16235 8996 16244
rect 8944 16201 8953 16235
rect 8953 16201 8987 16235
rect 8987 16201 8996 16235
rect 8944 16192 8996 16201
rect 9680 16124 9732 16176
rect 11060 16235 11112 16244
rect 11060 16201 11069 16235
rect 11069 16201 11103 16235
rect 11103 16201 11112 16235
rect 11060 16192 11112 16201
rect 13820 16192 13872 16244
rect 16028 16192 16080 16244
rect 18420 16192 18472 16244
rect 11152 16124 11204 16176
rect 21272 16192 21324 16244
rect 23664 16192 23716 16244
rect 18972 16124 19024 16176
rect 8576 16056 8628 16108
rect 11612 16099 11664 16108
rect 11612 16065 11621 16099
rect 11621 16065 11655 16099
rect 11655 16065 11664 16099
rect 11612 16056 11664 16065
rect 12624 16099 12676 16108
rect 12624 16065 12633 16099
rect 12633 16065 12667 16099
rect 12667 16065 12676 16099
rect 12624 16056 12676 16065
rect 13268 16056 13320 16108
rect 13728 16099 13780 16108
rect 13728 16065 13737 16099
rect 13737 16065 13771 16099
rect 13771 16065 13780 16099
rect 13728 16056 13780 16065
rect 4620 15988 4672 16040
rect 7932 15988 7984 16040
rect 8024 15988 8076 16040
rect 9680 15988 9732 16040
rect 13360 15988 13412 16040
rect 13912 16099 13964 16108
rect 13912 16065 13926 16099
rect 13926 16065 13960 16099
rect 13960 16065 13964 16099
rect 13912 16056 13964 16065
rect 15108 16056 15160 16108
rect 15476 16056 15528 16108
rect 16580 16056 16632 16108
rect 18236 16056 18288 16108
rect 18604 16056 18656 16108
rect 19524 16056 19576 16108
rect 21732 16124 21784 16176
rect 22284 16124 22336 16176
rect 23480 16167 23532 16176
rect 23480 16133 23489 16167
rect 23489 16133 23523 16167
rect 23523 16133 23532 16167
rect 23480 16124 23532 16133
rect 20720 16056 20772 16108
rect 20996 16056 21048 16108
rect 21180 16099 21232 16108
rect 21180 16065 21189 16099
rect 21189 16065 21223 16099
rect 21223 16065 21232 16099
rect 21180 16056 21232 16065
rect 21456 16056 21508 16108
rect 22192 16099 22244 16108
rect 22192 16065 22201 16099
rect 22201 16065 22235 16099
rect 22235 16065 22244 16099
rect 22192 16056 22244 16065
rect 23112 16099 23164 16108
rect 23112 16065 23121 16099
rect 23121 16065 23155 16099
rect 23155 16065 23164 16099
rect 23112 16056 23164 16065
rect 23204 16056 23256 16108
rect 15844 15988 15896 16040
rect 17040 15988 17092 16040
rect 17316 15988 17368 16040
rect 18788 16031 18840 16040
rect 18788 15997 18797 16031
rect 18797 15997 18831 16031
rect 18831 15997 18840 16031
rect 18788 15988 18840 15997
rect 19340 16031 19392 16040
rect 19340 15997 19349 16031
rect 19349 15997 19383 16031
rect 19383 15997 19392 16031
rect 19340 15988 19392 15997
rect 19892 16031 19944 16040
rect 19892 15997 19901 16031
rect 19901 15997 19935 16031
rect 19935 15997 19944 16031
rect 19892 15988 19944 15997
rect 5356 15920 5408 15972
rect 10324 15920 10376 15972
rect 5448 15852 5500 15904
rect 10140 15852 10192 15904
rect 12900 15963 12952 15972
rect 12900 15929 12909 15963
rect 12909 15929 12943 15963
rect 12943 15929 12952 15963
rect 12900 15920 12952 15929
rect 18696 15920 18748 15972
rect 11980 15852 12032 15904
rect 15568 15895 15620 15904
rect 15568 15861 15577 15895
rect 15577 15861 15611 15895
rect 15611 15861 15620 15895
rect 15568 15852 15620 15861
rect 15660 15852 15712 15904
rect 19800 15920 19852 15972
rect 19984 15895 20036 15904
rect 19984 15861 19993 15895
rect 19993 15861 20027 15895
rect 20027 15861 20036 15895
rect 19984 15852 20036 15861
rect 20996 15852 21048 15904
rect 21180 15852 21232 15904
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 23296 15852 23348 15904
rect 24676 16056 24728 16108
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 12214 15750 12266 15802
rect 12278 15750 12330 15802
rect 12342 15750 12394 15802
rect 12406 15750 12458 15802
rect 12470 15750 12522 15802
rect 20214 15750 20266 15802
rect 20278 15750 20330 15802
rect 20342 15750 20394 15802
rect 20406 15750 20458 15802
rect 20470 15750 20522 15802
rect 4620 15648 4672 15700
rect 5264 15648 5316 15700
rect 5908 15648 5960 15700
rect 7932 15691 7984 15700
rect 7932 15657 7941 15691
rect 7941 15657 7975 15691
rect 7975 15657 7984 15691
rect 7932 15648 7984 15657
rect 14832 15691 14884 15700
rect 14832 15657 14841 15691
rect 14841 15657 14875 15691
rect 14875 15657 14884 15691
rect 14832 15648 14884 15657
rect 15200 15648 15252 15700
rect 2688 15555 2740 15564
rect 2688 15521 2697 15555
rect 2697 15521 2731 15555
rect 2731 15521 2740 15555
rect 2688 15512 2740 15521
rect 4988 15555 5040 15564
rect 4988 15521 4997 15555
rect 4997 15521 5031 15555
rect 5031 15521 5040 15555
rect 4988 15512 5040 15521
rect 5448 15580 5500 15632
rect 13820 15580 13872 15632
rect 15016 15580 15068 15632
rect 16120 15648 16172 15700
rect 7196 15512 7248 15564
rect 8576 15512 8628 15564
rect 9036 15512 9088 15564
rect 11612 15555 11664 15564
rect 11612 15521 11621 15555
rect 11621 15521 11655 15555
rect 11655 15521 11664 15555
rect 11612 15512 11664 15521
rect 11980 15512 12032 15564
rect 15108 15512 15160 15564
rect 5356 15444 5408 15496
rect 6000 15444 6052 15496
rect 6736 15444 6788 15496
rect 8944 15444 8996 15496
rect 10232 15487 10284 15496
rect 10232 15453 10241 15487
rect 10241 15453 10275 15487
rect 10275 15453 10284 15487
rect 10232 15444 10284 15453
rect 10324 15487 10376 15496
rect 10324 15453 10334 15487
rect 10334 15453 10368 15487
rect 10368 15453 10376 15487
rect 10324 15444 10376 15453
rect 10600 15487 10652 15496
rect 10600 15453 10609 15487
rect 10609 15453 10643 15487
rect 10643 15453 10652 15487
rect 10600 15444 10652 15453
rect 10876 15444 10928 15496
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 14924 15444 14976 15496
rect 5724 15419 5776 15428
rect 5724 15385 5733 15419
rect 5733 15385 5767 15419
rect 5767 15385 5776 15419
rect 5724 15376 5776 15385
rect 6828 15376 6880 15428
rect 1400 15308 1452 15360
rect 1768 15308 1820 15360
rect 2688 15308 2740 15360
rect 4804 15351 4856 15360
rect 4804 15317 4813 15351
rect 4813 15317 4847 15351
rect 4847 15317 4856 15351
rect 4804 15308 4856 15317
rect 5632 15308 5684 15360
rect 6736 15308 6788 15360
rect 7932 15308 7984 15360
rect 8852 15308 8904 15360
rect 10416 15308 10468 15360
rect 14648 15376 14700 15428
rect 14740 15376 14792 15428
rect 15384 15444 15436 15496
rect 15476 15487 15528 15496
rect 15476 15453 15485 15487
rect 15485 15453 15519 15487
rect 15519 15453 15528 15487
rect 15476 15444 15528 15453
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 16580 15648 16632 15700
rect 17132 15648 17184 15700
rect 18788 15648 18840 15700
rect 20628 15648 20680 15700
rect 16764 15623 16816 15632
rect 16764 15589 16773 15623
rect 16773 15589 16807 15623
rect 16807 15589 16816 15623
rect 16764 15580 16816 15589
rect 18604 15623 18656 15632
rect 18604 15589 18613 15623
rect 18613 15589 18647 15623
rect 18647 15589 18656 15623
rect 18604 15580 18656 15589
rect 18696 15580 18748 15632
rect 22468 15580 22520 15632
rect 19340 15512 19392 15564
rect 21180 15512 21232 15564
rect 21732 15555 21784 15564
rect 21732 15521 21741 15555
rect 21741 15521 21775 15555
rect 21775 15521 21784 15555
rect 21732 15512 21784 15521
rect 23388 15512 23440 15564
rect 16580 15487 16632 15496
rect 16580 15453 16625 15487
rect 16625 15453 16632 15487
rect 16580 15444 16632 15453
rect 10876 15351 10928 15360
rect 10876 15317 10885 15351
rect 10885 15317 10919 15351
rect 10919 15317 10928 15351
rect 10876 15308 10928 15317
rect 14832 15351 14884 15360
rect 14832 15317 14841 15351
rect 14841 15317 14875 15351
rect 14875 15317 14884 15351
rect 14832 15308 14884 15317
rect 15108 15308 15160 15360
rect 16028 15308 16080 15360
rect 17316 15487 17368 15496
rect 17316 15453 17325 15487
rect 17325 15453 17359 15487
rect 17359 15453 17368 15487
rect 17316 15444 17368 15453
rect 18144 15444 18196 15496
rect 19892 15487 19944 15496
rect 19892 15453 19901 15487
rect 19901 15453 19935 15487
rect 19935 15453 19944 15487
rect 19892 15444 19944 15453
rect 16948 15376 17000 15428
rect 18972 15376 19024 15428
rect 19248 15376 19300 15428
rect 19524 15308 19576 15360
rect 19984 15308 20036 15360
rect 20904 15444 20956 15496
rect 21456 15487 21508 15496
rect 21456 15453 21465 15487
rect 21465 15453 21499 15487
rect 21499 15453 21508 15487
rect 21456 15444 21508 15453
rect 20628 15376 20680 15428
rect 21640 15444 21692 15496
rect 22100 15444 22152 15496
rect 23204 15444 23256 15496
rect 23480 15487 23532 15496
rect 23480 15453 23489 15487
rect 23489 15453 23523 15487
rect 23523 15453 23532 15487
rect 23480 15444 23532 15453
rect 23572 15444 23624 15496
rect 20812 15308 20864 15360
rect 22008 15308 22060 15360
rect 23940 15351 23992 15360
rect 23940 15317 23949 15351
rect 23949 15317 23983 15351
rect 23983 15317 23992 15351
rect 23940 15308 23992 15317
rect 8214 15206 8266 15258
rect 8278 15206 8330 15258
rect 8342 15206 8394 15258
rect 8406 15206 8458 15258
rect 8470 15206 8522 15258
rect 16214 15206 16266 15258
rect 16278 15206 16330 15258
rect 16342 15206 16394 15258
rect 16406 15206 16458 15258
rect 16470 15206 16522 15258
rect 24214 15206 24266 15258
rect 24278 15206 24330 15258
rect 24342 15206 24394 15258
rect 24406 15206 24458 15258
rect 24470 15206 24522 15258
rect 2044 15104 2096 15156
rect 2320 15147 2372 15156
rect 2320 15113 2345 15147
rect 2345 15113 2372 15147
rect 2320 15104 2372 15113
rect 2136 15079 2188 15088
rect 2136 15045 2145 15079
rect 2145 15045 2179 15079
rect 2179 15045 2188 15079
rect 2136 15036 2188 15045
rect 4068 15104 4120 15156
rect 4804 15104 4856 15156
rect 5172 15104 5224 15156
rect 3976 15036 4028 15088
rect 1400 14968 1452 15020
rect 2964 15011 3016 15020
rect 2964 14977 2973 15011
rect 2973 14977 3007 15011
rect 3007 14977 3016 15011
rect 2964 14968 3016 14977
rect 6000 15036 6052 15088
rect 7656 15036 7708 15088
rect 7012 14968 7064 15020
rect 7104 15011 7156 15020
rect 7104 14977 7113 15011
rect 7113 14977 7147 15011
rect 7147 14977 7156 15011
rect 7104 14968 7156 14977
rect 8852 15147 8904 15156
rect 8852 15113 8861 15147
rect 8861 15113 8895 15147
rect 8895 15113 8904 15147
rect 8852 15104 8904 15113
rect 10232 15104 10284 15156
rect 10600 15036 10652 15088
rect 11704 15036 11756 15088
rect 13084 15104 13136 15156
rect 9864 15011 9916 15020
rect 9864 14977 9873 15011
rect 9873 14977 9907 15011
rect 9907 14977 9916 15011
rect 9864 14968 9916 14977
rect 3884 14900 3936 14952
rect 7840 14900 7892 14952
rect 10140 15011 10192 15020
rect 10140 14977 10149 15011
rect 10149 14977 10183 15011
rect 10183 14977 10192 15011
rect 10140 14968 10192 14977
rect 10416 14900 10468 14952
rect 11336 14968 11388 15020
rect 11612 15011 11664 15020
rect 11612 14977 11621 15011
rect 11621 14977 11655 15011
rect 11655 14977 11664 15011
rect 11612 14968 11664 14977
rect 11796 15011 11848 15020
rect 11796 14977 11805 15011
rect 11805 14977 11839 15011
rect 11839 14977 11848 15011
rect 11796 14968 11848 14977
rect 11980 14968 12032 15020
rect 13728 15036 13780 15088
rect 12716 15011 12768 15020
rect 12716 14977 12733 15011
rect 12733 14977 12768 15011
rect 12716 14968 12768 14977
rect 12808 15011 12860 15020
rect 12808 14977 12817 15011
rect 12817 14977 12851 15011
rect 12851 14977 12860 15011
rect 12808 14968 12860 14977
rect 13268 14968 13320 15020
rect 13360 14968 13412 15020
rect 13820 14968 13872 15020
rect 14740 15036 14792 15088
rect 15016 15104 15068 15156
rect 15660 15104 15712 15156
rect 16028 15104 16080 15156
rect 16948 15104 17000 15156
rect 17316 15147 17368 15156
rect 17316 15113 17325 15147
rect 17325 15113 17359 15147
rect 17359 15113 17368 15147
rect 17316 15104 17368 15113
rect 15568 15036 15620 15088
rect 18788 15104 18840 15156
rect 19248 15104 19300 15156
rect 19432 15147 19484 15156
rect 19432 15113 19441 15147
rect 19441 15113 19475 15147
rect 19475 15113 19484 15147
rect 19432 15104 19484 15113
rect 19708 15104 19760 15156
rect 15292 14968 15344 15020
rect 14648 14900 14700 14952
rect 14924 14900 14976 14952
rect 15476 14900 15528 14952
rect 15844 14900 15896 14952
rect 16120 15011 16172 15020
rect 16120 14977 16129 15011
rect 16129 14977 16163 15011
rect 16163 14977 16172 15011
rect 16120 14968 16172 14977
rect 18144 15036 18196 15088
rect 18420 15079 18472 15088
rect 18420 15045 18429 15079
rect 18429 15045 18463 15079
rect 18463 15045 18472 15079
rect 18420 15036 18472 15045
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 17224 14968 17276 15020
rect 17316 14900 17368 14952
rect 1952 14764 2004 14816
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 5816 14807 5868 14816
rect 5816 14773 5825 14807
rect 5825 14773 5859 14807
rect 5859 14773 5868 14807
rect 5816 14764 5868 14773
rect 6000 14807 6052 14816
rect 6000 14773 6009 14807
rect 6009 14773 6043 14807
rect 6043 14773 6052 14807
rect 6000 14764 6052 14773
rect 10600 14832 10652 14884
rect 11152 14832 11204 14884
rect 10508 14764 10560 14816
rect 10784 14807 10836 14816
rect 10784 14773 10793 14807
rect 10793 14773 10827 14807
rect 10827 14773 10836 14807
rect 10784 14764 10836 14773
rect 10968 14807 11020 14816
rect 10968 14773 10977 14807
rect 10977 14773 11011 14807
rect 11011 14773 11020 14807
rect 10968 14764 11020 14773
rect 17776 14832 17828 14884
rect 15016 14764 15068 14816
rect 15200 14764 15252 14816
rect 17040 14764 17092 14816
rect 17592 14764 17644 14816
rect 19340 14968 19392 15020
rect 19616 15011 19668 15020
rect 19616 14977 19625 15011
rect 19625 14977 19659 15011
rect 19659 14977 19668 15011
rect 19616 14968 19668 14977
rect 19892 14968 19944 15020
rect 20628 15104 20680 15156
rect 20904 15036 20956 15088
rect 20628 14968 20680 15020
rect 20996 15011 21048 15020
rect 20996 14977 21005 15011
rect 21005 14977 21039 15011
rect 21039 14977 21048 15011
rect 20996 14968 21048 14977
rect 21180 15011 21232 15020
rect 21180 14977 21189 15011
rect 21189 14977 21223 15011
rect 21223 14977 21232 15011
rect 21180 14968 21232 14977
rect 21272 15011 21324 15020
rect 21272 14977 21281 15011
rect 21281 14977 21315 15011
rect 21315 14977 21324 15011
rect 21272 14968 21324 14977
rect 22100 15104 22152 15156
rect 22192 15104 22244 15156
rect 21732 15036 21784 15088
rect 21548 14968 21600 15020
rect 23388 15079 23440 15088
rect 23388 15045 23397 15079
rect 23397 15045 23431 15079
rect 23431 15045 23440 15079
rect 23388 15036 23440 15045
rect 23572 15036 23624 15088
rect 22100 14968 22152 15020
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 22376 15011 22428 15020
rect 22376 14977 22390 15011
rect 22390 14977 22424 15011
rect 22424 14977 22428 15011
rect 22376 14968 22428 14977
rect 23756 14968 23808 15020
rect 24124 14968 24176 15020
rect 22468 14900 22520 14952
rect 18052 14832 18104 14884
rect 22284 14832 22336 14884
rect 25044 14832 25096 14884
rect 23020 14764 23072 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 12214 14662 12266 14714
rect 12278 14662 12330 14714
rect 12342 14662 12394 14714
rect 12406 14662 12458 14714
rect 12470 14662 12522 14714
rect 20214 14662 20266 14714
rect 20278 14662 20330 14714
rect 20342 14662 20394 14714
rect 20406 14662 20458 14714
rect 20470 14662 20522 14714
rect 3884 14603 3936 14612
rect 3884 14569 3893 14603
rect 3893 14569 3927 14603
rect 3927 14569 3936 14603
rect 3884 14560 3936 14569
rect 4068 14492 4120 14544
rect 7656 14560 7708 14612
rect 7840 14603 7892 14612
rect 7840 14569 7849 14603
rect 7849 14569 7883 14603
rect 7883 14569 7892 14603
rect 7840 14560 7892 14569
rect 8668 14560 8720 14612
rect 9312 14603 9364 14612
rect 9312 14569 9321 14603
rect 9321 14569 9355 14603
rect 9355 14569 9364 14603
rect 9312 14560 9364 14569
rect 9956 14560 10008 14612
rect 11796 14560 11848 14612
rect 12808 14560 12860 14612
rect 13268 14560 13320 14612
rect 15476 14560 15528 14612
rect 16948 14603 17000 14612
rect 16948 14569 16957 14603
rect 16957 14569 16991 14603
rect 16991 14569 17000 14603
rect 16948 14560 17000 14569
rect 17316 14603 17368 14612
rect 17316 14569 17325 14603
rect 17325 14569 17359 14603
rect 17359 14569 17368 14603
rect 17316 14560 17368 14569
rect 19340 14560 19392 14612
rect 19616 14560 19668 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 21364 14560 21416 14612
rect 1492 14467 1544 14476
rect 1492 14433 1501 14467
rect 1501 14433 1535 14467
rect 1535 14433 1544 14467
rect 1492 14424 1544 14433
rect 2964 14424 3016 14476
rect 4896 14424 4948 14476
rect 10968 14492 11020 14544
rect 11888 14492 11940 14544
rect 12072 14492 12124 14544
rect 12900 14492 12952 14544
rect 13544 14492 13596 14544
rect 7104 14424 7156 14476
rect 7932 14424 7984 14476
rect 4804 14356 4856 14408
rect 9128 14424 9180 14476
rect 8576 14356 8628 14408
rect 9772 14356 9824 14408
rect 10416 14399 10468 14408
rect 10416 14365 10425 14399
rect 10425 14365 10459 14399
rect 10459 14365 10468 14399
rect 10416 14356 10468 14365
rect 10784 14356 10836 14408
rect 1768 14331 1820 14340
rect 1768 14297 1777 14331
rect 1777 14297 1811 14331
rect 1811 14297 1820 14331
rect 1768 14288 1820 14297
rect 2504 14288 2556 14340
rect 5540 14288 5592 14340
rect 6000 14288 6052 14340
rect 7012 14288 7064 14340
rect 8024 14288 8076 14340
rect 8116 14288 8168 14340
rect 9220 14288 9272 14340
rect 2688 14220 2740 14272
rect 3332 14220 3384 14272
rect 6736 14263 6788 14272
rect 6736 14229 6745 14263
rect 6745 14229 6779 14263
rect 6779 14229 6788 14263
rect 6736 14220 6788 14229
rect 6920 14220 6972 14272
rect 8760 14220 8812 14272
rect 9036 14220 9088 14272
rect 9864 14288 9916 14340
rect 11244 14399 11296 14408
rect 11244 14365 11253 14399
rect 11253 14365 11287 14399
rect 11287 14365 11296 14399
rect 11244 14356 11296 14365
rect 11428 14399 11480 14408
rect 11428 14365 11437 14399
rect 11437 14365 11471 14399
rect 11471 14365 11480 14399
rect 11428 14356 11480 14365
rect 11796 14356 11848 14408
rect 11336 14288 11388 14340
rect 12072 14399 12124 14408
rect 12072 14365 12081 14399
rect 12081 14365 12115 14399
rect 12115 14365 12124 14399
rect 12072 14356 12124 14365
rect 12900 14356 12952 14408
rect 13268 14399 13320 14408
rect 13268 14365 13277 14399
rect 13277 14365 13311 14399
rect 13311 14365 13320 14399
rect 13268 14356 13320 14365
rect 15384 14467 15436 14476
rect 15384 14433 15393 14467
rect 15393 14433 15427 14467
rect 15427 14433 15436 14467
rect 15384 14424 15436 14433
rect 14096 14288 14148 14340
rect 15016 14356 15068 14408
rect 15108 14399 15160 14408
rect 15108 14365 15117 14399
rect 15117 14365 15151 14399
rect 15151 14365 15160 14399
rect 15108 14356 15160 14365
rect 14648 14288 14700 14340
rect 9680 14220 9732 14272
rect 11244 14220 11296 14272
rect 11980 14220 12032 14272
rect 12992 14220 13044 14272
rect 13360 14220 13412 14272
rect 13452 14263 13504 14272
rect 13452 14229 13461 14263
rect 13461 14229 13495 14263
rect 13495 14229 13504 14263
rect 13452 14220 13504 14229
rect 13912 14220 13964 14272
rect 15476 14288 15528 14340
rect 16948 14399 17000 14408
rect 16948 14365 16957 14399
rect 16957 14365 16991 14399
rect 16991 14365 17000 14399
rect 16948 14356 17000 14365
rect 17132 14399 17184 14408
rect 17132 14365 17141 14399
rect 17141 14365 17175 14399
rect 17175 14365 17184 14399
rect 17132 14356 17184 14365
rect 15752 14220 15804 14272
rect 17684 14288 17736 14340
rect 19432 14424 19484 14476
rect 18512 14331 18564 14340
rect 18512 14297 18521 14331
rect 18521 14297 18555 14331
rect 18555 14297 18564 14331
rect 18512 14288 18564 14297
rect 19340 14288 19392 14340
rect 20628 14356 20680 14408
rect 21088 14356 21140 14408
rect 23112 14492 23164 14544
rect 23756 14535 23808 14544
rect 23756 14501 23765 14535
rect 23765 14501 23799 14535
rect 23799 14501 23808 14535
rect 23756 14492 23808 14501
rect 22284 14399 22336 14408
rect 22284 14365 22293 14399
rect 22293 14365 22327 14399
rect 22327 14365 22336 14399
rect 22284 14356 22336 14365
rect 22560 14356 22612 14408
rect 16764 14220 16816 14272
rect 23664 14288 23716 14340
rect 20076 14220 20128 14272
rect 23756 14220 23808 14272
rect 8214 14118 8266 14170
rect 8278 14118 8330 14170
rect 8342 14118 8394 14170
rect 8406 14118 8458 14170
rect 8470 14118 8522 14170
rect 16214 14118 16266 14170
rect 16278 14118 16330 14170
rect 16342 14118 16394 14170
rect 16406 14118 16458 14170
rect 16470 14118 16522 14170
rect 24214 14118 24266 14170
rect 24278 14118 24330 14170
rect 24342 14118 24394 14170
rect 24406 14118 24458 14170
rect 24470 14118 24522 14170
rect 2136 14016 2188 14068
rect 2872 13948 2924 14000
rect 3332 14059 3384 14068
rect 3332 14025 3341 14059
rect 3341 14025 3375 14059
rect 3375 14025 3384 14059
rect 3332 14016 3384 14025
rect 3976 14059 4028 14068
rect 3976 14025 3985 14059
rect 3985 14025 4019 14059
rect 4019 14025 4028 14059
rect 3976 14016 4028 14025
rect 5908 14016 5960 14068
rect 6920 14016 6972 14068
rect 8116 14016 8168 14068
rect 9220 14016 9272 14068
rect 10968 14016 11020 14068
rect 12072 14016 12124 14068
rect 13360 14059 13412 14068
rect 13360 14025 13377 14059
rect 13377 14025 13412 14059
rect 13360 14016 13412 14025
rect 14096 14016 14148 14068
rect 15660 14059 15712 14068
rect 15660 14025 15669 14059
rect 15669 14025 15703 14059
rect 15703 14025 15712 14059
rect 15660 14016 15712 14025
rect 16672 14016 16724 14068
rect 16764 14059 16816 14068
rect 16764 14025 16773 14059
rect 16773 14025 16807 14059
rect 16807 14025 16816 14059
rect 16764 14016 16816 14025
rect 17040 14016 17092 14068
rect 20812 14016 20864 14068
rect 21088 14059 21140 14068
rect 21088 14025 21097 14059
rect 21097 14025 21131 14059
rect 21131 14025 21140 14059
rect 21088 14016 21140 14025
rect 21916 14016 21968 14068
rect 1492 13880 1544 13932
rect 6828 13991 6880 14000
rect 6828 13957 6837 13991
rect 6837 13957 6871 13991
rect 6871 13957 6880 13991
rect 6828 13948 6880 13957
rect 9036 13948 9088 14000
rect 4068 13880 4120 13932
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 8944 13880 8996 13932
rect 11060 13948 11112 14000
rect 10324 13880 10376 13932
rect 10508 13923 10560 13932
rect 10508 13889 10517 13923
rect 10517 13889 10551 13923
rect 10551 13889 10560 13923
rect 10508 13880 10560 13889
rect 10784 13923 10836 13932
rect 10784 13889 10793 13923
rect 10793 13889 10827 13923
rect 10827 13889 10836 13923
rect 10784 13880 10836 13889
rect 1860 13855 1912 13864
rect 1860 13821 1869 13855
rect 1869 13821 1903 13855
rect 1903 13821 1912 13855
rect 1860 13812 1912 13821
rect 7380 13855 7432 13864
rect 7380 13821 7389 13855
rect 7389 13821 7423 13855
rect 7423 13821 7432 13855
rect 7380 13812 7432 13821
rect 9680 13812 9732 13864
rect 10600 13812 10652 13864
rect 10968 13855 11020 13864
rect 10968 13821 10977 13855
rect 10977 13821 11011 13855
rect 11011 13821 11020 13855
rect 10968 13812 11020 13821
rect 11612 13880 11664 13932
rect 11888 13923 11940 13932
rect 11888 13889 11897 13923
rect 11897 13889 11931 13923
rect 11931 13889 11940 13923
rect 11888 13880 11940 13889
rect 12072 13880 12124 13932
rect 12808 13880 12860 13932
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 14096 13923 14148 13932
rect 14096 13889 14105 13923
rect 14105 13889 14139 13923
rect 14139 13889 14148 13923
rect 14096 13880 14148 13889
rect 1952 13676 2004 13728
rect 11152 13744 11204 13796
rect 11336 13744 11388 13796
rect 12624 13812 12676 13864
rect 12992 13812 13044 13864
rect 14004 13812 14056 13864
rect 15016 13923 15068 13932
rect 15016 13889 15025 13923
rect 15025 13889 15059 13923
rect 15059 13889 15068 13923
rect 15016 13880 15068 13889
rect 15200 13923 15252 13932
rect 15200 13889 15209 13923
rect 15209 13889 15243 13923
rect 15243 13889 15252 13923
rect 15200 13880 15252 13889
rect 16120 13880 16172 13932
rect 16948 13923 17000 13932
rect 16948 13889 16957 13923
rect 16957 13889 16991 13923
rect 16991 13889 17000 13923
rect 16948 13880 17000 13889
rect 17132 13923 17184 13932
rect 17132 13889 17141 13923
rect 17141 13889 17175 13923
rect 17175 13889 17184 13923
rect 17132 13880 17184 13889
rect 14924 13812 14976 13864
rect 16672 13812 16724 13864
rect 17592 13923 17644 13932
rect 17592 13889 17601 13923
rect 17601 13889 17635 13923
rect 17635 13889 17644 13923
rect 17592 13880 17644 13889
rect 19432 13991 19484 14000
rect 19432 13957 19441 13991
rect 19441 13957 19475 13991
rect 19475 13957 19484 13991
rect 19432 13948 19484 13957
rect 22560 13991 22612 14000
rect 22560 13957 22569 13991
rect 22569 13957 22603 13991
rect 22603 13957 22612 13991
rect 22560 13948 22612 13957
rect 18328 13880 18380 13932
rect 19340 13923 19392 13932
rect 19340 13889 19349 13923
rect 19349 13889 19383 13923
rect 19383 13889 19392 13923
rect 19340 13880 19392 13889
rect 17316 13812 17368 13864
rect 19984 13880 20036 13932
rect 22100 13880 22152 13932
rect 22192 13923 22244 13932
rect 22192 13889 22201 13923
rect 22201 13889 22235 13923
rect 22235 13889 22244 13923
rect 22192 13880 22244 13889
rect 23756 13991 23808 14000
rect 23756 13957 23765 13991
rect 23765 13957 23799 13991
rect 23799 13957 23808 13991
rect 23756 13948 23808 13957
rect 23940 13948 23992 14000
rect 11980 13744 12032 13796
rect 17132 13744 17184 13796
rect 24032 13812 24084 13864
rect 21548 13744 21600 13796
rect 3976 13676 4028 13728
rect 6184 13676 6236 13728
rect 8760 13676 8812 13728
rect 9312 13719 9364 13728
rect 9312 13685 9321 13719
rect 9321 13685 9355 13719
rect 9355 13685 9364 13719
rect 9312 13676 9364 13685
rect 9496 13719 9548 13728
rect 9496 13685 9505 13719
rect 9505 13685 9539 13719
rect 9539 13685 9548 13719
rect 9496 13676 9548 13685
rect 10140 13719 10192 13728
rect 10140 13685 10149 13719
rect 10149 13685 10183 13719
rect 10183 13685 10192 13719
rect 10140 13676 10192 13685
rect 11796 13719 11848 13728
rect 11796 13685 11805 13719
rect 11805 13685 11839 13719
rect 11839 13685 11848 13719
rect 11796 13676 11848 13685
rect 11888 13676 11940 13728
rect 13820 13676 13872 13728
rect 14832 13676 14884 13728
rect 15016 13676 15068 13728
rect 20628 13676 20680 13728
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 12214 13574 12266 13626
rect 12278 13574 12330 13626
rect 12342 13574 12394 13626
rect 12406 13574 12458 13626
rect 12470 13574 12522 13626
rect 20214 13574 20266 13626
rect 20278 13574 20330 13626
rect 20342 13574 20394 13626
rect 20406 13574 20458 13626
rect 20470 13574 20522 13626
rect 1952 13472 2004 13524
rect 2872 13472 2924 13524
rect 6184 13515 6236 13524
rect 6184 13481 6193 13515
rect 6193 13481 6227 13515
rect 6227 13481 6236 13515
rect 6184 13472 6236 13481
rect 7380 13472 7432 13524
rect 9312 13515 9364 13524
rect 9312 13481 9321 13515
rect 9321 13481 9355 13515
rect 9355 13481 9364 13515
rect 9312 13472 9364 13481
rect 11980 13472 12032 13524
rect 14464 13472 14516 13524
rect 15200 13472 15252 13524
rect 16120 13472 16172 13524
rect 16948 13515 17000 13524
rect 16948 13481 16957 13515
rect 16957 13481 16991 13515
rect 16991 13481 17000 13515
rect 16948 13472 17000 13481
rect 1860 13404 1912 13456
rect 10876 13404 10928 13456
rect 22468 13472 22520 13524
rect 19432 13404 19484 13456
rect 22192 13404 22244 13456
rect 1952 13336 2004 13388
rect 2228 13336 2280 13388
rect 3424 13336 3476 13388
rect 4896 13336 4948 13388
rect 6736 13336 6788 13388
rect 8116 13336 8168 13388
rect 2136 13268 2188 13320
rect 3332 13268 3384 13320
rect 8576 13336 8628 13388
rect 10784 13336 10836 13388
rect 13176 13336 13228 13388
rect 9864 13268 9916 13320
rect 1860 13243 1912 13252
rect 1860 13209 1869 13243
rect 1869 13209 1903 13243
rect 1903 13209 1912 13243
rect 1860 13200 1912 13209
rect 3976 13200 4028 13252
rect 8116 13200 8168 13252
rect 8944 13200 8996 13252
rect 9312 13243 9364 13252
rect 1308 13132 1360 13184
rect 2044 13175 2096 13184
rect 2044 13141 2069 13175
rect 2069 13141 2096 13175
rect 2044 13132 2096 13141
rect 3608 13132 3660 13184
rect 9128 13175 9180 13184
rect 9128 13141 9137 13175
rect 9137 13141 9171 13175
rect 9171 13141 9180 13175
rect 9128 13132 9180 13141
rect 9312 13209 9339 13243
rect 9339 13209 9364 13243
rect 9312 13200 9364 13209
rect 10324 13268 10376 13320
rect 11152 13268 11204 13320
rect 10692 13200 10744 13252
rect 11704 13243 11756 13252
rect 11704 13209 11731 13243
rect 11731 13209 11756 13243
rect 11704 13200 11756 13209
rect 12624 13311 12676 13320
rect 12624 13277 12633 13311
rect 12633 13277 12667 13311
rect 12667 13277 12676 13311
rect 12624 13268 12676 13277
rect 12900 13268 12952 13320
rect 15292 13336 15344 13388
rect 15752 13336 15804 13388
rect 13636 13311 13688 13320
rect 13636 13277 13645 13311
rect 13645 13277 13679 13311
rect 13679 13277 13688 13311
rect 13636 13268 13688 13277
rect 13912 13268 13964 13320
rect 15016 13268 15068 13320
rect 15936 13268 15988 13320
rect 16672 13379 16724 13388
rect 16672 13345 16681 13379
rect 16681 13345 16715 13379
rect 16715 13345 16724 13379
rect 16672 13336 16724 13345
rect 17500 13336 17552 13388
rect 18328 13379 18380 13388
rect 18328 13345 18337 13379
rect 18337 13345 18371 13379
rect 18371 13345 18380 13379
rect 18328 13336 18380 13345
rect 18420 13336 18472 13388
rect 19708 13336 19760 13388
rect 20076 13379 20128 13388
rect 20076 13345 20085 13379
rect 20085 13345 20119 13379
rect 20119 13345 20128 13379
rect 20076 13336 20128 13345
rect 21456 13336 21508 13388
rect 12992 13200 13044 13252
rect 13452 13200 13504 13252
rect 17960 13311 18012 13320
rect 17960 13277 17969 13311
rect 17969 13277 18003 13311
rect 18003 13277 18012 13311
rect 17960 13268 18012 13277
rect 19340 13268 19392 13320
rect 10968 13132 11020 13184
rect 11520 13175 11572 13184
rect 11520 13141 11529 13175
rect 11529 13141 11563 13175
rect 11563 13141 11572 13175
rect 11520 13132 11572 13141
rect 12072 13132 12124 13184
rect 14648 13132 14700 13184
rect 16764 13200 16816 13252
rect 18512 13200 18564 13252
rect 18880 13243 18932 13252
rect 18880 13209 18889 13243
rect 18889 13209 18923 13243
rect 18923 13209 18932 13243
rect 18880 13200 18932 13209
rect 19984 13243 20036 13252
rect 19984 13209 19993 13243
rect 19993 13209 20027 13243
rect 20027 13209 20036 13243
rect 19984 13200 20036 13209
rect 22836 13311 22888 13320
rect 22836 13277 22845 13311
rect 22845 13277 22879 13311
rect 22879 13277 22888 13311
rect 22836 13268 22888 13277
rect 23480 13268 23532 13320
rect 20720 13200 20772 13252
rect 23020 13200 23072 13252
rect 23664 13243 23716 13252
rect 23664 13209 23673 13243
rect 23673 13209 23707 13243
rect 23707 13209 23716 13243
rect 23664 13200 23716 13209
rect 21272 13132 21324 13184
rect 22192 13132 22244 13184
rect 24124 13175 24176 13184
rect 24124 13141 24133 13175
rect 24133 13141 24167 13175
rect 24167 13141 24176 13175
rect 24124 13132 24176 13141
rect 8214 13030 8266 13082
rect 8278 13030 8330 13082
rect 8342 13030 8394 13082
rect 8406 13030 8458 13082
rect 8470 13030 8522 13082
rect 16214 13030 16266 13082
rect 16278 13030 16330 13082
rect 16342 13030 16394 13082
rect 16406 13030 16458 13082
rect 16470 13030 16522 13082
rect 24214 13030 24266 13082
rect 24278 13030 24330 13082
rect 24342 13030 24394 13082
rect 24406 13030 24458 13082
rect 24470 13030 24522 13082
rect 9772 12928 9824 12980
rect 10600 12928 10652 12980
rect 11704 12928 11756 12980
rect 1860 12860 1912 12912
rect 2136 12860 2188 12912
rect 1308 12792 1360 12844
rect 3240 12860 3292 12912
rect 4068 12903 4120 12912
rect 4068 12869 4077 12903
rect 4077 12869 4111 12903
rect 4111 12869 4120 12903
rect 4068 12860 4120 12869
rect 5724 12903 5776 12912
rect 5724 12869 5733 12903
rect 5733 12869 5767 12903
rect 5767 12869 5776 12903
rect 5724 12860 5776 12869
rect 5908 12903 5960 12912
rect 5908 12869 5933 12903
rect 5933 12869 5960 12903
rect 5908 12860 5960 12869
rect 6552 12860 6604 12912
rect 4620 12792 4672 12844
rect 8576 12860 8628 12912
rect 9496 12860 9548 12912
rect 10324 12860 10376 12912
rect 11612 12835 11664 12844
rect 11612 12801 11621 12835
rect 11621 12801 11655 12835
rect 11655 12801 11664 12835
rect 11612 12792 11664 12801
rect 11704 12835 11756 12844
rect 11704 12801 11713 12835
rect 11713 12801 11747 12835
rect 11747 12801 11756 12835
rect 11704 12792 11756 12801
rect 2228 12724 2280 12776
rect 2780 12656 2832 12708
rect 3148 12767 3200 12776
rect 3148 12733 3157 12767
rect 3157 12733 3191 12767
rect 3191 12733 3200 12767
rect 3148 12724 3200 12733
rect 3424 12724 3476 12776
rect 7104 12724 7156 12776
rect 9496 12724 9548 12776
rect 2228 12631 2280 12640
rect 2228 12597 2237 12631
rect 2237 12597 2271 12631
rect 2271 12597 2280 12631
rect 2228 12588 2280 12597
rect 2320 12588 2372 12640
rect 3700 12631 3752 12640
rect 3700 12597 3709 12631
rect 3709 12597 3743 12631
rect 3743 12597 3752 12631
rect 3700 12588 3752 12597
rect 4712 12588 4764 12640
rect 5816 12588 5868 12640
rect 6736 12656 6788 12708
rect 6184 12588 6236 12640
rect 8668 12588 8720 12640
rect 8944 12588 8996 12640
rect 11336 12724 11388 12776
rect 11888 12928 11940 12980
rect 12072 12928 12124 12980
rect 11980 12860 12032 12912
rect 13912 12928 13964 12980
rect 11888 12835 11940 12844
rect 11888 12801 11897 12835
rect 11897 12801 11931 12835
rect 11931 12801 11940 12835
rect 11888 12792 11940 12801
rect 12072 12835 12124 12844
rect 12072 12801 12081 12835
rect 12081 12801 12115 12835
rect 12115 12801 12124 12835
rect 12072 12792 12124 12801
rect 12992 12835 13044 12844
rect 12992 12801 13002 12835
rect 13002 12801 13036 12835
rect 13036 12801 13044 12835
rect 12992 12792 13044 12801
rect 13268 12792 13320 12844
rect 12624 12724 12676 12776
rect 11796 12656 11848 12708
rect 14096 12767 14148 12776
rect 14096 12733 14105 12767
rect 14105 12733 14139 12767
rect 14139 12733 14148 12767
rect 14096 12724 14148 12733
rect 14648 12835 14700 12844
rect 14648 12801 14657 12835
rect 14657 12801 14691 12835
rect 14691 12801 14700 12835
rect 14648 12792 14700 12801
rect 14832 12792 14884 12844
rect 14924 12835 14976 12844
rect 14924 12801 14933 12835
rect 14933 12801 14967 12835
rect 14967 12801 14976 12835
rect 14924 12792 14976 12801
rect 15936 12928 15988 12980
rect 16764 12928 16816 12980
rect 20996 12928 21048 12980
rect 21548 12928 21600 12980
rect 16672 12860 16724 12912
rect 16120 12792 16172 12844
rect 16948 12860 17000 12912
rect 18052 12860 18104 12912
rect 21456 12860 21508 12912
rect 15660 12724 15712 12776
rect 15844 12724 15896 12776
rect 15752 12656 15804 12708
rect 14924 12588 14976 12640
rect 15108 12631 15160 12640
rect 15108 12597 15117 12631
rect 15117 12597 15151 12631
rect 15151 12597 15160 12631
rect 15108 12588 15160 12597
rect 15936 12588 15988 12640
rect 17776 12724 17828 12776
rect 20628 12792 20680 12844
rect 21088 12792 21140 12844
rect 21640 12792 21692 12844
rect 22100 12792 22152 12844
rect 21272 12767 21324 12776
rect 21272 12733 21281 12767
rect 21281 12733 21315 12767
rect 21315 12733 21324 12767
rect 21272 12724 21324 12733
rect 21364 12656 21416 12708
rect 22836 12835 22888 12844
rect 22836 12801 22845 12835
rect 22845 12801 22879 12835
rect 22879 12801 22888 12835
rect 22836 12792 22888 12801
rect 23112 12767 23164 12776
rect 23112 12733 23121 12767
rect 23121 12733 23155 12767
rect 23155 12733 23164 12767
rect 23112 12724 23164 12733
rect 19800 12588 19852 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 12214 12486 12266 12538
rect 12278 12486 12330 12538
rect 12342 12486 12394 12538
rect 12406 12486 12458 12538
rect 12470 12486 12522 12538
rect 20214 12486 20266 12538
rect 20278 12486 20330 12538
rect 20342 12486 20394 12538
rect 20406 12486 20458 12538
rect 20470 12486 20522 12538
rect 2320 12248 2372 12300
rect 4896 12384 4948 12436
rect 1492 12223 1544 12232
rect 1492 12189 1501 12223
rect 1501 12189 1535 12223
rect 1535 12189 1544 12223
rect 1492 12180 1544 12189
rect 3148 12180 3200 12232
rect 4068 12180 4120 12232
rect 2780 12112 2832 12164
rect 3424 12112 3476 12164
rect 7104 12248 7156 12300
rect 9496 12384 9548 12436
rect 11980 12384 12032 12436
rect 7472 12291 7524 12300
rect 7472 12257 7481 12291
rect 7481 12257 7515 12291
rect 7515 12257 7524 12291
rect 7472 12248 7524 12257
rect 10968 12248 11020 12300
rect 11428 12248 11480 12300
rect 8668 12180 8720 12232
rect 9772 12180 9824 12232
rect 9956 12180 10008 12232
rect 11060 12180 11112 12232
rect 11244 12180 11296 12232
rect 11888 12180 11940 12232
rect 12072 12180 12124 12232
rect 12900 12248 12952 12300
rect 14004 12316 14056 12368
rect 12624 12223 12676 12232
rect 12624 12189 12633 12223
rect 12633 12189 12667 12223
rect 12667 12189 12676 12223
rect 12624 12180 12676 12189
rect 12808 12180 12860 12232
rect 14832 12248 14884 12300
rect 13452 12223 13504 12232
rect 13452 12189 13461 12223
rect 13461 12189 13495 12223
rect 13495 12189 13504 12223
rect 13452 12180 13504 12189
rect 13544 12223 13596 12232
rect 13544 12189 13553 12223
rect 13553 12189 13587 12223
rect 13587 12189 13596 12223
rect 13544 12180 13596 12189
rect 14648 12180 14700 12232
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 15016 12223 15068 12232
rect 15016 12189 15025 12223
rect 15025 12189 15059 12223
rect 15059 12189 15068 12223
rect 15016 12180 15068 12189
rect 3240 12087 3292 12096
rect 3240 12053 3249 12087
rect 3249 12053 3283 12087
rect 3283 12053 3292 12087
rect 3240 12044 3292 12053
rect 3884 12087 3936 12096
rect 3884 12053 3893 12087
rect 3893 12053 3927 12087
rect 3927 12053 3936 12087
rect 3884 12044 3936 12053
rect 5172 12155 5224 12164
rect 5172 12121 5181 12155
rect 5181 12121 5215 12155
rect 5215 12121 5224 12155
rect 5172 12112 5224 12121
rect 6184 12112 6236 12164
rect 5540 12044 5592 12096
rect 5816 12044 5868 12096
rect 9496 12155 9548 12164
rect 9496 12121 9505 12155
rect 9505 12121 9539 12155
rect 9539 12121 9548 12155
rect 9496 12112 9548 12121
rect 10140 12112 10192 12164
rect 10416 12155 10468 12164
rect 10416 12121 10425 12155
rect 10425 12121 10459 12155
rect 10459 12121 10468 12155
rect 10416 12112 10468 12121
rect 10600 12155 10652 12164
rect 10600 12121 10609 12155
rect 10609 12121 10643 12155
rect 10643 12121 10652 12155
rect 10600 12112 10652 12121
rect 13268 12112 13320 12164
rect 14832 12112 14884 12164
rect 15752 12384 15804 12436
rect 15844 12427 15896 12436
rect 15844 12393 15853 12427
rect 15853 12393 15887 12427
rect 15887 12393 15896 12427
rect 15844 12384 15896 12393
rect 16120 12384 16172 12436
rect 17592 12384 17644 12436
rect 21456 12427 21508 12436
rect 21456 12393 21465 12427
rect 21465 12393 21499 12427
rect 21499 12393 21508 12427
rect 21456 12384 21508 12393
rect 18052 12316 18104 12368
rect 20076 12316 20128 12368
rect 15936 12291 15988 12300
rect 15936 12257 15945 12291
rect 15945 12257 15979 12291
rect 15979 12257 15988 12291
rect 15936 12248 15988 12257
rect 16120 12248 16172 12300
rect 17132 12248 17184 12300
rect 17684 12248 17736 12300
rect 15292 12180 15344 12232
rect 15752 12223 15804 12232
rect 15752 12189 15761 12223
rect 15761 12189 15795 12223
rect 15795 12189 15804 12223
rect 15752 12180 15804 12189
rect 16028 12180 16080 12232
rect 17224 12180 17276 12232
rect 18328 12223 18380 12232
rect 18328 12189 18337 12223
rect 18337 12189 18371 12223
rect 18371 12189 18380 12223
rect 18328 12180 18380 12189
rect 6920 12087 6972 12096
rect 6920 12053 6929 12087
rect 6929 12053 6963 12087
rect 6963 12053 6972 12087
rect 6920 12044 6972 12053
rect 8576 12044 8628 12096
rect 10232 12044 10284 12096
rect 10324 12087 10376 12096
rect 10324 12053 10333 12087
rect 10333 12053 10367 12087
rect 10367 12053 10376 12087
rect 10324 12044 10376 12053
rect 10968 12044 11020 12096
rect 12072 12044 12124 12096
rect 12808 12087 12860 12096
rect 12808 12053 12817 12087
rect 12817 12053 12851 12087
rect 12851 12053 12860 12087
rect 12808 12044 12860 12053
rect 13728 12087 13780 12096
rect 13728 12053 13737 12087
rect 13737 12053 13771 12087
rect 13771 12053 13780 12087
rect 13728 12044 13780 12053
rect 14096 12044 14148 12096
rect 15016 12044 15068 12096
rect 17500 12112 17552 12164
rect 19800 12248 19852 12300
rect 23664 12316 23716 12368
rect 19340 12223 19392 12232
rect 19340 12189 19349 12223
rect 19349 12189 19383 12223
rect 19383 12189 19392 12223
rect 19340 12180 19392 12189
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 20628 12180 20680 12232
rect 19432 12112 19484 12164
rect 15844 12044 15896 12096
rect 17684 12044 17736 12096
rect 17960 12087 18012 12096
rect 17960 12053 17969 12087
rect 17969 12053 18003 12087
rect 18003 12053 18012 12087
rect 17960 12044 18012 12053
rect 20628 12044 20680 12096
rect 22100 12291 22152 12300
rect 22100 12257 22109 12291
rect 22109 12257 22143 12291
rect 22143 12257 22152 12291
rect 22100 12248 22152 12257
rect 20996 12223 21048 12232
rect 20996 12189 21005 12223
rect 21005 12189 21039 12223
rect 21039 12189 21048 12223
rect 20996 12180 21048 12189
rect 21088 12223 21140 12232
rect 21088 12189 21097 12223
rect 21097 12189 21131 12223
rect 21131 12189 21140 12223
rect 21088 12180 21140 12189
rect 21456 12180 21508 12232
rect 21916 12223 21968 12232
rect 21916 12189 21925 12223
rect 21925 12189 21959 12223
rect 21959 12189 21968 12223
rect 21916 12180 21968 12189
rect 22468 12223 22520 12232
rect 22468 12189 22477 12223
rect 22477 12189 22511 12223
rect 22511 12189 22520 12223
rect 22468 12180 22520 12189
rect 23848 12223 23900 12232
rect 23848 12189 23857 12223
rect 23857 12189 23891 12223
rect 23891 12189 23900 12223
rect 23848 12180 23900 12189
rect 8214 11942 8266 11994
rect 8278 11942 8330 11994
rect 8342 11942 8394 11994
rect 8406 11942 8458 11994
rect 8470 11942 8522 11994
rect 16214 11942 16266 11994
rect 16278 11942 16330 11994
rect 16342 11942 16394 11994
rect 16406 11942 16458 11994
rect 16470 11942 16522 11994
rect 24214 11942 24266 11994
rect 24278 11942 24330 11994
rect 24342 11942 24394 11994
rect 24406 11942 24458 11994
rect 24470 11942 24522 11994
rect 3884 11840 3936 11892
rect 4068 11883 4120 11892
rect 4068 11849 4077 11883
rect 4077 11849 4111 11883
rect 4111 11849 4120 11883
rect 4068 11840 4120 11849
rect 4620 11840 4672 11892
rect 5172 11840 5224 11892
rect 5816 11840 5868 11892
rect 6644 11883 6696 11892
rect 6644 11849 6671 11883
rect 6671 11849 6696 11883
rect 6644 11840 6696 11849
rect 5540 11772 5592 11824
rect 7472 11840 7524 11892
rect 9496 11840 9548 11892
rect 10600 11840 10652 11892
rect 11704 11840 11756 11892
rect 1308 11704 1360 11756
rect 3700 11704 3752 11756
rect 5632 11704 5684 11756
rect 1492 11568 1544 11620
rect 5816 11679 5868 11688
rect 5816 11645 5825 11679
rect 5825 11645 5859 11679
rect 5859 11645 5868 11679
rect 5816 11636 5868 11645
rect 6000 11704 6052 11756
rect 7380 11815 7432 11824
rect 7380 11781 7389 11815
rect 7389 11781 7423 11815
rect 7423 11781 7432 11815
rect 7380 11772 7432 11781
rect 9128 11772 9180 11824
rect 9956 11815 10008 11824
rect 9956 11781 9965 11815
rect 9965 11781 9999 11815
rect 9999 11781 10008 11815
rect 9956 11772 10008 11781
rect 10692 11772 10744 11824
rect 6644 11636 6696 11688
rect 7104 11679 7156 11688
rect 7104 11645 7113 11679
rect 7113 11645 7147 11679
rect 7147 11645 7156 11679
rect 7104 11636 7156 11645
rect 5908 11500 5960 11552
rect 6736 11500 6788 11552
rect 7748 11500 7800 11552
rect 8116 11500 8168 11552
rect 10324 11747 10376 11756
rect 10324 11713 10333 11747
rect 10333 11713 10367 11747
rect 10367 11713 10376 11747
rect 10324 11704 10376 11713
rect 11428 11704 11480 11756
rect 13820 11840 13872 11892
rect 12072 11747 12124 11756
rect 12072 11713 12081 11747
rect 12081 11713 12115 11747
rect 12115 11713 12124 11747
rect 12072 11704 12124 11713
rect 13176 11747 13228 11756
rect 13176 11713 13185 11747
rect 13185 11713 13219 11747
rect 13219 11713 13228 11747
rect 13176 11704 13228 11713
rect 15476 11840 15528 11892
rect 16672 11840 16724 11892
rect 19984 11840 20036 11892
rect 20076 11840 20128 11892
rect 14648 11772 14700 11824
rect 10784 11679 10836 11688
rect 10784 11645 10793 11679
rect 10793 11645 10827 11679
rect 10827 11645 10836 11679
rect 10784 11636 10836 11645
rect 11796 11636 11848 11688
rect 11888 11636 11940 11688
rect 13452 11636 13504 11688
rect 14464 11636 14516 11688
rect 15108 11747 15160 11756
rect 15108 11713 15117 11747
rect 15117 11713 15151 11747
rect 15151 11713 15160 11747
rect 15108 11704 15160 11713
rect 18512 11772 18564 11824
rect 20996 11840 21048 11892
rect 20812 11772 20864 11824
rect 21732 11772 21784 11824
rect 15844 11747 15896 11756
rect 15844 11713 15853 11747
rect 15853 11713 15887 11747
rect 15887 11713 15896 11747
rect 15844 11704 15896 11713
rect 14648 11679 14700 11688
rect 14648 11645 14657 11679
rect 14657 11645 14691 11679
rect 14691 11645 14700 11679
rect 14648 11636 14700 11645
rect 15568 11636 15620 11688
rect 15936 11636 15988 11688
rect 19340 11704 19392 11756
rect 16948 11636 17000 11688
rect 9680 11568 9732 11620
rect 11152 11568 11204 11620
rect 11428 11568 11480 11620
rect 11980 11500 12032 11552
rect 12808 11568 12860 11620
rect 19800 11636 19852 11688
rect 20082 11636 20134 11688
rect 19432 11568 19484 11620
rect 20720 11704 20772 11756
rect 21456 11747 21508 11756
rect 21456 11713 21465 11747
rect 21465 11713 21499 11747
rect 21499 11713 21508 11747
rect 21456 11704 21508 11713
rect 22100 11815 22152 11824
rect 22100 11781 22109 11815
rect 22109 11781 22143 11815
rect 22143 11781 22152 11815
rect 22100 11772 22152 11781
rect 23848 11815 23900 11824
rect 23848 11781 23857 11815
rect 23857 11781 23891 11815
rect 23891 11781 23900 11815
rect 23848 11772 23900 11781
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 22744 11704 22796 11756
rect 23020 11704 23072 11756
rect 23388 11704 23440 11756
rect 21088 11636 21140 11688
rect 21364 11636 21416 11688
rect 22192 11568 22244 11620
rect 15108 11500 15160 11552
rect 15936 11500 15988 11552
rect 16028 11543 16080 11552
rect 16028 11509 16037 11543
rect 16037 11509 16071 11543
rect 16071 11509 16080 11543
rect 16028 11500 16080 11509
rect 21272 11500 21324 11552
rect 21548 11500 21600 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 12214 11398 12266 11450
rect 12278 11398 12330 11450
rect 12342 11398 12394 11450
rect 12406 11398 12458 11450
rect 12470 11398 12522 11450
rect 20214 11398 20266 11450
rect 20278 11398 20330 11450
rect 20342 11398 20394 11450
rect 20406 11398 20458 11450
rect 20470 11398 20522 11450
rect 2136 11296 2188 11348
rect 4712 11296 4764 11348
rect 4896 11339 4948 11348
rect 4896 11305 4905 11339
rect 4905 11305 4939 11339
rect 4939 11305 4948 11339
rect 4896 11296 4948 11305
rect 2964 11228 3016 11280
rect 7380 11339 7432 11348
rect 7380 11305 7389 11339
rect 7389 11305 7423 11339
rect 7423 11305 7432 11339
rect 7380 11296 7432 11305
rect 10784 11296 10836 11348
rect 13268 11296 13320 11348
rect 23112 11296 23164 11348
rect 3148 11203 3200 11212
rect 3148 11169 3157 11203
rect 3157 11169 3191 11203
rect 3191 11169 3200 11203
rect 3148 11160 3200 11169
rect 3424 11160 3476 11212
rect 3240 11092 3292 11144
rect 7840 11228 7892 11280
rect 8760 11228 8812 11280
rect 6920 11160 6972 11212
rect 7472 11160 7524 11212
rect 7932 11203 7984 11212
rect 7932 11169 7941 11203
rect 7941 11169 7975 11203
rect 7975 11169 7984 11203
rect 7932 11160 7984 11169
rect 6644 11135 6696 11144
rect 6644 11101 6653 11135
rect 6653 11101 6687 11135
rect 6687 11101 6696 11135
rect 6644 11092 6696 11101
rect 7748 11135 7800 11144
rect 7748 11101 7757 11135
rect 7757 11101 7791 11135
rect 7791 11101 7800 11135
rect 7748 11092 7800 11101
rect 9956 11160 10008 11212
rect 10416 11160 10468 11212
rect 11704 11228 11756 11280
rect 11612 11160 11664 11212
rect 13176 11160 13228 11212
rect 9680 11092 9732 11144
rect 9864 11135 9916 11144
rect 9864 11101 9873 11135
rect 9873 11101 9907 11135
rect 9907 11101 9916 11135
rect 9864 11092 9916 11101
rect 10140 11092 10192 11144
rect 10784 11135 10836 11144
rect 10784 11101 10793 11135
rect 10793 11101 10827 11135
rect 10827 11101 10836 11135
rect 10784 11092 10836 11101
rect 11428 11135 11480 11144
rect 11428 11101 11437 11135
rect 11437 11101 11471 11135
rect 11471 11101 11480 11135
rect 11428 11092 11480 11101
rect 1860 11067 1912 11076
rect 1860 11033 1869 11067
rect 1869 11033 1903 11067
rect 1903 11033 1912 11067
rect 1860 11024 1912 11033
rect 2044 11067 2096 11076
rect 2044 11033 2069 11067
rect 2069 11033 2096 11067
rect 2044 11024 2096 11033
rect 5908 11024 5960 11076
rect 8668 11024 8720 11076
rect 1952 10956 2004 11008
rect 2872 10999 2924 11008
rect 2872 10965 2881 10999
rect 2881 10965 2915 10999
rect 2915 10965 2924 10999
rect 2872 10956 2924 10965
rect 7012 10956 7064 11008
rect 8116 10956 8168 11008
rect 9404 11024 9456 11076
rect 10600 11024 10652 11076
rect 11152 11024 11204 11076
rect 11888 11092 11940 11144
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 15016 11160 15068 11212
rect 13636 11135 13688 11144
rect 13636 11101 13645 11135
rect 13645 11101 13679 11135
rect 13679 11101 13688 11135
rect 13636 11092 13688 11101
rect 13820 11092 13872 11144
rect 15660 11092 15712 11144
rect 16948 11160 17000 11212
rect 19708 11228 19760 11280
rect 20628 11228 20680 11280
rect 21180 11228 21232 11280
rect 22008 11228 22060 11280
rect 22100 11228 22152 11280
rect 12624 11024 12676 11076
rect 15384 11024 15436 11076
rect 10048 10999 10100 11008
rect 10048 10965 10057 10999
rect 10057 10965 10091 10999
rect 10091 10965 10100 10999
rect 10048 10956 10100 10965
rect 10324 10956 10376 11008
rect 11888 10956 11940 11008
rect 15660 10999 15712 11008
rect 15660 10965 15669 10999
rect 15669 10965 15703 10999
rect 15703 10965 15712 10999
rect 15660 10956 15712 10965
rect 15844 10956 15896 11008
rect 18052 11092 18104 11144
rect 19892 11092 19944 11144
rect 20628 11135 20680 11144
rect 20628 11101 20637 11135
rect 20637 11101 20671 11135
rect 20671 11101 20680 11135
rect 20628 11092 20680 11101
rect 23020 11203 23072 11212
rect 16580 11024 16632 11076
rect 20996 11092 21048 11144
rect 21732 11135 21784 11144
rect 21732 11101 21742 11135
rect 21742 11101 21776 11135
rect 21776 11101 21784 11135
rect 23020 11169 23029 11203
rect 23029 11169 23063 11203
rect 23063 11169 23072 11203
rect 23020 11160 23072 11169
rect 21732 11092 21784 11101
rect 22836 11092 22888 11144
rect 23664 11092 23716 11144
rect 22192 10956 22244 11008
rect 23112 10956 23164 11008
rect 23388 11024 23440 11076
rect 23572 11067 23624 11076
rect 23572 11033 23581 11067
rect 23581 11033 23615 11067
rect 23615 11033 23624 11067
rect 23572 11024 23624 11033
rect 23664 10956 23716 11008
rect 8214 10854 8266 10906
rect 8278 10854 8330 10906
rect 8342 10854 8394 10906
rect 8406 10854 8458 10906
rect 8470 10854 8522 10906
rect 16214 10854 16266 10906
rect 16278 10854 16330 10906
rect 16342 10854 16394 10906
rect 16406 10854 16458 10906
rect 16470 10854 16522 10906
rect 24214 10854 24266 10906
rect 24278 10854 24330 10906
rect 24342 10854 24394 10906
rect 24406 10854 24458 10906
rect 24470 10854 24522 10906
rect 2872 10752 2924 10804
rect 3240 10752 3292 10804
rect 5632 10752 5684 10804
rect 9128 10752 9180 10804
rect 9312 10752 9364 10804
rect 10048 10752 10100 10804
rect 10876 10795 10928 10804
rect 10876 10761 10885 10795
rect 10885 10761 10919 10795
rect 10919 10761 10928 10795
rect 10876 10752 10928 10761
rect 15568 10752 15620 10804
rect 1952 10727 2004 10736
rect 1952 10693 1961 10727
rect 1961 10693 1995 10727
rect 1995 10693 2004 10727
rect 1952 10684 2004 10693
rect 2964 10684 3016 10736
rect 5080 10684 5132 10736
rect 6552 10684 6604 10736
rect 1492 10548 1544 10600
rect 5356 10548 5408 10600
rect 7012 10548 7064 10600
rect 6644 10480 6696 10532
rect 7932 10684 7984 10736
rect 9864 10684 9916 10736
rect 10968 10727 11020 10736
rect 10968 10693 10977 10727
rect 10977 10693 11011 10727
rect 11011 10693 11020 10727
rect 10968 10684 11020 10693
rect 11796 10684 11848 10736
rect 8116 10616 8168 10668
rect 8576 10616 8628 10668
rect 9680 10616 9732 10668
rect 8944 10548 8996 10600
rect 12900 10684 12952 10736
rect 15108 10684 15160 10736
rect 12624 10616 12676 10668
rect 13268 10616 13320 10668
rect 13728 10659 13780 10668
rect 13728 10625 13737 10659
rect 13737 10625 13771 10659
rect 13771 10625 13780 10659
rect 13728 10616 13780 10625
rect 15292 10616 15344 10668
rect 16028 10752 16080 10804
rect 16580 10752 16632 10804
rect 18788 10795 18840 10804
rect 18788 10761 18797 10795
rect 18797 10761 18831 10795
rect 18831 10761 18840 10795
rect 18788 10752 18840 10761
rect 17960 10684 18012 10736
rect 20628 10795 20680 10804
rect 20628 10761 20637 10795
rect 20637 10761 20671 10795
rect 20671 10761 20680 10795
rect 20628 10752 20680 10761
rect 21456 10752 21508 10804
rect 23388 10752 23440 10804
rect 23572 10752 23624 10804
rect 23296 10684 23348 10736
rect 9036 10480 9088 10532
rect 10324 10548 10376 10600
rect 11888 10548 11940 10600
rect 9772 10480 9824 10532
rect 15936 10548 15988 10600
rect 15200 10480 15252 10532
rect 16948 10548 17000 10600
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 21548 10548 21600 10600
rect 22560 10591 22612 10600
rect 22560 10557 22569 10591
rect 22569 10557 22603 10591
rect 22603 10557 22612 10591
rect 22560 10548 22612 10557
rect 23388 10659 23440 10668
rect 23388 10625 23397 10659
rect 23397 10625 23431 10659
rect 23431 10625 23440 10659
rect 23388 10616 23440 10625
rect 23848 10616 23900 10668
rect 23480 10548 23532 10600
rect 22652 10480 22704 10532
rect 5448 10412 5500 10464
rect 5816 10412 5868 10464
rect 7288 10412 7340 10464
rect 7840 10412 7892 10464
rect 7932 10455 7984 10464
rect 7932 10421 7941 10455
rect 7941 10421 7975 10455
rect 7975 10421 7984 10455
rect 7932 10412 7984 10421
rect 13360 10455 13412 10464
rect 13360 10421 13369 10455
rect 13369 10421 13403 10455
rect 13403 10421 13412 10455
rect 13360 10412 13412 10421
rect 21916 10455 21968 10464
rect 21916 10421 21925 10455
rect 21925 10421 21959 10455
rect 21959 10421 21968 10455
rect 21916 10412 21968 10421
rect 22836 10412 22888 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 12214 10310 12266 10362
rect 12278 10310 12330 10362
rect 12342 10310 12394 10362
rect 12406 10310 12458 10362
rect 12470 10310 12522 10362
rect 20214 10310 20266 10362
rect 20278 10310 20330 10362
rect 20342 10310 20394 10362
rect 20406 10310 20458 10362
rect 20470 10310 20522 10362
rect 1952 10208 2004 10260
rect 2504 10072 2556 10124
rect 1492 10004 1544 10056
rect 2964 9936 3016 9988
rect 4712 10208 4764 10260
rect 5080 10251 5132 10260
rect 5080 10217 5089 10251
rect 5089 10217 5123 10251
rect 5123 10217 5132 10251
rect 5080 10208 5132 10217
rect 5356 10251 5408 10260
rect 5356 10217 5365 10251
rect 5365 10217 5399 10251
rect 5399 10217 5408 10251
rect 5356 10208 5408 10217
rect 7288 10208 7340 10260
rect 8576 10208 8628 10260
rect 12624 10251 12676 10260
rect 12624 10217 12633 10251
rect 12633 10217 12667 10251
rect 12667 10217 12676 10251
rect 12624 10208 12676 10217
rect 13268 10208 13320 10260
rect 17316 10208 17368 10260
rect 17592 10208 17644 10260
rect 6552 10140 6604 10192
rect 13544 10140 13596 10192
rect 15660 10140 15712 10192
rect 18052 10208 18104 10260
rect 18512 10251 18564 10260
rect 18512 10217 18521 10251
rect 18521 10217 18555 10251
rect 18555 10217 18564 10251
rect 18512 10208 18564 10217
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 2872 9868 2924 9920
rect 4620 9868 4672 9920
rect 5448 9868 5500 9920
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 7564 10072 7616 10124
rect 10324 10072 10376 10124
rect 6644 10047 6696 10056
rect 6644 10013 6653 10047
rect 6653 10013 6687 10047
rect 6687 10013 6696 10047
rect 6644 10004 6696 10013
rect 10876 10072 10928 10124
rect 13360 10072 13412 10124
rect 13636 10072 13688 10124
rect 6920 9979 6972 9988
rect 6920 9945 6929 9979
rect 6929 9945 6963 9979
rect 6963 9945 6972 9979
rect 6920 9936 6972 9945
rect 7932 9936 7984 9988
rect 9220 9936 9272 9988
rect 9312 9979 9364 9988
rect 9312 9945 9321 9979
rect 9321 9945 9355 9979
rect 9355 9945 9364 9979
rect 9312 9936 9364 9945
rect 9772 9936 9824 9988
rect 10968 9936 11020 9988
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 14004 10004 14056 10056
rect 15292 10115 15344 10124
rect 15292 10081 15301 10115
rect 15301 10081 15335 10115
rect 15335 10081 15344 10115
rect 15292 10072 15344 10081
rect 7104 9868 7156 9920
rect 10232 9868 10284 9920
rect 13820 9936 13872 9988
rect 12624 9868 12676 9920
rect 12900 9868 12952 9920
rect 15384 10047 15436 10056
rect 15384 10013 15393 10047
rect 15393 10013 15427 10047
rect 15427 10013 15436 10047
rect 15384 10004 15436 10013
rect 19892 10072 19944 10124
rect 22652 10208 22704 10260
rect 23296 10208 23348 10260
rect 24032 10208 24084 10260
rect 22468 10072 22520 10124
rect 22928 10072 22980 10124
rect 23112 10072 23164 10124
rect 16672 10004 16724 10056
rect 20628 10004 20680 10056
rect 23572 10004 23624 10056
rect 15292 9936 15344 9988
rect 17500 9979 17552 9988
rect 17500 9945 17509 9979
rect 17509 9945 17543 9979
rect 17543 9945 17552 9979
rect 17500 9936 17552 9945
rect 19800 9936 19852 9988
rect 15752 9868 15804 9920
rect 17684 9911 17736 9920
rect 17684 9877 17709 9911
rect 17709 9877 17736 9911
rect 17684 9868 17736 9877
rect 19616 9868 19668 9920
rect 19984 9868 20036 9920
rect 21548 9936 21600 9988
rect 21916 9979 21968 9988
rect 21916 9945 21925 9979
rect 21925 9945 21959 9979
rect 21959 9945 21968 9979
rect 21916 9936 21968 9945
rect 22652 9936 22704 9988
rect 21640 9868 21692 9920
rect 22100 9868 22152 9920
rect 8214 9766 8266 9818
rect 8278 9766 8330 9818
rect 8342 9766 8394 9818
rect 8406 9766 8458 9818
rect 8470 9766 8522 9818
rect 16214 9766 16266 9818
rect 16278 9766 16330 9818
rect 16342 9766 16394 9818
rect 16406 9766 16458 9818
rect 16470 9766 16522 9818
rect 24214 9766 24266 9818
rect 24278 9766 24330 9818
rect 24342 9766 24394 9818
rect 24406 9766 24458 9818
rect 24470 9766 24522 9818
rect 1860 9639 1912 9648
rect 1860 9605 1869 9639
rect 1869 9605 1903 9639
rect 1903 9605 1912 9639
rect 1860 9596 1912 9605
rect 2044 9639 2096 9648
rect 2044 9605 2069 9639
rect 2069 9605 2096 9639
rect 2504 9707 2556 9716
rect 2504 9673 2513 9707
rect 2513 9673 2547 9707
rect 2547 9673 2556 9707
rect 2504 9664 2556 9673
rect 2872 9707 2924 9716
rect 2872 9673 2881 9707
rect 2881 9673 2915 9707
rect 2915 9673 2924 9707
rect 2872 9664 2924 9673
rect 6920 9707 6972 9716
rect 6920 9673 6929 9707
rect 6929 9673 6963 9707
rect 6963 9673 6972 9707
rect 6920 9664 6972 9673
rect 7472 9664 7524 9716
rect 9036 9664 9088 9716
rect 10232 9664 10284 9716
rect 2044 9596 2096 9605
rect 2964 9596 3016 9648
rect 4988 9596 5040 9648
rect 6276 9596 6328 9648
rect 3240 9528 3292 9580
rect 6552 9528 6604 9580
rect 8944 9639 8996 9648
rect 8944 9605 8953 9639
rect 8953 9605 8987 9639
rect 8987 9605 8996 9639
rect 8944 9596 8996 9605
rect 9128 9639 9180 9648
rect 9128 9605 9153 9639
rect 9153 9605 9180 9639
rect 9128 9596 9180 9605
rect 7104 9571 7156 9580
rect 7104 9537 7113 9571
rect 7113 9537 7147 9571
rect 7147 9537 7156 9571
rect 7104 9528 7156 9537
rect 7472 9528 7524 9580
rect 9864 9528 9916 9580
rect 10324 9528 10376 9580
rect 10876 9571 10928 9580
rect 10876 9537 10885 9571
rect 10885 9537 10919 9571
rect 10919 9537 10928 9571
rect 10876 9528 10928 9537
rect 3148 9503 3200 9512
rect 3148 9469 3157 9503
rect 3157 9469 3191 9503
rect 3191 9469 3200 9503
rect 3148 9460 3200 9469
rect 1492 9392 1544 9444
rect 5264 9460 5316 9512
rect 5908 9460 5960 9512
rect 6368 9460 6420 9512
rect 7564 9460 7616 9512
rect 7840 9460 7892 9512
rect 10416 9460 10468 9512
rect 11520 9528 11572 9580
rect 12072 9528 12124 9580
rect 2136 9324 2188 9376
rect 6644 9392 6696 9444
rect 9772 9392 9824 9444
rect 5816 9324 5868 9376
rect 7380 9324 7432 9376
rect 8760 9324 8812 9376
rect 10508 9367 10560 9376
rect 10508 9333 10517 9367
rect 10517 9333 10551 9367
rect 10551 9333 10560 9367
rect 10508 9324 10560 9333
rect 11244 9503 11296 9512
rect 11244 9469 11253 9503
rect 11253 9469 11287 9503
rect 11287 9469 11296 9503
rect 11244 9460 11296 9469
rect 12624 9707 12676 9716
rect 12624 9673 12633 9707
rect 12633 9673 12667 9707
rect 12667 9673 12676 9707
rect 12624 9664 12676 9673
rect 13268 9664 13320 9716
rect 15752 9664 15804 9716
rect 12716 9528 12768 9580
rect 14004 9571 14056 9580
rect 14004 9537 14013 9571
rect 14013 9537 14047 9571
rect 14047 9537 14056 9571
rect 14004 9528 14056 9537
rect 14648 9596 14700 9648
rect 14464 9571 14516 9580
rect 14464 9537 14473 9571
rect 14473 9537 14507 9571
rect 14507 9537 14516 9571
rect 14464 9528 14516 9537
rect 15292 9528 15344 9580
rect 18052 9596 18104 9648
rect 18604 9596 18656 9648
rect 22192 9664 22244 9716
rect 22468 9664 22520 9716
rect 22560 9664 22612 9716
rect 23756 9664 23808 9716
rect 22100 9639 22152 9648
rect 12900 9392 12952 9444
rect 15108 9392 15160 9444
rect 13452 9367 13504 9376
rect 13452 9333 13461 9367
rect 13461 9333 13495 9367
rect 13495 9333 13504 9367
rect 13452 9324 13504 9333
rect 13728 9324 13780 9376
rect 15660 9528 15712 9580
rect 16120 9528 16172 9580
rect 18696 9528 18748 9580
rect 18880 9528 18932 9580
rect 19340 9528 19392 9580
rect 22100 9605 22127 9639
rect 22127 9605 22152 9639
rect 22100 9596 22152 9605
rect 15752 9503 15804 9512
rect 15752 9469 15761 9503
rect 15761 9469 15795 9503
rect 15795 9469 15804 9503
rect 15752 9460 15804 9469
rect 15844 9460 15896 9512
rect 18236 9460 18288 9512
rect 19984 9503 20036 9512
rect 19984 9469 19993 9503
rect 19993 9469 20027 9503
rect 20027 9469 20036 9503
rect 19984 9460 20036 9469
rect 21364 9528 21416 9580
rect 22836 9639 22888 9648
rect 22836 9605 22845 9639
rect 22845 9605 22879 9639
rect 22879 9605 22888 9639
rect 22836 9596 22888 9605
rect 23480 9596 23532 9648
rect 21548 9460 21600 9512
rect 23388 9460 23440 9512
rect 16580 9324 16632 9376
rect 17224 9324 17276 9376
rect 18788 9367 18840 9376
rect 18788 9333 18797 9367
rect 18797 9333 18831 9367
rect 18831 9333 18840 9367
rect 18788 9324 18840 9333
rect 18972 9367 19024 9376
rect 18972 9333 18981 9367
rect 18981 9333 19015 9367
rect 19015 9333 19024 9367
rect 18972 9324 19024 9333
rect 22284 9324 22336 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 12214 9222 12266 9274
rect 12278 9222 12330 9274
rect 12342 9222 12394 9274
rect 12406 9222 12458 9274
rect 12470 9222 12522 9274
rect 20214 9222 20266 9274
rect 20278 9222 20330 9274
rect 20342 9222 20394 9274
rect 20406 9222 20458 9274
rect 20470 9222 20522 9274
rect 4804 9163 4856 9172
rect 4804 9129 4813 9163
rect 4813 9129 4847 9163
rect 4847 9129 4856 9163
rect 4804 9120 4856 9129
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 5264 9163 5316 9172
rect 5264 9129 5273 9163
rect 5273 9129 5307 9163
rect 5307 9129 5316 9163
rect 5264 9120 5316 9129
rect 5356 9120 5408 9172
rect 1492 8916 1544 8968
rect 2136 8848 2188 8900
rect 8024 9052 8076 9104
rect 5448 8959 5500 8968
rect 5448 8925 5457 8959
rect 5457 8925 5491 8959
rect 5491 8925 5500 8959
rect 5448 8916 5500 8925
rect 5632 8984 5684 9036
rect 5816 8916 5868 8968
rect 6368 8959 6420 8968
rect 6368 8925 6377 8959
rect 6377 8925 6411 8959
rect 6411 8925 6420 8959
rect 6368 8916 6420 8925
rect 6460 8916 6512 8968
rect 7196 8984 7248 9036
rect 7472 8959 7524 8968
rect 7472 8925 7481 8959
rect 7481 8925 7515 8959
rect 7515 8925 7524 8959
rect 7472 8916 7524 8925
rect 2228 8780 2280 8832
rect 2504 8780 2556 8832
rect 4712 8848 4764 8900
rect 5356 8848 5408 8900
rect 3332 8823 3384 8832
rect 3332 8789 3341 8823
rect 3341 8789 3375 8823
rect 3375 8789 3384 8823
rect 3332 8780 3384 8789
rect 5540 8780 5592 8832
rect 6920 8780 6972 8832
rect 7104 8848 7156 8900
rect 7380 8891 7432 8900
rect 7380 8857 7389 8891
rect 7389 8857 7423 8891
rect 7423 8857 7432 8891
rect 7380 8848 7432 8857
rect 7840 8848 7892 8900
rect 8024 8848 8076 8900
rect 8668 9120 8720 9172
rect 9312 9120 9364 9172
rect 10508 9120 10560 9172
rect 18052 9163 18104 9172
rect 18052 9129 18061 9163
rect 18061 9129 18095 9163
rect 18095 9129 18104 9163
rect 18052 9120 18104 9129
rect 18972 9120 19024 9172
rect 19800 9120 19852 9172
rect 13452 9052 13504 9104
rect 9404 8959 9456 8968
rect 9404 8925 9413 8959
rect 9413 8925 9447 8959
rect 9447 8925 9456 8959
rect 9404 8916 9456 8925
rect 11244 8984 11296 9036
rect 15200 8984 15252 9036
rect 16948 8984 17000 9036
rect 19340 9027 19392 9036
rect 19340 8993 19349 9027
rect 19349 8993 19383 9027
rect 19383 8993 19392 9027
rect 19340 8984 19392 8993
rect 19616 8984 19668 9036
rect 22376 9120 22428 9172
rect 21916 9052 21968 9104
rect 22652 9120 22704 9172
rect 23204 9120 23256 9172
rect 23480 9163 23532 9172
rect 23480 9129 23489 9163
rect 23489 9129 23523 9163
rect 23523 9129 23532 9163
rect 23480 9120 23532 9129
rect 23664 9120 23716 9172
rect 10876 8916 10928 8968
rect 11060 8916 11112 8968
rect 12072 8916 12124 8968
rect 12716 8916 12768 8968
rect 10324 8891 10376 8900
rect 10324 8857 10333 8891
rect 10333 8857 10367 8891
rect 10367 8857 10376 8891
rect 10324 8848 10376 8857
rect 10416 8891 10468 8900
rect 10416 8857 10425 8891
rect 10425 8857 10459 8891
rect 10459 8857 10468 8891
rect 10416 8848 10468 8857
rect 10508 8848 10560 8900
rect 14096 8916 14148 8968
rect 14188 8959 14240 8968
rect 14188 8925 14197 8959
rect 14197 8925 14231 8959
rect 14231 8925 14240 8959
rect 14188 8916 14240 8925
rect 21456 8916 21508 8968
rect 7748 8780 7800 8832
rect 8760 8780 8812 8832
rect 9864 8780 9916 8832
rect 12992 8780 13044 8832
rect 14372 8848 14424 8900
rect 15200 8848 15252 8900
rect 16580 8891 16632 8900
rect 16580 8857 16589 8891
rect 16589 8857 16623 8891
rect 16623 8857 16632 8891
rect 16580 8848 16632 8857
rect 14648 8780 14700 8832
rect 14740 8780 14792 8832
rect 18880 8848 18932 8900
rect 19340 8848 19392 8900
rect 20076 8848 20128 8900
rect 18604 8780 18656 8832
rect 19708 8780 19760 8832
rect 20628 8780 20680 8832
rect 21272 8780 21324 8832
rect 21824 8916 21876 8968
rect 24124 8959 24176 8968
rect 24124 8925 24133 8959
rect 24133 8925 24167 8959
rect 24167 8925 24176 8959
rect 24124 8916 24176 8925
rect 24676 8848 24728 8900
rect 8214 8678 8266 8730
rect 8278 8678 8330 8730
rect 8342 8678 8394 8730
rect 8406 8678 8458 8730
rect 8470 8678 8522 8730
rect 16214 8678 16266 8730
rect 16278 8678 16330 8730
rect 16342 8678 16394 8730
rect 16406 8678 16458 8730
rect 16470 8678 16522 8730
rect 24214 8678 24266 8730
rect 24278 8678 24330 8730
rect 24342 8678 24394 8730
rect 24406 8678 24458 8730
rect 24470 8678 24522 8730
rect 2136 8619 2188 8628
rect 2136 8585 2145 8619
rect 2145 8585 2179 8619
rect 2179 8585 2188 8619
rect 2136 8576 2188 8585
rect 2228 8576 2280 8628
rect 2872 8576 2924 8628
rect 3332 8576 3384 8628
rect 1584 8508 1636 8560
rect 4712 8576 4764 8628
rect 3608 8508 3660 8560
rect 6368 8576 6420 8628
rect 6644 8576 6696 8628
rect 2136 8440 2188 8492
rect 2780 8440 2832 8492
rect 3424 8483 3476 8492
rect 3424 8449 3433 8483
rect 3433 8449 3467 8483
rect 3467 8449 3476 8483
rect 3424 8440 3476 8449
rect 6460 8508 6512 8560
rect 7288 8508 7340 8560
rect 6368 8440 6420 8492
rect 6828 8483 6880 8492
rect 6828 8449 6837 8483
rect 6837 8449 6871 8483
rect 6871 8449 6880 8483
rect 6828 8440 6880 8449
rect 6920 8483 6972 8492
rect 6920 8449 6929 8483
rect 6929 8449 6963 8483
rect 6963 8449 6972 8483
rect 6920 8440 6972 8449
rect 7012 8483 7064 8492
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 9220 8576 9272 8628
rect 10876 8576 10928 8628
rect 14372 8619 14424 8628
rect 14372 8585 14381 8619
rect 14381 8585 14415 8619
rect 14415 8585 14424 8619
rect 14372 8576 14424 8585
rect 15200 8619 15252 8628
rect 15200 8585 15209 8619
rect 15209 8585 15243 8619
rect 15243 8585 15252 8619
rect 15200 8576 15252 8585
rect 7748 8551 7800 8560
rect 7748 8517 7757 8551
rect 7757 8517 7791 8551
rect 7791 8517 7800 8551
rect 7748 8508 7800 8517
rect 8760 8508 8812 8560
rect 10232 8508 10284 8560
rect 10324 8508 10376 8560
rect 15844 8576 15896 8628
rect 18696 8619 18748 8628
rect 18696 8585 18705 8619
rect 18705 8585 18739 8619
rect 18739 8585 18748 8619
rect 18696 8576 18748 8585
rect 3148 8372 3200 8424
rect 3792 8304 3844 8356
rect 6460 8304 6512 8356
rect 7196 8415 7248 8424
rect 7196 8381 7205 8415
rect 7205 8381 7239 8415
rect 7239 8381 7248 8415
rect 7196 8372 7248 8381
rect 6920 8304 6972 8356
rect 10416 8483 10468 8492
rect 10416 8449 10425 8483
rect 10425 8449 10459 8483
rect 10459 8449 10468 8483
rect 10416 8440 10468 8449
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 10784 8483 10836 8492
rect 10784 8449 10793 8483
rect 10793 8449 10827 8483
rect 10827 8449 10836 8483
rect 10784 8440 10836 8449
rect 11060 8372 11112 8424
rect 11888 8483 11940 8492
rect 11888 8449 11897 8483
rect 11897 8449 11931 8483
rect 11931 8449 11940 8483
rect 11888 8440 11940 8449
rect 11980 8440 12032 8492
rect 12624 8440 12676 8492
rect 12808 8440 12860 8492
rect 13820 8440 13872 8492
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 15108 8440 15160 8492
rect 15476 8508 15528 8560
rect 16672 8508 16724 8560
rect 17224 8551 17276 8560
rect 17224 8517 17233 8551
rect 17233 8517 17267 8551
rect 17267 8517 17276 8551
rect 17224 8508 17276 8517
rect 18788 8508 18840 8560
rect 19340 8619 19392 8628
rect 19340 8585 19349 8619
rect 19349 8585 19383 8619
rect 19383 8585 19392 8619
rect 19340 8576 19392 8585
rect 19708 8619 19760 8628
rect 19708 8585 19717 8619
rect 19717 8585 19751 8619
rect 19751 8585 19760 8619
rect 19708 8576 19760 8585
rect 20076 8576 20128 8628
rect 21548 8576 21600 8628
rect 15752 8440 15804 8492
rect 20996 8551 21048 8560
rect 20996 8517 21005 8551
rect 21005 8517 21039 8551
rect 21039 8517 21048 8551
rect 20996 8508 21048 8517
rect 21732 8508 21784 8560
rect 11704 8304 11756 8356
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 14648 8415 14700 8424
rect 14648 8381 14657 8415
rect 14657 8381 14691 8415
rect 14691 8381 14700 8415
rect 21088 8440 21140 8492
rect 21364 8440 21416 8492
rect 22192 8508 22244 8560
rect 24676 8508 24728 8560
rect 14648 8372 14700 8381
rect 16120 8415 16172 8424
rect 16120 8381 16129 8415
rect 16129 8381 16163 8415
rect 16163 8381 16172 8415
rect 16120 8372 16172 8381
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 19708 8372 19760 8424
rect 19892 8415 19944 8424
rect 19892 8381 19901 8415
rect 19901 8381 19935 8415
rect 19935 8381 19944 8415
rect 19892 8372 19944 8381
rect 22284 8415 22336 8424
rect 22284 8381 22293 8415
rect 22293 8381 22327 8415
rect 22327 8381 22336 8415
rect 22284 8372 22336 8381
rect 15936 8347 15988 8356
rect 15936 8313 15945 8347
rect 15945 8313 15979 8347
rect 15979 8313 15988 8347
rect 15936 8304 15988 8313
rect 18788 8304 18840 8356
rect 1952 8279 2004 8288
rect 1952 8245 1961 8279
rect 1961 8245 1995 8279
rect 1995 8245 2004 8279
rect 1952 8236 2004 8245
rect 5540 8236 5592 8288
rect 6552 8236 6604 8288
rect 7288 8236 7340 8288
rect 10048 8236 10100 8288
rect 13452 8236 13504 8288
rect 13544 8236 13596 8288
rect 15016 8236 15068 8288
rect 16580 8236 16632 8288
rect 18880 8236 18932 8288
rect 20996 8304 21048 8356
rect 21364 8347 21416 8356
rect 21364 8313 21373 8347
rect 21373 8313 21407 8347
rect 21407 8313 21416 8347
rect 21364 8304 21416 8313
rect 23296 8304 23348 8356
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 21180 8236 21232 8245
rect 21640 8236 21692 8288
rect 23664 8236 23716 8288
rect 23848 8236 23900 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 12214 8134 12266 8186
rect 12278 8134 12330 8186
rect 12342 8134 12394 8186
rect 12406 8134 12458 8186
rect 12470 8134 12522 8186
rect 20214 8134 20266 8186
rect 20278 8134 20330 8186
rect 20342 8134 20394 8186
rect 20406 8134 20458 8186
rect 20470 8134 20522 8186
rect 1676 8075 1728 8084
rect 1676 8041 1685 8075
rect 1685 8041 1719 8075
rect 1719 8041 1728 8075
rect 1676 8032 1728 8041
rect 3148 8032 3200 8084
rect 6276 8032 6328 8084
rect 7104 8032 7156 8084
rect 7196 8032 7248 8084
rect 7472 8032 7524 8084
rect 7564 8032 7616 8084
rect 10508 8032 10560 8084
rect 11060 8032 11112 8084
rect 11980 8032 12032 8084
rect 12900 8032 12952 8084
rect 15936 8032 15988 8084
rect 16580 8032 16632 8084
rect 17684 8032 17736 8084
rect 18972 8032 19024 8084
rect 19524 8032 19576 8084
rect 2872 7939 2924 7948
rect 2872 7905 2881 7939
rect 2881 7905 2915 7939
rect 2915 7905 2924 7939
rect 2872 7896 2924 7905
rect 3148 7896 3200 7948
rect 3608 7896 3660 7948
rect 4068 7896 4120 7948
rect 6644 7896 6696 7948
rect 1400 7828 1452 7880
rect 1676 7828 1728 7880
rect 2688 7828 2740 7880
rect 6552 7828 6604 7880
rect 7288 7964 7340 8016
rect 7748 7964 7800 8016
rect 11152 7964 11204 8016
rect 7932 7896 7984 7948
rect 7104 7828 7156 7880
rect 4620 7760 4672 7812
rect 1768 7692 1820 7744
rect 2412 7735 2464 7744
rect 2412 7701 2421 7735
rect 2421 7701 2455 7735
rect 2455 7701 2464 7735
rect 2412 7692 2464 7701
rect 3240 7692 3292 7744
rect 6460 7692 6512 7744
rect 7840 7828 7892 7880
rect 8116 7828 8168 7880
rect 7656 7692 7708 7744
rect 9036 7871 9088 7880
rect 9036 7837 9045 7871
rect 9045 7837 9079 7871
rect 9079 7837 9088 7871
rect 9036 7828 9088 7837
rect 9588 7828 9640 7880
rect 11336 7896 11388 7948
rect 13728 7964 13780 8016
rect 12808 7896 12860 7948
rect 10692 7760 10744 7812
rect 9496 7692 9548 7744
rect 11060 7871 11112 7880
rect 11060 7837 11069 7871
rect 11069 7837 11103 7871
rect 11103 7837 11112 7871
rect 11060 7828 11112 7837
rect 11704 7828 11756 7880
rect 11888 7871 11940 7880
rect 11888 7837 11897 7871
rect 11897 7837 11931 7871
rect 11931 7837 11940 7871
rect 11888 7828 11940 7837
rect 12624 7828 12676 7880
rect 13176 7871 13228 7880
rect 13176 7837 13185 7871
rect 13185 7837 13219 7871
rect 13219 7837 13228 7871
rect 13176 7828 13228 7837
rect 13452 7896 13504 7948
rect 14924 7896 14976 7948
rect 15476 7896 15528 7948
rect 13728 7828 13780 7880
rect 14096 7828 14148 7880
rect 14188 7871 14240 7880
rect 14188 7837 14197 7871
rect 14197 7837 14231 7871
rect 14231 7837 14240 7871
rect 14188 7828 14240 7837
rect 19616 7964 19668 8016
rect 21180 8032 21232 8084
rect 21916 7964 21968 8016
rect 22284 8032 22336 8084
rect 23848 7964 23900 8016
rect 17500 7896 17552 7948
rect 18236 7939 18288 7948
rect 18236 7905 18245 7939
rect 18245 7905 18279 7939
rect 18279 7905 18288 7939
rect 18236 7896 18288 7905
rect 18696 7896 18748 7948
rect 17592 7828 17644 7880
rect 19708 7896 19760 7948
rect 22100 7896 22152 7948
rect 22652 7896 22704 7948
rect 23388 7939 23440 7948
rect 23388 7905 23397 7939
rect 23397 7905 23431 7939
rect 23431 7905 23440 7939
rect 23388 7896 23440 7905
rect 11704 7692 11756 7744
rect 14740 7760 14792 7812
rect 15752 7760 15804 7812
rect 15844 7692 15896 7744
rect 18696 7760 18748 7812
rect 18880 7760 18932 7812
rect 17132 7692 17184 7744
rect 17408 7692 17460 7744
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 18512 7692 18564 7744
rect 19432 7692 19484 7744
rect 23296 7871 23348 7880
rect 23296 7837 23305 7871
rect 23305 7837 23339 7871
rect 23339 7837 23348 7871
rect 23296 7828 23348 7837
rect 20812 7760 20864 7812
rect 22100 7760 22152 7812
rect 22928 7760 22980 7812
rect 23020 7760 23072 7812
rect 23664 7828 23716 7880
rect 24124 7871 24176 7880
rect 24124 7837 24133 7871
rect 24133 7837 24167 7871
rect 24167 7837 24176 7871
rect 24124 7828 24176 7837
rect 19800 7735 19852 7744
rect 19800 7701 19809 7735
rect 19809 7701 19843 7735
rect 19843 7701 19852 7735
rect 19800 7692 19852 7701
rect 20076 7692 20128 7744
rect 20904 7735 20956 7744
rect 20904 7701 20913 7735
rect 20913 7701 20947 7735
rect 20947 7701 20956 7735
rect 20904 7692 20956 7701
rect 21824 7692 21876 7744
rect 22560 7692 22612 7744
rect 22744 7692 22796 7744
rect 8214 7590 8266 7642
rect 8278 7590 8330 7642
rect 8342 7590 8394 7642
rect 8406 7590 8458 7642
rect 8470 7590 8522 7642
rect 16214 7590 16266 7642
rect 16278 7590 16330 7642
rect 16342 7590 16394 7642
rect 16406 7590 16458 7642
rect 16470 7590 16522 7642
rect 24214 7590 24266 7642
rect 24278 7590 24330 7642
rect 24342 7590 24394 7642
rect 24406 7590 24458 7642
rect 24470 7590 24522 7642
rect 2412 7488 2464 7540
rect 3240 7531 3292 7540
rect 3240 7497 3249 7531
rect 3249 7497 3283 7531
rect 3283 7497 3292 7531
rect 3240 7488 3292 7497
rect 4620 7488 4672 7540
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 7932 7531 7984 7540
rect 7932 7497 7941 7531
rect 7941 7497 7975 7531
rect 7975 7497 7984 7531
rect 7932 7488 7984 7497
rect 8116 7488 8168 7540
rect 12716 7488 12768 7540
rect 12992 7531 13044 7540
rect 12992 7497 13019 7531
rect 13019 7497 13044 7531
rect 2872 7352 2924 7404
rect 3792 7395 3844 7404
rect 3792 7361 3800 7395
rect 3800 7361 3834 7395
rect 3834 7361 3844 7395
rect 3792 7352 3844 7361
rect 3976 7352 4028 7404
rect 1492 7327 1544 7336
rect 1492 7293 1501 7327
rect 1501 7293 1535 7327
rect 1535 7293 1544 7327
rect 1492 7284 1544 7293
rect 2504 7284 2556 7336
rect 5816 7420 5868 7472
rect 6552 7420 6604 7472
rect 4712 7352 4764 7404
rect 5080 7352 5132 7404
rect 5172 7395 5224 7404
rect 5172 7361 5181 7395
rect 5181 7361 5215 7395
rect 5215 7361 5224 7395
rect 5172 7352 5224 7361
rect 5908 7395 5960 7404
rect 5908 7361 5917 7395
rect 5917 7361 5951 7395
rect 5951 7361 5960 7395
rect 5908 7352 5960 7361
rect 6092 7395 6144 7404
rect 6092 7361 6101 7395
rect 6101 7361 6135 7395
rect 6135 7361 6144 7395
rect 6092 7352 6144 7361
rect 6644 7395 6696 7404
rect 6644 7361 6653 7395
rect 6653 7361 6687 7395
rect 6687 7361 6696 7395
rect 6644 7352 6696 7361
rect 5632 7327 5684 7336
rect 5632 7293 5641 7327
rect 5641 7293 5675 7327
rect 5675 7293 5684 7327
rect 6828 7352 6880 7404
rect 7656 7463 7708 7472
rect 7656 7429 7665 7463
rect 7665 7429 7699 7463
rect 7699 7429 7708 7463
rect 7656 7420 7708 7429
rect 5632 7284 5684 7293
rect 3148 7216 3200 7268
rect 1952 7148 2004 7200
rect 4804 7216 4856 7268
rect 6368 7216 6420 7268
rect 8668 7420 8720 7472
rect 8760 7352 8812 7404
rect 4896 7191 4948 7200
rect 4896 7157 4905 7191
rect 4905 7157 4939 7191
rect 4939 7157 4948 7191
rect 4896 7148 4948 7157
rect 5356 7191 5408 7200
rect 5356 7157 5365 7191
rect 5365 7157 5399 7191
rect 5399 7157 5408 7191
rect 5356 7148 5408 7157
rect 5724 7148 5776 7200
rect 6736 7148 6788 7200
rect 6920 7148 6972 7200
rect 8576 7148 8628 7200
rect 8668 7191 8720 7200
rect 8668 7157 8677 7191
rect 8677 7157 8711 7191
rect 8711 7157 8720 7191
rect 8668 7148 8720 7157
rect 9496 7463 9548 7472
rect 9496 7429 9505 7463
rect 9505 7429 9539 7463
rect 9539 7429 9548 7463
rect 9496 7420 9548 7429
rect 12992 7488 13044 7497
rect 14280 7463 14332 7472
rect 14280 7429 14289 7463
rect 14289 7429 14323 7463
rect 14323 7429 14332 7463
rect 14280 7420 14332 7429
rect 14464 7463 14516 7472
rect 14464 7429 14489 7463
rect 14489 7429 14516 7463
rect 14740 7488 14792 7540
rect 14464 7420 14516 7429
rect 14924 7463 14976 7472
rect 14924 7429 14933 7463
rect 14933 7429 14967 7463
rect 14967 7429 14976 7463
rect 14924 7420 14976 7429
rect 15108 7463 15160 7472
rect 15108 7429 15133 7463
rect 15133 7429 15160 7463
rect 15108 7420 15160 7429
rect 15384 7420 15436 7472
rect 16028 7420 16080 7472
rect 9220 7327 9272 7336
rect 9220 7293 9229 7327
rect 9229 7293 9263 7327
rect 9263 7293 9272 7327
rect 9220 7284 9272 7293
rect 9588 7284 9640 7336
rect 9864 7284 9916 7336
rect 11612 7327 11664 7336
rect 11612 7293 11621 7327
rect 11621 7293 11655 7327
rect 11655 7293 11664 7327
rect 11612 7284 11664 7293
rect 11888 7327 11940 7336
rect 11888 7293 11897 7327
rect 11897 7293 11931 7327
rect 11931 7293 11940 7327
rect 11888 7284 11940 7293
rect 10508 7216 10560 7268
rect 13544 7395 13596 7404
rect 13544 7361 13553 7395
rect 13553 7361 13587 7395
rect 13587 7361 13596 7395
rect 13544 7352 13596 7361
rect 13728 7352 13780 7404
rect 16120 7352 16172 7404
rect 17408 7463 17460 7472
rect 17408 7429 17417 7463
rect 17417 7429 17451 7463
rect 17451 7429 17460 7463
rect 17408 7420 17460 7429
rect 19800 7488 19852 7540
rect 20812 7488 20864 7540
rect 19340 7420 19392 7472
rect 19432 7463 19484 7472
rect 19432 7429 19441 7463
rect 19441 7429 19475 7463
rect 19475 7429 19484 7463
rect 19432 7420 19484 7429
rect 12716 7284 12768 7336
rect 15108 7284 15160 7336
rect 15292 7284 15344 7336
rect 18512 7352 18564 7404
rect 16948 7284 17000 7336
rect 21732 7420 21784 7472
rect 22560 7463 22612 7472
rect 22560 7429 22569 7463
rect 22569 7429 22603 7463
rect 22603 7429 22612 7463
rect 22560 7420 22612 7429
rect 24032 7420 24084 7472
rect 22192 7352 22244 7404
rect 15016 7148 15068 7200
rect 15200 7148 15252 7200
rect 15568 7191 15620 7200
rect 15568 7157 15577 7191
rect 15577 7157 15611 7191
rect 15611 7157 15620 7191
rect 15568 7148 15620 7157
rect 22652 7284 22704 7336
rect 22928 7284 22980 7336
rect 15936 7148 15988 7200
rect 19248 7148 19300 7200
rect 21456 7148 21508 7200
rect 22376 7148 22428 7200
rect 23296 7148 23348 7200
rect 24584 7148 24636 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 12214 7046 12266 7098
rect 12278 7046 12330 7098
rect 12342 7046 12394 7098
rect 12406 7046 12458 7098
rect 12470 7046 12522 7098
rect 20214 7046 20266 7098
rect 20278 7046 20330 7098
rect 20342 7046 20394 7098
rect 20406 7046 20458 7098
rect 20470 7046 20522 7098
rect 1952 6944 2004 6996
rect 6092 6944 6144 6996
rect 8024 6944 8076 6996
rect 10508 6944 10560 6996
rect 3056 6876 3108 6928
rect 5816 6876 5868 6928
rect 1584 6672 1636 6724
rect 2504 6740 2556 6792
rect 3792 6808 3844 6860
rect 5632 6808 5684 6860
rect 6092 6808 6144 6860
rect 9680 6876 9732 6928
rect 16028 6944 16080 6996
rect 18052 6944 18104 6996
rect 18972 6944 19024 6996
rect 19616 6987 19668 6996
rect 19616 6953 19625 6987
rect 19625 6953 19659 6987
rect 19659 6953 19668 6987
rect 19616 6944 19668 6953
rect 20076 6944 20128 6996
rect 20904 6944 20956 6996
rect 12072 6876 12124 6928
rect 2136 6672 2188 6724
rect 2872 6672 2924 6724
rect 3056 6715 3108 6724
rect 3056 6681 3065 6715
rect 3065 6681 3099 6715
rect 3099 6681 3108 6715
rect 3056 6672 3108 6681
rect 2780 6647 2832 6656
rect 2780 6613 2789 6647
rect 2789 6613 2823 6647
rect 2823 6613 2832 6647
rect 2780 6604 2832 6613
rect 3516 6647 3568 6656
rect 3516 6613 3525 6647
rect 3525 6613 3559 6647
rect 3559 6613 3568 6647
rect 3516 6604 3568 6613
rect 3792 6672 3844 6724
rect 5908 6740 5960 6792
rect 6736 6808 6788 6860
rect 3976 6604 4028 6656
rect 5540 6604 5592 6656
rect 5816 6672 5868 6724
rect 6552 6672 6604 6724
rect 7840 6740 7892 6792
rect 11152 6808 11204 6860
rect 11704 6808 11756 6860
rect 13728 6876 13780 6928
rect 15476 6876 15528 6928
rect 15936 6876 15988 6928
rect 17592 6876 17644 6928
rect 19524 6876 19576 6928
rect 12624 6808 12676 6860
rect 16948 6808 17000 6860
rect 17040 6808 17092 6860
rect 22100 6808 22152 6860
rect 9680 6740 9732 6792
rect 8852 6672 8904 6724
rect 9312 6672 9364 6724
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 10416 6783 10468 6792
rect 10416 6749 10425 6783
rect 10425 6749 10459 6783
rect 10459 6749 10468 6783
rect 10416 6740 10468 6749
rect 10968 6783 11020 6792
rect 10968 6749 10977 6783
rect 10977 6749 11011 6783
rect 11011 6749 11020 6783
rect 10968 6740 11020 6749
rect 11612 6740 11664 6792
rect 11796 6740 11848 6792
rect 10600 6672 10652 6724
rect 12808 6740 12860 6792
rect 14096 6740 14148 6792
rect 18236 6740 18288 6792
rect 12992 6672 13044 6724
rect 13360 6672 13412 6724
rect 14464 6715 14516 6724
rect 14464 6681 14473 6715
rect 14473 6681 14507 6715
rect 14507 6681 14516 6715
rect 14464 6672 14516 6681
rect 15200 6672 15252 6724
rect 16764 6672 16816 6724
rect 18880 6740 18932 6792
rect 19340 6740 19392 6792
rect 19984 6740 20036 6792
rect 22284 6808 22336 6860
rect 23020 6808 23072 6860
rect 23756 6851 23808 6860
rect 23756 6817 23765 6851
rect 23765 6817 23799 6851
rect 23799 6817 23808 6851
rect 23756 6808 23808 6817
rect 6644 6604 6696 6656
rect 8116 6604 8168 6656
rect 8760 6604 8812 6656
rect 17224 6604 17276 6656
rect 19892 6672 19944 6724
rect 21364 6672 21416 6724
rect 18420 6647 18472 6656
rect 18420 6613 18437 6647
rect 18437 6613 18472 6647
rect 18420 6604 18472 6613
rect 18972 6647 19024 6656
rect 18972 6613 18981 6647
rect 18981 6613 19015 6647
rect 19015 6613 19024 6647
rect 18972 6604 19024 6613
rect 20076 6604 20128 6656
rect 22008 6604 22060 6656
rect 23020 6604 23072 6656
rect 23112 6647 23164 6656
rect 23112 6613 23121 6647
rect 23121 6613 23155 6647
rect 23155 6613 23164 6647
rect 23112 6604 23164 6613
rect 23296 6604 23348 6656
rect 8214 6502 8266 6554
rect 8278 6502 8330 6554
rect 8342 6502 8394 6554
rect 8406 6502 8458 6554
rect 8470 6502 8522 6554
rect 16214 6502 16266 6554
rect 16278 6502 16330 6554
rect 16342 6502 16394 6554
rect 16406 6502 16458 6554
rect 16470 6502 16522 6554
rect 24214 6502 24266 6554
rect 24278 6502 24330 6554
rect 24342 6502 24394 6554
rect 24406 6502 24458 6554
rect 24470 6502 24522 6554
rect 2320 6307 2372 6316
rect 2320 6273 2329 6307
rect 2329 6273 2363 6307
rect 2363 6273 2372 6307
rect 2320 6264 2372 6273
rect 2780 6332 2832 6384
rect 2412 6239 2464 6248
rect 2412 6205 2421 6239
rect 2421 6205 2455 6239
rect 2455 6205 2464 6239
rect 2412 6196 2464 6205
rect 3516 6264 3568 6316
rect 6644 6400 6696 6452
rect 7564 6400 7616 6452
rect 6736 6332 6788 6384
rect 8116 6400 8168 6452
rect 8576 6400 8628 6452
rect 8944 6443 8996 6452
rect 8944 6409 8953 6443
rect 8953 6409 8987 6443
rect 8987 6409 8996 6443
rect 8944 6400 8996 6409
rect 9404 6400 9456 6452
rect 10232 6400 10284 6452
rect 3148 6196 3200 6248
rect 4988 6307 5040 6316
rect 4988 6273 4997 6307
rect 4997 6273 5031 6307
rect 5031 6273 5040 6307
rect 4988 6264 5040 6273
rect 5356 6264 5408 6316
rect 6000 6264 6052 6316
rect 6552 6307 6604 6316
rect 6552 6273 6562 6307
rect 6562 6273 6596 6307
rect 6596 6273 6604 6307
rect 6552 6264 6604 6273
rect 7012 6264 7064 6316
rect 7196 6264 7248 6316
rect 7840 6375 7892 6384
rect 7840 6341 7849 6375
rect 7849 6341 7883 6375
rect 7883 6341 7892 6375
rect 7840 6332 7892 6341
rect 9220 6332 9272 6384
rect 14096 6400 14148 6452
rect 14464 6400 14516 6452
rect 15568 6400 15620 6452
rect 16764 6443 16816 6452
rect 16764 6409 16773 6443
rect 16773 6409 16807 6443
rect 16807 6409 16816 6443
rect 16764 6400 16816 6409
rect 17224 6443 17276 6452
rect 17224 6409 17233 6443
rect 17233 6409 17267 6443
rect 17267 6409 17276 6443
rect 17224 6400 17276 6409
rect 17868 6443 17920 6452
rect 17868 6409 17877 6443
rect 17877 6409 17911 6443
rect 17911 6409 17920 6443
rect 17868 6400 17920 6409
rect 20720 6400 20772 6452
rect 9404 6307 9456 6316
rect 9404 6273 9413 6307
rect 9413 6273 9447 6307
rect 9447 6273 9456 6307
rect 9404 6264 9456 6273
rect 9680 6264 9732 6316
rect 10600 6307 10652 6316
rect 10600 6273 10609 6307
rect 10609 6273 10643 6307
rect 10643 6273 10652 6307
rect 10600 6264 10652 6273
rect 10968 6307 11020 6316
rect 10968 6273 10977 6307
rect 10977 6273 11011 6307
rect 11011 6273 11020 6307
rect 10968 6264 11020 6273
rect 13360 6264 13412 6316
rect 5632 6196 5684 6248
rect 5908 6196 5960 6248
rect 5172 6128 5224 6180
rect 5448 6171 5500 6180
rect 5448 6137 5457 6171
rect 5457 6137 5491 6171
rect 5491 6137 5500 6171
rect 5448 6128 5500 6137
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 3056 6103 3108 6112
rect 3056 6069 3065 6103
rect 3065 6069 3099 6103
rect 3099 6069 3108 6103
rect 3056 6060 3108 6069
rect 6092 6103 6144 6112
rect 6092 6069 6101 6103
rect 6101 6069 6135 6103
rect 6135 6069 6144 6103
rect 6092 6060 6144 6069
rect 7564 6103 7616 6112
rect 7564 6069 7573 6103
rect 7573 6069 7607 6103
rect 7607 6069 7616 6103
rect 7564 6060 7616 6069
rect 8576 6060 8628 6112
rect 9036 6060 9088 6112
rect 12072 6239 12124 6248
rect 12072 6205 12081 6239
rect 12081 6205 12115 6239
rect 12115 6205 12124 6239
rect 12072 6196 12124 6205
rect 14372 6264 14424 6316
rect 15108 6307 15160 6316
rect 15108 6273 15117 6307
rect 15117 6273 15151 6307
rect 15151 6273 15160 6307
rect 15108 6264 15160 6273
rect 13912 6196 13964 6248
rect 15844 6307 15896 6316
rect 15844 6273 15853 6307
rect 15853 6273 15887 6307
rect 15887 6273 15896 6307
rect 15844 6264 15896 6273
rect 16948 6264 17000 6316
rect 18052 6332 18104 6384
rect 22100 6400 22152 6452
rect 21088 6332 21140 6384
rect 21548 6332 21600 6384
rect 23112 6400 23164 6452
rect 24032 6443 24084 6452
rect 24032 6409 24041 6443
rect 24041 6409 24075 6443
rect 24075 6409 24084 6443
rect 24032 6400 24084 6409
rect 23940 6332 23992 6384
rect 17960 6307 18012 6316
rect 17960 6273 17969 6307
rect 17969 6273 18003 6307
rect 18003 6273 18012 6307
rect 17960 6264 18012 6273
rect 17500 6196 17552 6248
rect 17776 6196 17828 6248
rect 18512 6307 18564 6316
rect 18512 6273 18521 6307
rect 18521 6273 18555 6307
rect 18555 6273 18564 6307
rect 18512 6264 18564 6273
rect 19708 6264 19760 6316
rect 20812 6264 20864 6316
rect 19064 6239 19116 6248
rect 19064 6205 19073 6239
rect 19073 6205 19107 6239
rect 19107 6205 19116 6239
rect 19064 6196 19116 6205
rect 19340 6196 19392 6248
rect 19800 6196 19852 6248
rect 22376 6196 22428 6248
rect 22652 6196 22704 6248
rect 24676 6332 24728 6384
rect 14004 6128 14056 6180
rect 16856 6128 16908 6180
rect 18972 6128 19024 6180
rect 13360 6060 13412 6112
rect 14280 6103 14332 6112
rect 14280 6069 14289 6103
rect 14289 6069 14323 6103
rect 14323 6069 14332 6103
rect 14280 6060 14332 6069
rect 16672 6060 16724 6112
rect 16948 6060 17000 6112
rect 19340 6060 19392 6112
rect 19524 6103 19576 6112
rect 19524 6069 19533 6103
rect 19533 6069 19567 6103
rect 19567 6069 19576 6103
rect 19524 6060 19576 6069
rect 21180 6060 21232 6112
rect 21640 6060 21692 6112
rect 23388 6128 23440 6180
rect 22284 6060 22336 6112
rect 23296 6060 23348 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 12214 5958 12266 6010
rect 12278 5958 12330 6010
rect 12342 5958 12394 6010
rect 12406 5958 12458 6010
rect 12470 5958 12522 6010
rect 20214 5958 20266 6010
rect 20278 5958 20330 6010
rect 20342 5958 20394 6010
rect 20406 5958 20458 6010
rect 20470 5958 20522 6010
rect 2320 5856 2372 5908
rect 4988 5856 5040 5908
rect 5448 5856 5500 5908
rect 3976 5788 4028 5840
rect 2228 5763 2280 5772
rect 2228 5729 2237 5763
rect 2237 5729 2271 5763
rect 2271 5729 2280 5763
rect 2228 5720 2280 5729
rect 1768 5695 1820 5704
rect 1768 5661 1777 5695
rect 1777 5661 1811 5695
rect 1811 5661 1820 5695
rect 1768 5652 1820 5661
rect 2044 5652 2096 5704
rect 3056 5652 3108 5704
rect 2412 5584 2464 5636
rect 5540 5788 5592 5840
rect 3792 5652 3844 5704
rect 4068 5652 4120 5704
rect 5172 5652 5224 5704
rect 5540 5695 5592 5704
rect 5540 5661 5550 5695
rect 5550 5661 5584 5695
rect 5584 5661 5592 5695
rect 5540 5652 5592 5661
rect 5724 5695 5776 5704
rect 5724 5661 5733 5695
rect 5733 5661 5767 5695
rect 5767 5661 5776 5695
rect 5724 5652 5776 5661
rect 5908 5695 5960 5704
rect 7840 5856 7892 5908
rect 5908 5661 5922 5695
rect 5922 5661 5956 5695
rect 5956 5661 5960 5695
rect 5908 5652 5960 5661
rect 6736 5652 6788 5704
rect 6460 5627 6512 5636
rect 6460 5593 6469 5627
rect 6469 5593 6503 5627
rect 6503 5593 6512 5627
rect 8116 5652 8168 5704
rect 9312 5856 9364 5908
rect 12072 5856 12124 5908
rect 17132 5856 17184 5908
rect 17684 5856 17736 5908
rect 19616 5856 19668 5908
rect 20076 5856 20128 5908
rect 8576 5788 8628 5840
rect 8852 5788 8904 5840
rect 11704 5788 11756 5840
rect 11980 5788 12032 5840
rect 8944 5652 8996 5704
rect 10324 5720 10376 5772
rect 11888 5720 11940 5772
rect 15660 5788 15712 5840
rect 17408 5788 17460 5840
rect 18328 5788 18380 5840
rect 20628 5856 20680 5908
rect 20996 5856 21048 5908
rect 6460 5584 6512 5593
rect 7840 5584 7892 5636
rect 9496 5695 9548 5704
rect 9496 5661 9505 5695
rect 9505 5661 9539 5695
rect 9539 5661 9548 5695
rect 9496 5652 9548 5661
rect 10232 5652 10284 5704
rect 10600 5584 10652 5636
rect 10876 5695 10928 5704
rect 10876 5661 10885 5695
rect 10885 5661 10919 5695
rect 10919 5661 10928 5695
rect 10876 5652 10928 5661
rect 11612 5695 11664 5704
rect 11612 5661 11620 5695
rect 11620 5661 11654 5695
rect 11654 5661 11664 5695
rect 11612 5652 11664 5661
rect 11980 5652 12032 5704
rect 12624 5652 12676 5704
rect 12716 5584 12768 5636
rect 12992 5584 13044 5636
rect 13360 5695 13412 5704
rect 13360 5661 13369 5695
rect 13369 5661 13403 5695
rect 13403 5661 13412 5695
rect 13360 5652 13412 5661
rect 13728 5652 13780 5704
rect 14280 5652 14332 5704
rect 15752 5763 15804 5772
rect 15752 5729 15761 5763
rect 15761 5729 15795 5763
rect 15795 5729 15804 5763
rect 15752 5720 15804 5729
rect 17316 5720 17368 5772
rect 20076 5720 20128 5772
rect 16580 5652 16632 5704
rect 18236 5695 18288 5704
rect 18236 5661 18245 5695
rect 18245 5661 18279 5695
rect 18279 5661 18288 5695
rect 18236 5652 18288 5661
rect 19248 5652 19300 5704
rect 19800 5652 19852 5704
rect 21272 5720 21324 5772
rect 22008 5788 22060 5840
rect 21916 5720 21968 5772
rect 22376 5763 22428 5772
rect 22376 5729 22385 5763
rect 22385 5729 22419 5763
rect 22419 5729 22428 5763
rect 22376 5720 22428 5729
rect 23020 5720 23072 5772
rect 22284 5652 22336 5704
rect 4620 5516 4672 5568
rect 7380 5516 7432 5568
rect 9588 5516 9640 5568
rect 10784 5516 10836 5568
rect 10968 5516 11020 5568
rect 11704 5516 11756 5568
rect 12808 5516 12860 5568
rect 13176 5516 13228 5568
rect 16672 5627 16724 5636
rect 16672 5593 16681 5627
rect 16681 5593 16715 5627
rect 16715 5593 16724 5627
rect 16672 5584 16724 5593
rect 16948 5584 17000 5636
rect 17408 5584 17460 5636
rect 14832 5559 14884 5568
rect 14832 5525 14841 5559
rect 14841 5525 14875 5559
rect 14875 5525 14884 5559
rect 14832 5516 14884 5525
rect 17040 5559 17092 5568
rect 17040 5525 17049 5559
rect 17049 5525 17083 5559
rect 17083 5525 17092 5559
rect 17040 5516 17092 5525
rect 17224 5516 17276 5568
rect 17960 5559 18012 5568
rect 17960 5525 17969 5559
rect 17969 5525 18003 5559
rect 18003 5525 18012 5559
rect 17960 5516 18012 5525
rect 19156 5516 19208 5568
rect 20904 5584 20956 5636
rect 22652 5627 22704 5636
rect 22652 5593 22661 5627
rect 22661 5593 22695 5627
rect 22695 5593 22704 5627
rect 22652 5584 22704 5593
rect 23664 5584 23716 5636
rect 21088 5516 21140 5568
rect 21364 5516 21416 5568
rect 24676 5516 24728 5568
rect 8214 5414 8266 5466
rect 8278 5414 8330 5466
rect 8342 5414 8394 5466
rect 8406 5414 8458 5466
rect 8470 5414 8522 5466
rect 16214 5414 16266 5466
rect 16278 5414 16330 5466
rect 16342 5414 16394 5466
rect 16406 5414 16458 5466
rect 16470 5414 16522 5466
rect 24214 5414 24266 5466
rect 24278 5414 24330 5466
rect 24342 5414 24394 5466
rect 24406 5414 24458 5466
rect 24470 5414 24522 5466
rect 2228 5312 2280 5364
rect 1676 5287 1728 5296
rect 1676 5253 1685 5287
rect 1685 5253 1719 5287
rect 1719 5253 1728 5287
rect 1676 5244 1728 5253
rect 7288 5355 7340 5364
rect 7288 5321 7297 5355
rect 7297 5321 7331 5355
rect 7331 5321 7340 5355
rect 7288 5312 7340 5321
rect 7380 5355 7432 5364
rect 7380 5321 7389 5355
rect 7389 5321 7423 5355
rect 7423 5321 7432 5355
rect 7380 5312 7432 5321
rect 7932 5312 7984 5364
rect 2412 5176 2464 5228
rect 3056 5219 3108 5228
rect 3056 5185 3065 5219
rect 3065 5185 3099 5219
rect 3099 5185 3108 5219
rect 3056 5176 3108 5185
rect 3976 5176 4028 5228
rect 4896 5176 4948 5228
rect 4620 5108 4672 5160
rect 4804 5151 4856 5160
rect 4804 5117 4813 5151
rect 4813 5117 4847 5151
rect 4847 5117 4856 5151
rect 4804 5108 4856 5117
rect 5540 5244 5592 5296
rect 6460 5244 6512 5296
rect 10324 5312 10376 5364
rect 9496 5244 9548 5296
rect 6276 5176 6328 5228
rect 7012 5219 7064 5228
rect 7012 5185 7021 5219
rect 7021 5185 7055 5219
rect 7055 5185 7064 5219
rect 7012 5176 7064 5185
rect 7564 5176 7616 5228
rect 7840 5219 7892 5228
rect 7840 5185 7849 5219
rect 7849 5185 7883 5219
rect 7883 5185 7892 5219
rect 7840 5176 7892 5185
rect 6184 5108 6236 5160
rect 2044 5083 2096 5092
rect 2044 5049 2053 5083
rect 2053 5049 2087 5083
rect 2087 5049 2096 5083
rect 2044 5040 2096 5049
rect 2320 5040 2372 5092
rect 8116 5108 8168 5160
rect 8668 5219 8720 5228
rect 8668 5185 8677 5219
rect 8677 5185 8711 5219
rect 8711 5185 8720 5219
rect 8668 5176 8720 5185
rect 10232 5219 10284 5228
rect 10232 5185 10241 5219
rect 10241 5185 10275 5219
rect 10275 5185 10284 5219
rect 10232 5176 10284 5185
rect 10416 5219 10468 5228
rect 10416 5185 10425 5219
rect 10425 5185 10459 5219
rect 10459 5185 10468 5219
rect 10416 5176 10468 5185
rect 10692 5219 10744 5228
rect 10692 5185 10701 5219
rect 10701 5185 10735 5219
rect 10735 5185 10744 5219
rect 10692 5176 10744 5185
rect 12624 5312 12676 5364
rect 12716 5312 12768 5364
rect 15108 5312 15160 5364
rect 15568 5312 15620 5364
rect 11612 5244 11664 5296
rect 11980 5219 12032 5228
rect 11980 5185 11988 5219
rect 11988 5185 12022 5219
rect 12022 5185 12032 5219
rect 11980 5176 12032 5185
rect 9128 5108 9180 5160
rect 9680 5151 9732 5160
rect 9680 5117 9689 5151
rect 9689 5117 9723 5151
rect 9723 5117 9732 5151
rect 9680 5108 9732 5117
rect 13544 5219 13596 5228
rect 13544 5185 13553 5219
rect 13553 5185 13587 5219
rect 13587 5185 13596 5219
rect 13544 5176 13596 5185
rect 3332 4972 3384 5024
rect 3516 5015 3568 5024
rect 3516 4981 3525 5015
rect 3525 4981 3559 5015
rect 3559 4981 3568 5015
rect 3516 4972 3568 4981
rect 5264 4972 5316 5024
rect 6460 5015 6512 5024
rect 6460 4981 6469 5015
rect 6469 4981 6503 5015
rect 6503 4981 6512 5015
rect 6460 4972 6512 4981
rect 7012 4972 7064 5024
rect 7380 4972 7432 5024
rect 11888 5040 11940 5092
rect 12716 5151 12768 5160
rect 12716 5117 12725 5151
rect 12725 5117 12759 5151
rect 12759 5117 12768 5151
rect 12716 5108 12768 5117
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 13452 5108 13504 5160
rect 13820 5219 13872 5228
rect 13820 5185 13829 5219
rect 13829 5185 13863 5219
rect 13863 5185 13872 5219
rect 13820 5176 13872 5185
rect 14372 5244 14424 5296
rect 14832 5287 14884 5296
rect 14832 5253 14841 5287
rect 14841 5253 14875 5287
rect 14875 5253 14884 5287
rect 14832 5244 14884 5253
rect 13912 5040 13964 5092
rect 15016 5176 15068 5228
rect 17960 5244 18012 5296
rect 18696 5355 18748 5364
rect 18696 5321 18705 5355
rect 18705 5321 18739 5355
rect 18739 5321 18748 5355
rect 18696 5312 18748 5321
rect 19064 5312 19116 5364
rect 19524 5244 19576 5296
rect 19708 5244 19760 5296
rect 16856 5176 16908 5228
rect 14740 5108 14792 5160
rect 15752 5108 15804 5160
rect 16120 5151 16172 5160
rect 16120 5117 16129 5151
rect 16129 5117 16163 5151
rect 16163 5117 16172 5151
rect 16120 5108 16172 5117
rect 16764 5108 16816 5160
rect 15384 5040 15436 5092
rect 11980 4972 12032 5024
rect 12808 4972 12860 5024
rect 16580 5040 16632 5092
rect 16672 4972 16724 5024
rect 17316 5108 17368 5160
rect 19984 5108 20036 5160
rect 20720 5355 20772 5364
rect 20720 5321 20729 5355
rect 20729 5321 20763 5355
rect 20763 5321 20772 5355
rect 20720 5312 20772 5321
rect 20904 5312 20956 5364
rect 21548 5312 21600 5364
rect 21364 5287 21416 5296
rect 21364 5253 21373 5287
rect 21373 5253 21407 5287
rect 21407 5253 21416 5287
rect 22652 5312 22704 5364
rect 23020 5312 23072 5364
rect 23296 5355 23348 5364
rect 23296 5321 23305 5355
rect 23305 5321 23339 5355
rect 23339 5321 23348 5355
rect 23296 5312 23348 5321
rect 23940 5312 23992 5364
rect 21364 5244 21416 5253
rect 20996 5176 21048 5228
rect 21732 5176 21784 5228
rect 21364 5108 21416 5160
rect 23388 5151 23440 5160
rect 23388 5117 23397 5151
rect 23397 5117 23431 5151
rect 23431 5117 23440 5151
rect 23388 5108 23440 5117
rect 20720 4972 20772 5024
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 22744 4972 22796 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 12214 4870 12266 4922
rect 12278 4870 12330 4922
rect 12342 4870 12394 4922
rect 12406 4870 12458 4922
rect 12470 4870 12522 4922
rect 20214 4870 20266 4922
rect 20278 4870 20330 4922
rect 20342 4870 20394 4922
rect 20406 4870 20458 4922
rect 20470 4870 20522 4922
rect 1400 4768 1452 4820
rect 2044 4768 2096 4820
rect 2688 4768 2740 4820
rect 1860 4743 1912 4752
rect 1860 4709 1869 4743
rect 1869 4709 1903 4743
rect 1903 4709 1912 4743
rect 1860 4700 1912 4709
rect 2780 4700 2832 4752
rect 4896 4768 4948 4820
rect 7288 4768 7340 4820
rect 8760 4768 8812 4820
rect 2964 4675 3016 4684
rect 2964 4641 2973 4675
rect 2973 4641 3007 4675
rect 3007 4641 3016 4675
rect 2964 4632 3016 4641
rect 4068 4632 4120 4684
rect 5540 4632 5592 4684
rect 6184 4675 6236 4684
rect 6184 4641 6193 4675
rect 6193 4641 6227 4675
rect 6227 4641 6236 4675
rect 6184 4632 6236 4641
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 7196 4632 7248 4684
rect 7380 4675 7432 4684
rect 7380 4641 7389 4675
rect 7389 4641 7423 4675
rect 7423 4641 7432 4675
rect 7380 4632 7432 4641
rect 9128 4632 9180 4684
rect 2320 4607 2372 4616
rect 2320 4573 2329 4607
rect 2329 4573 2363 4607
rect 2363 4573 2372 4607
rect 2320 4564 2372 4573
rect 2228 4471 2280 4480
rect 2228 4437 2237 4471
rect 2237 4437 2271 4471
rect 2271 4437 2280 4471
rect 2228 4428 2280 4437
rect 2504 4428 2556 4480
rect 3240 4564 3292 4616
rect 3516 4564 3568 4616
rect 3976 4564 4028 4616
rect 4620 4607 4672 4616
rect 4620 4573 4629 4607
rect 4629 4573 4663 4607
rect 4663 4573 4672 4607
rect 4620 4564 4672 4573
rect 4804 4564 4856 4616
rect 5448 4607 5500 4616
rect 5448 4573 5457 4607
rect 5457 4573 5491 4607
rect 5491 4573 5500 4607
rect 5448 4564 5500 4573
rect 7012 4607 7064 4616
rect 7012 4573 7021 4607
rect 7021 4573 7055 4607
rect 7055 4573 7064 4607
rect 7012 4564 7064 4573
rect 7104 4564 7156 4616
rect 7656 4564 7708 4616
rect 8668 4607 8720 4616
rect 8668 4573 8677 4607
rect 8677 4573 8711 4607
rect 8711 4573 8720 4607
rect 8668 4564 8720 4573
rect 10876 4768 10928 4820
rect 12716 4768 12768 4820
rect 13820 4768 13872 4820
rect 17316 4811 17368 4820
rect 17316 4777 17325 4811
rect 17325 4777 17359 4811
rect 17359 4777 17368 4811
rect 17316 4768 17368 4777
rect 9680 4564 9732 4616
rect 11704 4700 11756 4752
rect 12624 4743 12676 4752
rect 12624 4709 12633 4743
rect 12633 4709 12667 4743
rect 12667 4709 12676 4743
rect 12624 4700 12676 4709
rect 14280 4700 14332 4752
rect 15016 4700 15068 4752
rect 15108 4700 15160 4752
rect 10324 4564 10376 4616
rect 10692 4564 10744 4616
rect 9956 4496 10008 4548
rect 10048 4496 10100 4548
rect 2872 4428 2924 4480
rect 5356 4428 5408 4480
rect 6828 4428 6880 4480
rect 10416 4428 10468 4480
rect 10692 4428 10744 4480
rect 10968 4607 11020 4616
rect 10968 4573 10977 4607
rect 10977 4573 11011 4607
rect 11011 4573 11020 4607
rect 10968 4564 11020 4573
rect 11428 4607 11480 4616
rect 11428 4573 11437 4607
rect 11437 4573 11471 4607
rect 11471 4573 11480 4607
rect 11428 4564 11480 4573
rect 11980 4632 12032 4684
rect 11704 4607 11756 4616
rect 11704 4573 11713 4607
rect 11713 4573 11747 4607
rect 11747 4573 11756 4607
rect 11704 4564 11756 4573
rect 10876 4539 10928 4548
rect 10876 4505 10885 4539
rect 10885 4505 10919 4539
rect 10919 4505 10928 4539
rect 10876 4496 10928 4505
rect 11888 4496 11940 4548
rect 12808 4564 12860 4616
rect 14464 4632 14516 4684
rect 12900 4496 12952 4548
rect 13360 4607 13412 4616
rect 13360 4573 13369 4607
rect 13369 4573 13403 4607
rect 13403 4573 13412 4607
rect 13360 4564 13412 4573
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 13544 4607 13596 4616
rect 13544 4573 13589 4607
rect 13589 4573 13596 4607
rect 13544 4564 13596 4573
rect 13728 4607 13780 4616
rect 13728 4573 13737 4607
rect 13737 4573 13771 4607
rect 13771 4573 13780 4607
rect 13728 4564 13780 4573
rect 14280 4564 14332 4616
rect 14372 4607 14424 4616
rect 14372 4573 14381 4607
rect 14381 4573 14415 4607
rect 14415 4573 14424 4607
rect 14372 4564 14424 4573
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 14832 4564 14884 4616
rect 14924 4607 14976 4616
rect 14924 4573 14933 4607
rect 14933 4573 14967 4607
rect 14967 4573 14976 4607
rect 14924 4564 14976 4573
rect 15016 4564 15068 4616
rect 15660 4632 15712 4684
rect 19708 4811 19760 4820
rect 19708 4777 19717 4811
rect 19717 4777 19751 4811
rect 19751 4777 19760 4811
rect 19708 4768 19760 4777
rect 20720 4768 20772 4820
rect 22376 4811 22428 4820
rect 22376 4777 22385 4811
rect 22385 4777 22419 4811
rect 22419 4777 22428 4811
rect 22376 4768 22428 4777
rect 23020 4768 23072 4820
rect 23756 4768 23808 4820
rect 24124 4811 24176 4820
rect 24124 4777 24133 4811
rect 24133 4777 24167 4811
rect 24167 4777 24176 4811
rect 24124 4768 24176 4777
rect 17500 4632 17552 4684
rect 19616 4632 19668 4684
rect 11244 4471 11296 4480
rect 11244 4437 11253 4471
rect 11253 4437 11287 4471
rect 11287 4437 11296 4471
rect 11244 4428 11296 4437
rect 11704 4428 11756 4480
rect 13820 4428 13872 4480
rect 15384 4496 15436 4548
rect 18696 4564 18748 4616
rect 18880 4607 18932 4616
rect 18880 4573 18889 4607
rect 18889 4573 18923 4607
rect 18923 4573 18932 4607
rect 18880 4564 18932 4573
rect 19800 4564 19852 4616
rect 19340 4539 19392 4548
rect 19340 4505 19349 4539
rect 19349 4505 19383 4539
rect 19383 4505 19392 4539
rect 19340 4496 19392 4505
rect 19616 4496 19668 4548
rect 21548 4632 21600 4684
rect 23204 4675 23256 4684
rect 23204 4641 23213 4675
rect 23213 4641 23247 4675
rect 23247 4641 23256 4675
rect 23204 4632 23256 4641
rect 19984 4607 20036 4616
rect 19984 4573 19993 4607
rect 19993 4573 20027 4607
rect 20027 4573 20036 4607
rect 19984 4564 20036 4573
rect 15844 4428 15896 4480
rect 17592 4428 17644 4480
rect 20720 4496 20772 4548
rect 22100 4539 22152 4548
rect 22100 4505 22109 4539
rect 22109 4505 22143 4539
rect 22143 4505 22152 4539
rect 22100 4496 22152 4505
rect 20076 4428 20128 4480
rect 21732 4471 21784 4480
rect 21732 4437 21741 4471
rect 21741 4437 21775 4471
rect 21775 4437 21784 4471
rect 21732 4428 21784 4437
rect 23296 4471 23348 4480
rect 23296 4437 23305 4471
rect 23305 4437 23339 4471
rect 23339 4437 23348 4471
rect 23296 4428 23348 4437
rect 23388 4471 23440 4480
rect 23388 4437 23397 4471
rect 23397 4437 23431 4471
rect 23431 4437 23440 4471
rect 23388 4428 23440 4437
rect 23940 4428 23992 4480
rect 8214 4326 8266 4378
rect 8278 4326 8330 4378
rect 8342 4326 8394 4378
rect 8406 4326 8458 4378
rect 8470 4326 8522 4378
rect 16214 4326 16266 4378
rect 16278 4326 16330 4378
rect 16342 4326 16394 4378
rect 16406 4326 16458 4378
rect 16470 4326 16522 4378
rect 24214 4326 24266 4378
rect 24278 4326 24330 4378
rect 24342 4326 24394 4378
rect 24406 4326 24458 4378
rect 24470 4326 24522 4378
rect 2780 4224 2832 4276
rect 4620 4224 4672 4276
rect 2044 4156 2096 4208
rect 2412 4156 2464 4208
rect 7104 4224 7156 4276
rect 9680 4224 9732 4276
rect 10600 4224 10652 4276
rect 11244 4224 11296 4276
rect 13728 4224 13780 4276
rect 3976 4131 4028 4140
rect 3976 4097 3985 4131
rect 3985 4097 4019 4131
rect 4019 4097 4028 4131
rect 3976 4088 4028 4097
rect 4068 4088 4120 4140
rect 4896 4088 4948 4140
rect 5264 4131 5316 4140
rect 5264 4097 5273 4131
rect 5273 4097 5307 4131
rect 5307 4097 5316 4131
rect 5264 4088 5316 4097
rect 5356 4131 5408 4140
rect 5356 4097 5365 4131
rect 5365 4097 5399 4131
rect 5399 4097 5408 4131
rect 5356 4088 5408 4097
rect 1492 4020 1544 4072
rect 3148 4020 3200 4072
rect 4712 4020 4764 4072
rect 6828 4156 6880 4208
rect 7380 4156 7432 4208
rect 9588 4156 9640 4208
rect 9312 4088 9364 4140
rect 9772 4088 9824 4140
rect 6000 4020 6052 4072
rect 3332 3952 3384 4004
rect 3240 3884 3292 3936
rect 4896 3884 4948 3936
rect 5172 3884 5224 3936
rect 6552 3884 6604 3936
rect 7012 4020 7064 4072
rect 7472 4020 7524 4072
rect 7656 4020 7708 4072
rect 9680 4020 9732 4072
rect 9956 4131 10008 4140
rect 9956 4097 9965 4131
rect 9965 4097 9999 4131
rect 9999 4097 10008 4131
rect 9956 4088 10008 4097
rect 10324 4156 10376 4208
rect 10600 4088 10652 4140
rect 10692 4131 10744 4140
rect 10692 4097 10701 4131
rect 10701 4097 10735 4131
rect 10735 4097 10744 4131
rect 10692 4088 10744 4097
rect 10876 4156 10928 4208
rect 13912 4224 13964 4276
rect 14924 4224 14976 4276
rect 10784 4020 10836 4072
rect 11980 4088 12032 4140
rect 12716 4088 12768 4140
rect 11888 4020 11940 4072
rect 12072 4063 12124 4072
rect 12072 4029 12081 4063
rect 12081 4029 12115 4063
rect 12115 4029 12124 4063
rect 12072 4020 12124 4029
rect 7104 3884 7156 3936
rect 7472 3884 7524 3936
rect 8760 3952 8812 4004
rect 12808 4020 12860 4072
rect 12716 3952 12768 4004
rect 13544 4088 13596 4140
rect 15016 4088 15068 4140
rect 15936 4224 15988 4276
rect 16120 4267 16172 4276
rect 16120 4233 16129 4267
rect 16129 4233 16163 4267
rect 16163 4233 16172 4267
rect 16120 4224 16172 4233
rect 17684 4224 17736 4276
rect 15568 4156 15620 4208
rect 15660 4131 15712 4140
rect 15660 4097 15669 4131
rect 15669 4097 15703 4131
rect 15703 4097 15712 4131
rect 15660 4088 15712 4097
rect 17040 4156 17092 4208
rect 15476 4020 15528 4072
rect 15568 4063 15620 4072
rect 15568 4029 15577 4063
rect 15577 4029 15611 4063
rect 15611 4029 15620 4063
rect 15568 4020 15620 4029
rect 13636 3952 13688 4004
rect 8668 3884 8720 3936
rect 9680 3927 9732 3936
rect 9680 3893 9689 3927
rect 9689 3893 9723 3927
rect 9723 3893 9732 3927
rect 9680 3884 9732 3893
rect 11888 3884 11940 3936
rect 13452 3884 13504 3936
rect 15200 3952 15252 4004
rect 14188 3884 14240 3936
rect 15752 3884 15804 3936
rect 16120 3884 16172 3936
rect 16764 4063 16816 4072
rect 16764 4029 16773 4063
rect 16773 4029 16807 4063
rect 16807 4029 16816 4063
rect 16764 4020 16816 4029
rect 17040 4063 17092 4072
rect 17040 4029 17049 4063
rect 17049 4029 17083 4063
rect 17083 4029 17092 4063
rect 17040 4020 17092 4029
rect 18880 4156 18932 4208
rect 18880 4020 18932 4072
rect 19616 4224 19668 4276
rect 20076 4224 20128 4276
rect 20996 4224 21048 4276
rect 21548 4267 21600 4276
rect 21548 4233 21557 4267
rect 21557 4233 21591 4267
rect 21591 4233 21600 4267
rect 21548 4224 21600 4233
rect 19340 4156 19392 4208
rect 21732 4156 21784 4208
rect 20812 4088 20864 4140
rect 21088 4088 21140 4140
rect 23480 4224 23532 4276
rect 24124 4156 24176 4208
rect 24584 4088 24636 4140
rect 21180 4020 21232 4072
rect 22008 4020 22060 4072
rect 18972 3952 19024 4004
rect 18236 3884 18288 3936
rect 19984 3952 20036 4004
rect 21916 3952 21968 4004
rect 22560 4020 22612 4072
rect 23204 4020 23256 4072
rect 19800 3884 19852 3936
rect 20720 3884 20772 3936
rect 23848 3952 23900 4004
rect 23756 3884 23808 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 12214 3782 12266 3834
rect 12278 3782 12330 3834
rect 12342 3782 12394 3834
rect 12406 3782 12458 3834
rect 12470 3782 12522 3834
rect 20214 3782 20266 3834
rect 20278 3782 20330 3834
rect 20342 3782 20394 3834
rect 20406 3782 20458 3834
rect 20470 3782 20522 3834
rect 2044 3680 2096 3732
rect 2412 3680 2464 3732
rect 2596 3655 2648 3664
rect 2596 3621 2605 3655
rect 2605 3621 2639 3655
rect 2639 3621 2648 3655
rect 2596 3612 2648 3621
rect 2320 3544 2372 3596
rect 3976 3612 4028 3664
rect 6368 3680 6420 3732
rect 7012 3680 7064 3732
rect 7380 3723 7432 3732
rect 7380 3689 7389 3723
rect 7389 3689 7423 3723
rect 7423 3689 7432 3723
rect 7380 3680 7432 3689
rect 9864 3680 9916 3732
rect 9956 3680 10008 3732
rect 10416 3680 10468 3732
rect 11612 3680 11664 3732
rect 12716 3680 12768 3732
rect 7656 3612 7708 3664
rect 1400 3476 1452 3528
rect 2228 3476 2280 3528
rect 2136 3383 2188 3392
rect 2136 3349 2161 3383
rect 2161 3349 2188 3383
rect 2412 3408 2464 3460
rect 3148 3587 3200 3596
rect 3148 3553 3157 3587
rect 3157 3553 3191 3587
rect 3191 3553 3200 3587
rect 3148 3544 3200 3553
rect 3240 3544 3292 3596
rect 7104 3544 7156 3596
rect 7196 3544 7248 3596
rect 3332 3476 3384 3528
rect 3056 3408 3108 3460
rect 4804 3408 4856 3460
rect 2136 3340 2188 3349
rect 3700 3340 3752 3392
rect 3792 3340 3844 3392
rect 4712 3340 4764 3392
rect 7288 3476 7340 3528
rect 7932 3519 7984 3528
rect 7932 3485 7941 3519
rect 7941 3485 7975 3519
rect 7975 3485 7984 3519
rect 7932 3476 7984 3485
rect 8116 3519 8168 3528
rect 8116 3485 8125 3519
rect 8125 3485 8159 3519
rect 8159 3485 8168 3519
rect 8116 3476 8168 3485
rect 10692 3612 10744 3664
rect 17040 3680 17092 3732
rect 18512 3680 18564 3732
rect 19892 3680 19944 3732
rect 21364 3680 21416 3732
rect 21916 3680 21968 3732
rect 22560 3723 22612 3732
rect 22560 3689 22569 3723
rect 22569 3689 22603 3723
rect 22603 3689 22612 3723
rect 22560 3680 22612 3689
rect 24032 3680 24084 3732
rect 9680 3544 9732 3596
rect 11060 3544 11112 3596
rect 5172 3451 5224 3460
rect 5172 3417 5181 3451
rect 5181 3417 5215 3451
rect 5215 3417 5224 3451
rect 5172 3408 5224 3417
rect 6184 3408 6236 3460
rect 6736 3408 6788 3460
rect 5540 3340 5592 3392
rect 6000 3340 6052 3392
rect 6920 3340 6972 3392
rect 7564 3408 7616 3460
rect 10876 3476 10928 3528
rect 13544 3587 13596 3596
rect 13544 3553 13553 3587
rect 13553 3553 13587 3587
rect 13587 3553 13596 3587
rect 13544 3544 13596 3553
rect 13636 3544 13688 3596
rect 13820 3587 13872 3596
rect 13820 3553 13829 3587
rect 13829 3553 13863 3587
rect 13863 3553 13872 3587
rect 13820 3544 13872 3553
rect 15844 3612 15896 3664
rect 19064 3612 19116 3664
rect 8024 3340 8076 3392
rect 9220 3408 9272 3460
rect 9404 3340 9456 3392
rect 11428 3451 11480 3460
rect 11428 3417 11437 3451
rect 11437 3417 11471 3451
rect 11471 3417 11480 3451
rect 11428 3408 11480 3417
rect 14096 3476 14148 3528
rect 14280 3519 14332 3528
rect 14280 3485 14289 3519
rect 14289 3485 14323 3519
rect 14323 3485 14332 3519
rect 14280 3476 14332 3485
rect 12900 3408 12952 3460
rect 14740 3519 14792 3528
rect 14740 3485 14749 3519
rect 14749 3485 14783 3519
rect 14783 3485 14792 3519
rect 14740 3476 14792 3485
rect 15292 3476 15344 3528
rect 15752 3476 15804 3528
rect 19984 3544 20036 3596
rect 16580 3476 16632 3528
rect 16948 3476 17000 3528
rect 17224 3476 17276 3528
rect 19248 3476 19300 3528
rect 19432 3476 19484 3528
rect 20076 3476 20128 3528
rect 20720 3612 20772 3664
rect 21548 3612 21600 3664
rect 23480 3612 23532 3664
rect 24124 3612 24176 3664
rect 21180 3587 21232 3596
rect 21180 3553 21189 3587
rect 21189 3553 21223 3587
rect 21223 3553 21232 3587
rect 21180 3544 21232 3553
rect 21364 3544 21416 3596
rect 21732 3544 21784 3596
rect 23112 3587 23164 3596
rect 23112 3553 23121 3587
rect 23121 3553 23155 3587
rect 23155 3553 23164 3587
rect 23112 3544 23164 3553
rect 22100 3476 22152 3528
rect 22192 3519 22244 3528
rect 22192 3485 22201 3519
rect 22201 3485 22235 3519
rect 22235 3485 22244 3519
rect 22192 3476 22244 3485
rect 23296 3476 23348 3528
rect 23572 3476 23624 3528
rect 24584 3476 24636 3528
rect 12072 3340 12124 3392
rect 15200 3383 15252 3392
rect 15200 3349 15209 3383
rect 15209 3349 15243 3383
rect 15243 3349 15252 3383
rect 15200 3340 15252 3349
rect 15384 3383 15436 3392
rect 15384 3349 15411 3383
rect 15411 3349 15436 3383
rect 15384 3340 15436 3349
rect 16028 3451 16080 3460
rect 16028 3417 16037 3451
rect 16037 3417 16071 3451
rect 16071 3417 16080 3451
rect 16028 3408 16080 3417
rect 16856 3383 16908 3392
rect 16856 3349 16865 3383
rect 16865 3349 16899 3383
rect 16899 3349 16908 3383
rect 16856 3340 16908 3349
rect 18236 3408 18288 3460
rect 18696 3451 18748 3460
rect 18696 3417 18705 3451
rect 18705 3417 18739 3451
rect 18739 3417 18748 3451
rect 18696 3408 18748 3417
rect 18788 3408 18840 3460
rect 18604 3340 18656 3392
rect 20628 3383 20680 3392
rect 20628 3349 20637 3383
rect 20637 3349 20671 3383
rect 20671 3349 20680 3383
rect 20628 3340 20680 3349
rect 20996 3383 21048 3392
rect 20996 3349 21005 3383
rect 21005 3349 21039 3383
rect 21039 3349 21048 3383
rect 20996 3340 21048 3349
rect 21088 3383 21140 3392
rect 21088 3349 21097 3383
rect 21097 3349 21131 3383
rect 21131 3349 21140 3383
rect 21088 3340 21140 3349
rect 21364 3408 21416 3460
rect 22376 3408 22428 3460
rect 24676 3408 24728 3460
rect 23572 3340 23624 3392
rect 24768 3340 24820 3392
rect 8214 3238 8266 3290
rect 8278 3238 8330 3290
rect 8342 3238 8394 3290
rect 8406 3238 8458 3290
rect 8470 3238 8522 3290
rect 16214 3238 16266 3290
rect 16278 3238 16330 3290
rect 16342 3238 16394 3290
rect 16406 3238 16458 3290
rect 16470 3238 16522 3290
rect 24214 3238 24266 3290
rect 24278 3238 24330 3290
rect 24342 3238 24394 3290
rect 24406 3238 24458 3290
rect 24470 3238 24522 3290
rect 2044 3136 2096 3188
rect 2228 3136 2280 3188
rect 5724 3136 5776 3188
rect 5816 3179 5868 3188
rect 5816 3145 5841 3179
rect 5841 3145 5868 3179
rect 5816 3136 5868 3145
rect 6184 3136 6236 3188
rect 6552 3136 6604 3188
rect 1584 3000 1636 3052
rect 2412 3068 2464 3120
rect 3056 3068 3108 3120
rect 3148 3000 3200 3052
rect 3516 3000 3568 3052
rect 3976 3000 4028 3052
rect 4804 3068 4856 3120
rect 2504 2932 2556 2984
rect 3332 2932 3384 2984
rect 4068 2864 4120 2916
rect 4620 2932 4672 2984
rect 4896 3000 4948 3052
rect 5448 3068 5500 3120
rect 6276 3068 6328 3120
rect 4804 2932 4856 2984
rect 6552 2975 6604 2984
rect 6552 2941 6561 2975
rect 6561 2941 6595 2975
rect 6595 2941 6604 2975
rect 6552 2932 6604 2941
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 7288 3043 7340 3052
rect 7288 3009 7297 3043
rect 7297 3009 7331 3043
rect 7331 3009 7340 3043
rect 7288 3000 7340 3009
rect 8024 3000 8076 3052
rect 10600 3136 10652 3188
rect 13360 3136 13412 3188
rect 16028 3179 16080 3188
rect 16028 3145 16037 3179
rect 16037 3145 16071 3179
rect 16071 3145 16080 3179
rect 16028 3136 16080 3145
rect 16856 3136 16908 3188
rect 17684 3136 17736 3188
rect 9680 3000 9732 3052
rect 10416 3043 10468 3052
rect 10416 3009 10425 3043
rect 10425 3009 10459 3043
rect 10459 3009 10468 3043
rect 10416 3000 10468 3009
rect 10876 3043 10928 3052
rect 10876 3009 10885 3043
rect 10885 3009 10919 3043
rect 10919 3009 10928 3043
rect 10876 3000 10928 3009
rect 11152 3000 11204 3052
rect 12716 3068 12768 3120
rect 13452 3068 13504 3120
rect 8576 2932 8628 2984
rect 5356 2907 5408 2916
rect 5356 2873 5365 2907
rect 5365 2873 5399 2907
rect 5399 2873 5408 2907
rect 5356 2864 5408 2873
rect 2320 2796 2372 2848
rect 2780 2839 2832 2848
rect 2780 2805 2789 2839
rect 2789 2805 2823 2839
rect 2823 2805 2832 2839
rect 2780 2796 2832 2805
rect 6368 2796 6420 2848
rect 7472 2907 7524 2916
rect 7472 2873 7481 2907
rect 7481 2873 7515 2907
rect 7515 2873 7524 2907
rect 7472 2864 7524 2873
rect 9588 2932 9640 2984
rect 10784 2975 10836 2984
rect 10784 2941 10793 2975
rect 10793 2941 10827 2975
rect 10827 2941 10836 2975
rect 10784 2932 10836 2941
rect 11888 2932 11940 2984
rect 12808 3043 12860 3052
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 17592 3111 17644 3120
rect 17592 3077 17601 3111
rect 17601 3077 17635 3111
rect 17635 3077 17644 3111
rect 17592 3068 17644 3077
rect 18696 3136 18748 3188
rect 18972 3136 19024 3188
rect 18512 3068 18564 3120
rect 18604 3111 18656 3120
rect 18604 3077 18613 3111
rect 18613 3077 18647 3111
rect 18647 3077 18656 3111
rect 18604 3068 18656 3077
rect 20996 3136 21048 3188
rect 14004 3043 14056 3052
rect 14004 3009 14013 3043
rect 14013 3009 14047 3043
rect 14047 3009 14056 3043
rect 14004 3000 14056 3009
rect 14188 3043 14240 3052
rect 14188 3009 14197 3043
rect 14197 3009 14231 3043
rect 14231 3009 14240 3043
rect 14188 3000 14240 3009
rect 12716 2932 12768 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 13268 2975 13320 2984
rect 13268 2941 13277 2975
rect 13277 2941 13311 2975
rect 13311 2941 13320 2975
rect 13268 2932 13320 2941
rect 15108 3000 15160 3052
rect 15200 3043 15252 3052
rect 15200 3009 15209 3043
rect 15209 3009 15243 3043
rect 15243 3009 15252 3043
rect 15200 3000 15252 3009
rect 15476 3000 15528 3052
rect 16856 3000 16908 3052
rect 17316 3000 17368 3052
rect 17500 3000 17552 3052
rect 19984 3068 20036 3120
rect 22560 3179 22612 3188
rect 22560 3145 22569 3179
rect 22569 3145 22603 3179
rect 22603 3145 22612 3179
rect 22560 3136 22612 3145
rect 23388 3136 23440 3188
rect 22100 3111 22152 3120
rect 22100 3077 22127 3111
rect 22127 3077 22152 3111
rect 22100 3068 22152 3077
rect 22376 3068 22428 3120
rect 23756 3068 23808 3120
rect 19340 3000 19392 3052
rect 19800 3043 19852 3052
rect 19800 3009 19809 3043
rect 19809 3009 19843 3043
rect 19843 3009 19852 3043
rect 19800 3000 19852 3009
rect 21640 3000 21692 3052
rect 14924 2932 14976 2984
rect 15752 2932 15804 2984
rect 16120 2932 16172 2984
rect 17224 2932 17276 2984
rect 9312 2864 9364 2916
rect 7564 2796 7616 2848
rect 7748 2796 7800 2848
rect 9036 2796 9088 2848
rect 9956 2839 10008 2848
rect 9956 2805 9965 2839
rect 9965 2805 9999 2839
rect 9999 2805 10008 2839
rect 9956 2796 10008 2805
rect 10968 2864 11020 2916
rect 11336 2864 11388 2916
rect 14832 2864 14884 2916
rect 19616 2864 19668 2916
rect 13544 2796 13596 2848
rect 15016 2796 15068 2848
rect 15476 2796 15528 2848
rect 17684 2796 17736 2848
rect 18236 2796 18288 2848
rect 18972 2796 19024 2848
rect 19524 2796 19576 2848
rect 20628 2932 20680 2984
rect 20812 2932 20864 2984
rect 21272 2932 21324 2984
rect 21180 2796 21232 2848
rect 23940 2932 23992 2984
rect 24032 2796 24084 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 12214 2694 12266 2746
rect 12278 2694 12330 2746
rect 12342 2694 12394 2746
rect 12406 2694 12458 2746
rect 12470 2694 12522 2746
rect 20214 2694 20266 2746
rect 20278 2694 20330 2746
rect 20342 2694 20394 2746
rect 20406 2694 20458 2746
rect 20470 2694 20522 2746
rect 3148 2592 3200 2644
rect 2780 2524 2832 2576
rect 6552 2592 6604 2644
rect 7196 2592 7248 2644
rect 2688 2499 2740 2508
rect 2688 2465 2697 2499
rect 2697 2465 2731 2499
rect 2731 2465 2740 2499
rect 2688 2456 2740 2465
rect 1308 2320 1360 2372
rect 2320 2431 2372 2440
rect 2320 2397 2329 2431
rect 2329 2397 2363 2431
rect 2363 2397 2372 2431
rect 2320 2388 2372 2397
rect 3056 2388 3108 2440
rect 3332 2388 3384 2440
rect 2872 2320 2924 2372
rect 3976 2431 4028 2440
rect 3976 2397 3985 2431
rect 3985 2397 4019 2431
rect 4019 2397 4028 2431
rect 3976 2388 4028 2397
rect 7748 2524 7800 2576
rect 10692 2592 10744 2644
rect 11520 2592 11572 2644
rect 17776 2592 17828 2644
rect 17960 2592 18012 2644
rect 18788 2592 18840 2644
rect 20076 2592 20128 2644
rect 22468 2592 22520 2644
rect 5356 2456 5408 2508
rect 4804 2388 4856 2440
rect 5724 2388 5776 2440
rect 6736 2499 6788 2508
rect 6736 2465 6745 2499
rect 6745 2465 6779 2499
rect 6779 2465 6788 2499
rect 6736 2456 6788 2465
rect 7840 2499 7892 2508
rect 7840 2465 7849 2499
rect 7849 2465 7883 2499
rect 7883 2465 7892 2499
rect 7840 2456 7892 2465
rect 8116 2456 8168 2508
rect 9036 2524 9088 2576
rect 8852 2456 8904 2508
rect 9864 2456 9916 2508
rect 12624 2524 12676 2576
rect 13176 2524 13228 2576
rect 14004 2524 14056 2576
rect 6828 2431 6880 2440
rect 6828 2397 6837 2431
rect 6837 2397 6871 2431
rect 6871 2397 6880 2431
rect 6828 2388 6880 2397
rect 7012 2388 7064 2440
rect 7656 2388 7708 2440
rect 7932 2431 7984 2440
rect 7932 2397 7941 2431
rect 7941 2397 7975 2431
rect 7975 2397 7984 2431
rect 7932 2388 7984 2397
rect 8024 2388 8076 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 6644 2252 6696 2304
rect 8116 2320 8168 2372
rect 9036 2252 9088 2304
rect 9680 2252 9732 2304
rect 10416 2252 10468 2304
rect 10692 2388 10744 2440
rect 11152 2431 11204 2440
rect 11152 2397 11161 2431
rect 11161 2397 11195 2431
rect 11195 2397 11204 2431
rect 11152 2388 11204 2397
rect 11336 2320 11388 2372
rect 12624 2388 12676 2440
rect 12992 2388 13044 2440
rect 14740 2499 14792 2508
rect 14740 2465 14749 2499
rect 14749 2465 14783 2499
rect 14783 2465 14792 2499
rect 14740 2456 14792 2465
rect 15384 2456 15436 2508
rect 18696 2567 18748 2576
rect 18696 2533 18705 2567
rect 18705 2533 18739 2567
rect 18739 2533 18748 2567
rect 18696 2524 18748 2533
rect 15936 2456 15988 2508
rect 16672 2499 16724 2508
rect 16672 2465 16681 2499
rect 16681 2465 16715 2499
rect 16715 2465 16724 2499
rect 16672 2456 16724 2465
rect 16856 2456 16908 2508
rect 17040 2456 17092 2508
rect 17224 2499 17276 2508
rect 17224 2465 17233 2499
rect 17233 2465 17267 2499
rect 17267 2465 17276 2499
rect 17224 2456 17276 2465
rect 17592 2456 17644 2508
rect 17776 2456 17828 2508
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 15752 2431 15804 2440
rect 15752 2397 15761 2431
rect 15761 2397 15795 2431
rect 15795 2397 15804 2431
rect 15752 2388 15804 2397
rect 16028 2431 16080 2440
rect 16028 2397 16037 2431
rect 16037 2397 16071 2431
rect 16071 2397 16080 2431
rect 16028 2388 16080 2397
rect 12808 2320 12860 2372
rect 15936 2363 15988 2372
rect 15936 2329 15945 2363
rect 15945 2329 15979 2363
rect 15979 2329 15988 2363
rect 15936 2320 15988 2329
rect 17684 2388 17736 2440
rect 18144 2388 18196 2440
rect 19248 2388 19300 2440
rect 17592 2320 17644 2372
rect 18972 2363 19024 2372
rect 18972 2329 18981 2363
rect 18981 2329 19015 2363
rect 19015 2329 19024 2363
rect 18972 2320 19024 2329
rect 11428 2252 11480 2304
rect 11980 2252 12032 2304
rect 15476 2252 15528 2304
rect 20904 2524 20956 2576
rect 19524 2499 19576 2508
rect 19524 2465 19533 2499
rect 19533 2465 19567 2499
rect 19567 2465 19576 2499
rect 19524 2456 19576 2465
rect 22560 2456 22612 2508
rect 23112 2456 23164 2508
rect 19616 2388 19668 2440
rect 20628 2431 20680 2440
rect 20628 2397 20637 2431
rect 20637 2397 20671 2431
rect 20671 2397 20680 2431
rect 20628 2388 20680 2397
rect 22192 2388 22244 2440
rect 23020 2388 23072 2440
rect 21088 2320 21140 2372
rect 20076 2252 20128 2304
rect 8214 2150 8266 2202
rect 8278 2150 8330 2202
rect 8342 2150 8394 2202
rect 8406 2150 8458 2202
rect 8470 2150 8522 2202
rect 16214 2150 16266 2202
rect 16278 2150 16330 2202
rect 16342 2150 16394 2202
rect 16406 2150 16458 2202
rect 16470 2150 16522 2202
rect 24214 2150 24266 2202
rect 24278 2150 24330 2202
rect 24342 2150 24394 2202
rect 24406 2150 24458 2202
rect 24470 2150 24522 2202
rect 1584 2048 1636 2100
rect 3976 2091 4028 2100
rect 3976 2057 3985 2091
rect 3985 2057 4019 2091
rect 4019 2057 4028 2091
rect 3976 2048 4028 2057
rect 4804 2048 4856 2100
rect 5172 2091 5224 2100
rect 5172 2057 5197 2091
rect 5197 2057 5224 2091
rect 5172 2048 5224 2057
rect 1952 1980 2004 2032
rect 2688 1980 2740 2032
rect 5448 1980 5500 2032
rect 3240 1955 3292 1964
rect 3240 1921 3249 1955
rect 3249 1921 3283 1955
rect 3283 1921 3292 1955
rect 3240 1912 3292 1921
rect 3332 1912 3384 1964
rect 5080 1912 5132 1964
rect 2320 1844 2372 1896
rect 6736 2023 6788 2032
rect 6736 1989 6745 2023
rect 6745 1989 6779 2023
rect 6779 1989 6788 2023
rect 6736 1980 6788 1989
rect 7564 1980 7616 2032
rect 9036 2048 9088 2100
rect 10140 2048 10192 2100
rect 11612 2048 11664 2100
rect 11980 2048 12032 2100
rect 9680 1980 9732 2032
rect 14096 2048 14148 2100
rect 5632 1887 5684 1896
rect 5632 1853 5641 1887
rect 5641 1853 5675 1887
rect 5675 1853 5684 1887
rect 5632 1844 5684 1853
rect 3884 1776 3936 1828
rect 7380 1955 7432 1964
rect 7380 1921 7389 1955
rect 7389 1921 7423 1955
rect 7423 1921 7432 1955
rect 7380 1912 7432 1921
rect 9588 1912 9640 1964
rect 3148 1708 3200 1760
rect 3608 1751 3660 1760
rect 3608 1717 3617 1751
rect 3617 1717 3651 1751
rect 3651 1717 3660 1751
rect 6736 1819 6788 1828
rect 6736 1785 6745 1819
rect 6745 1785 6779 1819
rect 6779 1785 6788 1819
rect 6736 1776 6788 1785
rect 7104 1844 7156 1896
rect 8116 1844 8168 1896
rect 9680 1844 9732 1896
rect 10048 1955 10100 1964
rect 10048 1921 10057 1955
rect 10057 1921 10091 1955
rect 10091 1921 10100 1955
rect 10048 1912 10100 1921
rect 11060 1912 11112 1964
rect 11152 1912 11204 1964
rect 12072 1912 12124 1964
rect 7472 1776 7524 1828
rect 3608 1708 3660 1717
rect 5172 1751 5224 1760
rect 5172 1717 5181 1751
rect 5181 1717 5215 1751
rect 5215 1717 5224 1751
rect 5172 1708 5224 1717
rect 7012 1708 7064 1760
rect 7104 1708 7156 1760
rect 9680 1708 9732 1760
rect 9956 1708 10008 1760
rect 11796 1708 11848 1760
rect 12072 1776 12124 1828
rect 13268 1776 13320 1828
rect 13544 1955 13596 1964
rect 13544 1921 13553 1955
rect 13553 1921 13587 1955
rect 13587 1921 13596 1955
rect 13544 1912 13596 1921
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 14280 1912 14332 1964
rect 14740 1912 14792 1964
rect 17868 2048 17920 2100
rect 18696 2048 18748 2100
rect 19064 2048 19116 2100
rect 15476 1980 15528 2032
rect 16580 1980 16632 2032
rect 17040 2023 17092 2032
rect 17040 1989 17049 2023
rect 17049 1989 17083 2023
rect 17083 1989 17092 2023
rect 17040 1980 17092 1989
rect 17500 1980 17552 2032
rect 18420 1980 18472 2032
rect 20720 1980 20772 2032
rect 15568 1912 15620 1964
rect 16764 1955 16816 1964
rect 16764 1921 16773 1955
rect 16773 1921 16807 1955
rect 16807 1921 16816 1955
rect 16764 1912 16816 1921
rect 18788 1844 18840 1896
rect 13636 1776 13688 1828
rect 15200 1776 15252 1828
rect 18144 1776 18196 1828
rect 13820 1708 13872 1760
rect 15936 1708 15988 1760
rect 19892 1844 19944 1896
rect 19984 1844 20036 1896
rect 23664 2048 23716 2100
rect 23848 1980 23900 2032
rect 23756 1955 23808 1964
rect 23756 1921 23765 1955
rect 23765 1921 23799 1955
rect 23799 1921 23808 1955
rect 23756 1912 23808 1921
rect 19800 1708 19852 1760
rect 22100 1844 22152 1896
rect 24768 2048 24820 2100
rect 24676 1980 24728 2032
rect 20812 1708 20864 1760
rect 22008 1751 22060 1760
rect 22008 1717 22017 1751
rect 22017 1717 22051 1751
rect 22051 1717 22060 1751
rect 22008 1708 22060 1717
rect 23940 1708 23992 1760
rect 4214 1606 4266 1658
rect 4278 1606 4330 1658
rect 4342 1606 4394 1658
rect 4406 1606 4458 1658
rect 4470 1606 4522 1658
rect 12214 1606 12266 1658
rect 12278 1606 12330 1658
rect 12342 1606 12394 1658
rect 12406 1606 12458 1658
rect 12470 1606 12522 1658
rect 20214 1606 20266 1658
rect 20278 1606 20330 1658
rect 20342 1606 20394 1658
rect 20406 1606 20458 1658
rect 20470 1606 20522 1658
rect 1952 1547 2004 1556
rect 1952 1513 1961 1547
rect 1961 1513 1995 1547
rect 1995 1513 2004 1547
rect 1952 1504 2004 1513
rect 2228 1504 2280 1556
rect 5172 1504 5224 1556
rect 7288 1504 7340 1556
rect 7472 1504 7524 1556
rect 7840 1504 7892 1556
rect 8668 1504 8720 1556
rect 9496 1504 9548 1556
rect 10692 1504 10744 1556
rect 10784 1547 10836 1556
rect 10784 1513 10793 1547
rect 10793 1513 10827 1547
rect 10827 1513 10836 1547
rect 10784 1504 10836 1513
rect 3056 1479 3108 1488
rect 3056 1445 3065 1479
rect 3065 1445 3099 1479
rect 3099 1445 3108 1479
rect 3056 1436 3108 1445
rect 3332 1436 3384 1488
rect 1584 1368 1636 1420
rect 1492 1343 1544 1352
rect 1492 1309 1501 1343
rect 1501 1309 1535 1343
rect 1535 1309 1544 1343
rect 1492 1300 1544 1309
rect 1676 1300 1728 1352
rect 2136 1275 2188 1284
rect 2136 1241 2163 1275
rect 2163 1241 2188 1275
rect 2136 1232 2188 1241
rect 3608 1300 3660 1352
rect 3884 1368 3936 1420
rect 4068 1300 4120 1352
rect 4620 1368 4672 1420
rect 4804 1300 4856 1352
rect 5172 1343 5224 1352
rect 5172 1309 5181 1343
rect 5181 1309 5215 1343
rect 5215 1309 5224 1343
rect 5172 1300 5224 1309
rect 7196 1436 7248 1488
rect 7380 1436 7432 1488
rect 15936 1504 15988 1556
rect 17132 1504 17184 1556
rect 17408 1504 17460 1556
rect 17592 1504 17644 1556
rect 18236 1504 18288 1556
rect 18788 1547 18840 1556
rect 18788 1513 18797 1547
rect 18797 1513 18831 1547
rect 18831 1513 18840 1547
rect 18788 1504 18840 1513
rect 20076 1547 20128 1556
rect 20076 1513 20106 1547
rect 20106 1513 20128 1547
rect 20076 1504 20128 1513
rect 21088 1504 21140 1556
rect 21916 1547 21968 1556
rect 21916 1513 21925 1547
rect 21925 1513 21959 1547
rect 21959 1513 21968 1547
rect 21916 1504 21968 1513
rect 22008 1504 22060 1556
rect 11980 1436 12032 1488
rect 12072 1436 12124 1488
rect 16028 1436 16080 1488
rect 1676 1207 1728 1216
rect 1676 1173 1685 1207
rect 1685 1173 1719 1207
rect 1719 1173 1728 1207
rect 1676 1164 1728 1173
rect 3608 1164 3660 1216
rect 3976 1232 4028 1284
rect 6828 1368 6880 1420
rect 7932 1368 7984 1420
rect 6092 1300 6144 1352
rect 6368 1300 6420 1352
rect 6000 1232 6052 1284
rect 7840 1343 7892 1352
rect 7840 1309 7849 1343
rect 7849 1309 7883 1343
rect 7883 1309 7892 1343
rect 7840 1300 7892 1309
rect 9588 1300 9640 1352
rect 9956 1343 10008 1352
rect 9956 1309 9965 1343
rect 9965 1309 9999 1343
rect 9999 1309 10008 1343
rect 9956 1300 10008 1309
rect 10876 1368 10928 1420
rect 13176 1411 13228 1420
rect 13176 1377 13185 1411
rect 13185 1377 13219 1411
rect 13219 1377 13228 1411
rect 13176 1368 13228 1377
rect 14740 1368 14792 1420
rect 15200 1368 15252 1420
rect 17408 1368 17460 1420
rect 11060 1343 11112 1352
rect 11060 1309 11069 1343
rect 11069 1309 11103 1343
rect 11103 1309 11112 1343
rect 11060 1300 11112 1309
rect 11520 1300 11572 1352
rect 11888 1300 11940 1352
rect 11980 1300 12032 1352
rect 12624 1300 12676 1352
rect 12716 1300 12768 1352
rect 13452 1300 13504 1352
rect 14004 1300 14056 1352
rect 15752 1343 15804 1352
rect 15752 1309 15761 1343
rect 15761 1309 15795 1343
rect 15795 1309 15804 1343
rect 15752 1300 15804 1309
rect 4620 1164 4672 1216
rect 5632 1164 5684 1216
rect 8576 1275 8628 1284
rect 8576 1241 8585 1275
rect 8585 1241 8619 1275
rect 8619 1241 8628 1275
rect 8576 1232 8628 1241
rect 8760 1232 8812 1284
rect 13820 1232 13872 1284
rect 14280 1232 14332 1284
rect 16856 1275 16908 1284
rect 16856 1241 16865 1275
rect 16865 1241 16899 1275
rect 16899 1241 16908 1275
rect 16856 1232 16908 1241
rect 16948 1232 17000 1284
rect 17316 1300 17368 1352
rect 17684 1343 17736 1352
rect 17684 1309 17705 1343
rect 17705 1309 17736 1343
rect 17684 1300 17736 1309
rect 18696 1300 18748 1352
rect 18972 1343 19024 1352
rect 18972 1309 18981 1343
rect 18981 1309 19015 1343
rect 19015 1309 19024 1343
rect 18972 1300 19024 1309
rect 19340 1343 19392 1352
rect 19340 1309 19349 1343
rect 19349 1309 19383 1343
rect 19383 1309 19392 1343
rect 19340 1300 19392 1309
rect 19800 1411 19852 1420
rect 19800 1377 19809 1411
rect 19809 1377 19843 1411
rect 19843 1377 19852 1411
rect 19800 1368 19852 1377
rect 23756 1368 23808 1420
rect 22100 1343 22152 1352
rect 22100 1309 22109 1343
rect 22109 1309 22143 1343
rect 22143 1309 22152 1343
rect 22100 1300 22152 1309
rect 22744 1300 22796 1352
rect 17868 1232 17920 1284
rect 6644 1207 6696 1216
rect 6644 1173 6653 1207
rect 6653 1173 6687 1207
rect 6687 1173 6696 1207
rect 6644 1164 6696 1173
rect 14004 1164 14056 1216
rect 18420 1164 18472 1216
rect 20076 1232 20128 1284
rect 19064 1164 19116 1216
rect 19984 1164 20036 1216
rect 8214 1062 8266 1114
rect 8278 1062 8330 1114
rect 8342 1062 8394 1114
rect 8406 1062 8458 1114
rect 8470 1062 8522 1114
rect 16214 1062 16266 1114
rect 16278 1062 16330 1114
rect 16342 1062 16394 1114
rect 16406 1062 16458 1114
rect 16470 1062 16522 1114
rect 24214 1062 24266 1114
rect 24278 1062 24330 1114
rect 24342 1062 24394 1114
rect 24406 1062 24458 1114
rect 24470 1062 24522 1114
rect 1676 960 1728 1012
rect 13084 960 13136 1012
rect 18512 960 18564 1012
rect 20076 960 20128 1012
rect 6644 892 6696 944
rect 13728 892 13780 944
rect 18236 892 18288 944
rect 21456 892 21508 944
rect 22100 892 22152 944
rect 4804 824 4856 876
rect 6460 824 6512 876
rect 7564 824 7616 876
rect 8576 824 8628 876
rect 19340 824 19392 876
rect 19708 756 19760 808
rect 17684 688 17736 740
rect 19340 688 19392 740
<< metal2 >>
rect 1306 19200 1362 20000
rect 3882 19200 3938 20000
rect 6458 19200 6514 20000
rect 9034 19200 9090 20000
rect 11610 19200 11666 20000
rect 13820 19304 13872 19310
rect 13820 19246 13872 19252
rect 1320 18290 1348 19200
rect 2962 18592 3018 18601
rect 2962 18527 3018 18536
rect 1860 18352 1912 18358
rect 1860 18294 1912 18300
rect 2412 18352 2464 18358
rect 2412 18294 2464 18300
rect 1308 18284 1360 18290
rect 1308 18226 1360 18232
rect 1676 18080 1728 18086
rect 1676 18022 1728 18028
rect 1688 17882 1716 18022
rect 1676 17876 1728 17882
rect 1676 17818 1728 17824
rect 1872 17270 1900 18294
rect 1952 17604 2004 17610
rect 1952 17546 2004 17552
rect 1964 17338 1992 17546
rect 1952 17332 2004 17338
rect 1952 17274 2004 17280
rect 2424 17270 2452 18294
rect 2976 18290 3004 18527
rect 3896 18290 3924 19200
rect 2964 18284 3016 18290
rect 2964 18226 3016 18232
rect 3884 18284 3936 18290
rect 3884 18226 3936 18232
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2596 18080 2648 18086
rect 2596 18022 2648 18028
rect 1860 17264 1912 17270
rect 2412 17264 2464 17270
rect 1860 17206 1912 17212
rect 2332 17212 2412 17218
rect 2332 17206 2464 17212
rect 1872 17082 1900 17206
rect 2332 17190 2452 17206
rect 1872 17054 2084 17082
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1768 16516 1820 16522
rect 1768 16458 1820 16464
rect 1780 16250 1808 16458
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1490 16144 1546 16153
rect 1490 16079 1492 16088
rect 1544 16079 1546 16088
rect 1492 16050 1544 16056
rect 1400 15360 1452 15366
rect 1400 15302 1452 15308
rect 1768 15360 1820 15366
rect 1768 15302 1820 15308
rect 1412 15026 1440 15302
rect 1400 15020 1452 15026
rect 1400 14962 1452 14968
rect 1412 14249 1440 14962
rect 1492 14476 1544 14482
rect 1492 14418 1544 14424
rect 1398 14240 1454 14249
rect 1398 14175 1454 14184
rect 1504 13938 1532 14418
rect 1780 14346 1808 15302
rect 1964 14822 1992 16934
rect 2056 16574 2084 17054
rect 2056 16546 2176 16574
rect 2148 16182 2176 16546
rect 2136 16176 2188 16182
rect 2136 16118 2188 16124
rect 2044 15156 2096 15162
rect 2044 15098 2096 15104
rect 1952 14816 2004 14822
rect 1952 14758 2004 14764
rect 1768 14340 1820 14346
rect 1768 14282 1820 14288
rect 1492 13932 1544 13938
rect 1492 13874 1544 13880
rect 1860 13864 1912 13870
rect 1860 13806 1912 13812
rect 1872 13462 1900 13806
rect 1964 13734 1992 14758
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 1964 13530 1992 13670
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1860 13456 1912 13462
rect 1860 13398 1912 13404
rect 1964 13394 1992 13466
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 1860 13252 1912 13258
rect 1860 13194 1912 13200
rect 1308 13184 1360 13190
rect 1308 13126 1360 13132
rect 1320 12850 1348 13126
rect 1872 12918 1900 13194
rect 2056 13190 2084 15098
rect 2148 15094 2176 16118
rect 2332 15162 2360 17190
rect 2516 16998 2544 18022
rect 2608 17610 2636 18022
rect 4208 17978 4528 18544
rect 6472 18290 6500 19200
rect 8208 18522 8528 18544
rect 8208 18470 8214 18522
rect 8266 18470 8278 18522
rect 8330 18470 8342 18522
rect 8394 18470 8406 18522
rect 8458 18470 8470 18522
rect 8522 18470 8528 18522
rect 5264 18284 5316 18290
rect 5264 18226 5316 18232
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 5172 18148 5224 18154
rect 5172 18090 5224 18096
rect 4620 18080 4672 18086
rect 4620 18022 4672 18028
rect 4208 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 4528 17978
rect 4068 17672 4120 17678
rect 4068 17614 4120 17620
rect 2596 17604 2648 17610
rect 2596 17546 2648 17552
rect 3332 17536 3384 17542
rect 3332 17478 3384 17484
rect 3344 17338 3372 17478
rect 2872 17332 2924 17338
rect 2872 17274 2924 17280
rect 3332 17332 3384 17338
rect 3332 17274 3384 17280
rect 2780 17060 2832 17066
rect 2780 17002 2832 17008
rect 2504 16992 2556 16998
rect 2504 16934 2556 16940
rect 2792 16522 2820 17002
rect 2780 16516 2832 16522
rect 2780 16458 2832 16464
rect 2688 16448 2740 16454
rect 2688 16390 2740 16396
rect 2700 16250 2728 16390
rect 2884 16250 2912 17274
rect 3976 17128 4028 17134
rect 4080 17082 4108 17614
rect 4028 17076 4108 17082
rect 3976 17070 4108 17076
rect 3988 17054 4108 17070
rect 4080 16658 4108 17054
rect 4208 16890 4528 17926
rect 4632 17746 4660 18022
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4208 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 4528 16890
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 3056 16516 3108 16522
rect 3056 16458 3108 16464
rect 2688 16244 2740 16250
rect 2688 16186 2740 16192
rect 2872 16244 2924 16250
rect 2872 16186 2924 16192
rect 2700 15570 2728 16186
rect 2872 16108 2924 16114
rect 3068 16096 3096 16458
rect 4080 16182 4108 16594
rect 4068 16176 4120 16182
rect 4068 16118 4120 16124
rect 2924 16068 3096 16096
rect 2872 16050 2924 16056
rect 2688 15564 2740 15570
rect 2688 15506 2740 15512
rect 2688 15360 2740 15366
rect 2688 15302 2740 15308
rect 2320 15156 2372 15162
rect 2320 15098 2372 15104
rect 2136 15088 2188 15094
rect 2136 15030 2188 15036
rect 2148 14074 2176 15030
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 14346 2544 14758
rect 2504 14340 2556 14346
rect 2504 14282 2556 14288
rect 2700 14278 2728 15302
rect 4080 15162 4108 16118
rect 4208 15802 4528 16838
rect 4724 16794 4752 17070
rect 4712 16788 4764 16794
rect 4712 16730 4764 16736
rect 4816 16726 4844 17206
rect 4988 16992 5040 16998
rect 4988 16934 5040 16940
rect 4804 16720 4856 16726
rect 4804 16662 4856 16668
rect 5000 16658 5028 16934
rect 4988 16652 5040 16658
rect 4988 16594 5040 16600
rect 5000 16250 5028 16594
rect 5080 16448 5132 16454
rect 5080 16390 5132 16396
rect 5092 16250 5120 16390
rect 4988 16244 5040 16250
rect 4988 16186 5040 16192
rect 5080 16244 5132 16250
rect 5080 16186 5132 16192
rect 4620 16040 4672 16046
rect 4620 15982 4672 15988
rect 4208 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 4528 15802
rect 4068 15156 4120 15162
rect 4068 15098 4120 15104
rect 3976 15088 4028 15094
rect 3976 15030 4028 15036
rect 2964 15020 3016 15026
rect 2964 14962 3016 14968
rect 2976 14482 3004 14962
rect 3884 14952 3936 14958
rect 3884 14894 3936 14900
rect 3896 14618 3924 14894
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 2964 14476 3016 14482
rect 2964 14418 3016 14424
rect 2688 14272 2740 14278
rect 2688 14214 2740 14220
rect 3332 14272 3384 14278
rect 3332 14214 3384 14220
rect 2136 14068 2188 14074
rect 2136 14010 2188 14016
rect 2148 13326 2176 14010
rect 2228 13388 2280 13394
rect 2228 13330 2280 13336
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1860 12912 1912 12918
rect 1860 12854 1912 12860
rect 2056 12866 2084 13126
rect 2136 12912 2188 12918
rect 2056 12860 2136 12866
rect 2056 12854 2188 12860
rect 1308 12844 1360 12850
rect 1308 12786 1360 12792
rect 1320 12073 1348 12786
rect 1492 12232 1544 12238
rect 1492 12174 1544 12180
rect 1306 12064 1362 12073
rect 1306 11999 1362 12008
rect 1308 11756 1360 11762
rect 1308 11698 1360 11704
rect 1320 9897 1348 11698
rect 1504 11626 1532 12174
rect 1492 11620 1544 11626
rect 1492 11562 1544 11568
rect 1504 10606 1532 11562
rect 1872 11082 1900 12854
rect 2056 12838 2176 12854
rect 2056 11082 2084 12838
rect 2240 12782 2268 13330
rect 2228 12776 2280 12782
rect 2228 12718 2280 12724
rect 2240 12646 2268 12718
rect 2228 12640 2280 12646
rect 2228 12582 2280 12588
rect 2320 12640 2372 12646
rect 2320 12582 2372 12588
rect 2240 12434 2268 12582
rect 2148 12406 2268 12434
rect 2148 11354 2176 12406
rect 2332 12306 2360 12582
rect 2320 12300 2372 12306
rect 2320 12242 2372 12248
rect 2136 11348 2188 11354
rect 2136 11290 2188 11296
rect 1860 11076 1912 11082
rect 1860 11018 1912 11024
rect 2044 11076 2096 11082
rect 2044 11018 2096 11024
rect 1492 10600 1544 10606
rect 1492 10542 1544 10548
rect 1504 10062 1532 10542
rect 1872 10282 1900 11018
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1964 10742 1992 10950
rect 1952 10736 2004 10742
rect 1952 10678 2004 10684
rect 1872 10266 1992 10282
rect 1872 10260 2004 10266
rect 1872 10254 1952 10260
rect 1492 10056 1544 10062
rect 1492 9998 1544 10004
rect 1306 9888 1362 9897
rect 1306 9823 1362 9832
rect 1504 9450 1532 9998
rect 1872 9654 1900 10254
rect 1952 10202 2004 10208
rect 2056 9654 2084 11018
rect 1860 9648 1912 9654
rect 1860 9590 1912 9596
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 1492 9444 1544 9450
rect 1492 9386 1544 9392
rect 1504 8974 1532 9386
rect 2148 9382 2176 11290
rect 2504 10124 2556 10130
rect 2504 10066 2556 10072
rect 2516 9722 2544 10066
rect 2504 9716 2556 9722
rect 2504 9658 2556 9664
rect 2136 9376 2188 9382
rect 2136 9318 2188 9324
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1400 7880 1452 7886
rect 1400 7822 1452 7828
rect 1412 7721 1440 7822
rect 1398 7712 1454 7721
rect 1398 7647 1454 7656
rect 1504 7342 1532 8910
rect 2136 8900 2188 8906
rect 2136 8842 2188 8848
rect 2148 8634 2176 8842
rect 2228 8832 2280 8838
rect 2228 8774 2280 8780
rect 2504 8832 2556 8838
rect 2504 8774 2556 8780
rect 2240 8634 2268 8774
rect 2136 8628 2188 8634
rect 2136 8570 2188 8576
rect 2228 8628 2280 8634
rect 2228 8570 2280 8576
rect 1584 8560 1636 8566
rect 1584 8502 1636 8508
rect 1492 7336 1544 7342
rect 1492 7278 1544 7284
rect 1398 5536 1454 5545
rect 1398 5471 1454 5480
rect 1412 4826 1440 5471
rect 1400 4820 1452 4826
rect 1400 4762 1452 4768
rect 1412 3534 1440 4762
rect 1504 4078 1532 7278
rect 1596 6730 1624 8502
rect 2136 8492 2188 8498
rect 2136 8434 2188 8440
rect 1952 8288 2004 8294
rect 1952 8230 2004 8236
rect 1674 8120 1730 8129
rect 1674 8055 1676 8064
rect 1728 8055 1730 8064
rect 1676 8026 1728 8032
rect 1676 7880 1728 7886
rect 1676 7822 1728 7828
rect 1584 6724 1636 6730
rect 1584 6666 1636 6672
rect 1596 5114 1624 6666
rect 1688 5302 1716 7822
rect 1768 7744 1820 7750
rect 1768 7686 1820 7692
rect 1780 5710 1808 7686
rect 1964 7206 1992 8230
rect 1952 7200 2004 7206
rect 1952 7142 2004 7148
rect 1964 7002 1992 7142
rect 1952 6996 2004 7002
rect 1952 6938 2004 6944
rect 1768 5704 1820 5710
rect 1768 5646 1820 5652
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1596 5086 1716 5114
rect 1492 4072 1544 4078
rect 1492 4014 1544 4020
rect 1400 3528 1452 3534
rect 1400 3470 1452 3476
rect 1490 3360 1546 3369
rect 1490 3295 1546 3304
rect 1308 2372 1360 2378
rect 1308 2314 1360 2320
rect 1320 800 1348 2314
rect 1504 1358 1532 3295
rect 1584 3052 1636 3058
rect 1584 2994 1636 3000
rect 1596 2106 1624 2994
rect 1584 2100 1636 2106
rect 1584 2042 1636 2048
rect 1596 1426 1624 2042
rect 1584 1420 1636 1426
rect 1584 1362 1636 1368
rect 1688 1358 1716 5086
rect 1860 4752 1912 4758
rect 1858 4720 1860 4729
rect 1912 4720 1914 4729
rect 1858 4655 1914 4664
rect 1964 4060 1992 6938
rect 2148 6730 2176 8434
rect 2412 7744 2464 7750
rect 2412 7686 2464 7692
rect 2424 7546 2452 7686
rect 2412 7540 2464 7546
rect 2412 7482 2464 7488
rect 2516 7342 2544 8774
rect 2700 7886 2728 14214
rect 3344 14074 3372 14214
rect 3988 14074 4016 15030
rect 4080 14550 4108 15098
rect 4208 14714 4528 15750
rect 4632 15706 4660 15982
rect 4620 15700 4672 15706
rect 4620 15642 4672 15648
rect 5000 15570 5028 16186
rect 4988 15564 5040 15570
rect 4908 15524 4988 15552
rect 4804 15360 4856 15366
rect 4804 15302 4856 15308
rect 4816 15162 4844 15302
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4208 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 4528 14714
rect 4068 14544 4120 14550
rect 4068 14486 4120 14492
rect 3332 14068 3384 14074
rect 3332 14010 3384 14016
rect 3976 14068 4028 14074
rect 3976 14010 4028 14016
rect 2872 14000 2924 14006
rect 2872 13942 2924 13948
rect 2884 13530 2912 13942
rect 2872 13524 2924 13530
rect 2872 13466 2924 13472
rect 3344 13326 3372 14010
rect 4068 13932 4120 13938
rect 4068 13874 4120 13880
rect 3976 13728 4028 13734
rect 3976 13670 4028 13676
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3332 13320 3384 13326
rect 3332 13262 3384 13268
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3148 12776 3200 12782
rect 3148 12718 3200 12724
rect 2780 12708 2832 12714
rect 2780 12650 2832 12656
rect 2792 12170 2820 12650
rect 3160 12238 3188 12718
rect 3148 12232 3200 12238
rect 3148 12174 3200 12180
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 3252 12102 3280 12854
rect 3436 12782 3464 13330
rect 3988 13258 4016 13670
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 3608 13184 3660 13190
rect 3608 13126 3660 13132
rect 3424 12776 3476 12782
rect 3424 12718 3476 12724
rect 3436 12170 3464 12718
rect 3424 12164 3476 12170
rect 3424 12106 3476 12112
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 2964 11280 3016 11286
rect 2964 11222 3016 11228
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2884 10810 2912 10950
rect 2872 10804 2924 10810
rect 2872 10746 2924 10752
rect 2976 10742 3004 11222
rect 3148 11212 3200 11218
rect 3148 11154 3200 11160
rect 2964 10736 3016 10742
rect 2964 10678 3016 10684
rect 2964 9988 3016 9994
rect 2964 9930 3016 9936
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9722 2912 9862
rect 2872 9716 2924 9722
rect 2792 9676 2872 9704
rect 2792 8498 2820 9676
rect 2872 9658 2924 9664
rect 2976 9654 3004 9930
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 3160 9518 3188 11154
rect 3252 11150 3280 12038
rect 3436 11218 3464 12106
rect 3424 11212 3476 11218
rect 3424 11154 3476 11160
rect 3240 11144 3292 11150
rect 3240 11086 3292 11092
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3252 9586 3280 10746
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 3148 9512 3200 9518
rect 3148 9454 3200 9460
rect 3332 8832 3384 8838
rect 3332 8774 3384 8780
rect 3344 8634 3372 8774
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 3332 8628 3384 8634
rect 3332 8570 3384 8576
rect 2780 8492 2832 8498
rect 2780 8434 2832 8440
rect 2884 7954 2912 8570
rect 3620 8566 3648 13126
rect 3700 12640 3752 12646
rect 3700 12582 3752 12588
rect 3712 11762 3740 12582
rect 3884 12096 3936 12102
rect 3884 12038 3936 12044
rect 3896 11898 3924 12038
rect 3884 11892 3936 11898
rect 3884 11834 3936 11840
rect 3700 11756 3752 11762
rect 3700 11698 3752 11704
rect 3608 8560 3660 8566
rect 3608 8502 3660 8508
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3148 8424 3200 8430
rect 3148 8366 3200 8372
rect 3160 8090 3188 8366
rect 3148 8084 3200 8090
rect 3148 8026 3200 8032
rect 3160 7954 3188 8026
rect 2872 7948 2924 7954
rect 2872 7890 2924 7896
rect 3148 7948 3200 7954
rect 3148 7890 3200 7896
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 3160 7426 3188 7890
rect 3240 7744 3292 7750
rect 3240 7686 3292 7692
rect 3252 7546 3280 7686
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 2872 7404 2924 7410
rect 3160 7398 3280 7426
rect 2872 7346 2924 7352
rect 2504 7336 2556 7342
rect 2504 7278 2556 7284
rect 2516 6798 2544 7278
rect 2504 6792 2556 6798
rect 2504 6734 2556 6740
rect 2884 6730 2912 7346
rect 3148 7268 3200 7274
rect 3148 7210 3200 7216
rect 3056 6928 3108 6934
rect 3056 6870 3108 6876
rect 3068 6730 3096 6870
rect 2136 6724 2188 6730
rect 2136 6666 2188 6672
rect 2872 6724 2924 6730
rect 2872 6666 2924 6672
rect 3056 6724 3108 6730
rect 3056 6666 3108 6672
rect 2044 5704 2096 5710
rect 2044 5646 2096 5652
rect 2056 5098 2084 5646
rect 2044 5092 2096 5098
rect 2044 5034 2096 5040
rect 2044 4820 2096 4826
rect 2044 4762 2096 4768
rect 2056 4214 2084 4762
rect 2044 4208 2096 4214
rect 2044 4150 2096 4156
rect 1964 4032 2084 4060
rect 2056 3738 2084 4032
rect 2044 3732 2096 3738
rect 2044 3674 2096 3680
rect 2056 3194 2084 3674
rect 2148 3398 2176 6666
rect 2780 6656 2832 6662
rect 2780 6598 2832 6604
rect 2792 6390 2820 6598
rect 2780 6384 2832 6390
rect 2780 6326 2832 6332
rect 2320 6316 2372 6322
rect 2320 6258 2372 6264
rect 2332 5914 2360 6258
rect 3160 6254 3188 7210
rect 2412 6248 2464 6254
rect 2412 6190 2464 6196
rect 3148 6248 3200 6254
rect 3148 6190 3200 6196
rect 2320 5908 2372 5914
rect 2320 5850 2372 5856
rect 2228 5772 2280 5778
rect 2228 5714 2280 5720
rect 2240 5370 2268 5714
rect 2424 5642 2452 6190
rect 3056 6112 3108 6118
rect 3056 6054 3108 6060
rect 3068 5710 3096 6054
rect 3056 5704 3108 5710
rect 3056 5646 3108 5652
rect 2412 5636 2464 5642
rect 2412 5578 2464 5584
rect 2228 5364 2280 5370
rect 2228 5306 2280 5312
rect 2240 4486 2268 5306
rect 2424 5234 2452 5578
rect 3068 5234 3096 5646
rect 2412 5228 2464 5234
rect 2412 5170 2464 5176
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 2320 5092 2372 5098
rect 2320 5034 2372 5040
rect 2332 4622 2360 5034
rect 2688 4820 2740 4826
rect 2688 4762 2740 4768
rect 2320 4616 2372 4622
rect 2320 4558 2372 4564
rect 2228 4480 2280 4486
rect 2228 4422 2280 4428
rect 2240 3534 2268 4422
rect 2332 3602 2360 4558
rect 2504 4480 2556 4486
rect 2504 4422 2556 4428
rect 2412 4208 2464 4214
rect 2412 4150 2464 4156
rect 2424 3738 2452 4150
rect 2412 3732 2464 3738
rect 2412 3674 2464 3680
rect 2320 3596 2372 3602
rect 2320 3538 2372 3544
rect 2228 3528 2280 3534
rect 2228 3470 2280 3476
rect 2412 3460 2464 3466
rect 2412 3402 2464 3408
rect 2136 3392 2188 3398
rect 2136 3334 2188 3340
rect 2044 3188 2096 3194
rect 2044 3130 2096 3136
rect 1952 2032 2004 2038
rect 1952 1974 2004 1980
rect 1964 1562 1992 1974
rect 1952 1556 2004 1562
rect 1952 1498 2004 1504
rect 1492 1352 1544 1358
rect 1492 1294 1544 1300
rect 1676 1352 1728 1358
rect 1676 1294 1728 1300
rect 2148 1290 2176 3334
rect 2228 3188 2280 3194
rect 2228 3130 2280 3136
rect 2240 1562 2268 3130
rect 2424 3126 2452 3402
rect 2412 3120 2464 3126
rect 2412 3062 2464 3068
rect 2516 2990 2544 4422
rect 2596 3664 2648 3670
rect 2700 3652 2728 4762
rect 2780 4752 2832 4758
rect 2780 4694 2832 4700
rect 2962 4720 3018 4729
rect 2792 4282 2820 4694
rect 2962 4655 2964 4664
rect 3016 4655 3018 4664
rect 2964 4626 3016 4632
rect 3252 4622 3280 7398
rect 3332 5024 3384 5030
rect 3332 4966 3384 4972
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 2872 4480 2924 4486
rect 2872 4422 2924 4428
rect 2780 4276 2832 4282
rect 2780 4218 2832 4224
rect 2648 3624 2728 3652
rect 2596 3606 2648 3612
rect 2504 2984 2556 2990
rect 2504 2926 2556 2932
rect 2320 2848 2372 2854
rect 2320 2790 2372 2796
rect 2780 2848 2832 2854
rect 2780 2790 2832 2796
rect 2332 2446 2360 2790
rect 2792 2582 2820 2790
rect 2780 2576 2832 2582
rect 2780 2518 2832 2524
rect 2688 2508 2740 2514
rect 2688 2450 2740 2456
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 2332 1902 2360 2382
rect 2700 2038 2728 2450
rect 2884 2378 2912 4422
rect 3148 4072 3200 4078
rect 3148 4014 3200 4020
rect 3160 3602 3188 4014
rect 3344 4010 3372 4966
rect 3332 4004 3384 4010
rect 3332 3946 3384 3952
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3252 3602 3280 3878
rect 3148 3596 3200 3602
rect 3148 3538 3200 3544
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3056 3460 3108 3466
rect 3056 3402 3108 3408
rect 3068 3126 3096 3402
rect 3056 3120 3108 3126
rect 3056 3062 3108 3068
rect 3160 3058 3188 3538
rect 3148 3052 3200 3058
rect 3148 2994 3200 3000
rect 3148 2644 3200 2650
rect 3148 2586 3200 2592
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 2688 2032 2740 2038
rect 2688 1974 2740 1980
rect 2320 1896 2372 1902
rect 2320 1838 2372 1844
rect 2228 1556 2280 1562
rect 2228 1498 2280 1504
rect 3068 1494 3096 2382
rect 3160 1766 3188 2586
rect 3252 1970 3280 3538
rect 3344 3534 3372 3946
rect 3332 3528 3384 3534
rect 3332 3470 3384 3476
rect 3344 2990 3372 3470
rect 3332 2984 3384 2990
rect 3332 2926 3384 2932
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 3344 1970 3372 2382
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3148 1760 3200 1766
rect 3148 1702 3200 1708
rect 3344 1494 3372 1906
rect 3056 1488 3108 1494
rect 3056 1430 3108 1436
rect 3332 1488 3384 1494
rect 3332 1430 3384 1436
rect 2136 1284 2188 1290
rect 2136 1226 2188 1232
rect 1676 1216 1728 1222
rect 1676 1158 1728 1164
rect 1688 1018 1716 1158
rect 1676 1012 1728 1018
rect 1676 954 1728 960
rect 3436 800 3464 8434
rect 3620 7954 3648 8502
rect 3792 8356 3844 8362
rect 3844 8316 3924 8344
rect 3792 8298 3844 8304
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3792 7404 3844 7410
rect 3792 7346 3844 7352
rect 3804 6866 3832 7346
rect 3792 6860 3844 6866
rect 3792 6802 3844 6808
rect 3792 6724 3844 6730
rect 3792 6666 3844 6672
rect 3516 6656 3568 6662
rect 3516 6598 3568 6604
rect 3528 6322 3556 6598
rect 3516 6316 3568 6322
rect 3516 6258 3568 6264
rect 3804 5710 3832 6666
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3528 4622 3556 4966
rect 3516 4616 3568 4622
rect 3516 4558 3568 4564
rect 3804 3398 3832 5646
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3792 3392 3844 3398
rect 3792 3334 3844 3340
rect 3712 3233 3740 3334
rect 3698 3224 3754 3233
rect 3698 3159 3754 3168
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 3528 1170 3556 2994
rect 3896 1834 3924 8316
rect 3988 7410 4016 13194
rect 4080 12918 4108 13874
rect 4208 13626 4528 14662
rect 4816 14414 4844 15098
rect 4908 14482 4936 15524
rect 4988 15506 5040 15512
rect 5184 15162 5212 18090
rect 5276 17746 5304 18226
rect 5356 18216 5408 18222
rect 5356 18158 5408 18164
rect 5448 18216 5500 18222
rect 5448 18158 5500 18164
rect 5264 17740 5316 17746
rect 5264 17682 5316 17688
rect 5276 17338 5304 17682
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 5368 17066 5396 18158
rect 5356 17060 5408 17066
rect 5356 17002 5408 17008
rect 5368 16590 5396 17002
rect 5460 16658 5488 18158
rect 7932 18080 7984 18086
rect 7932 18022 7984 18028
rect 5724 17672 5776 17678
rect 5724 17614 5776 17620
rect 5736 16794 5764 17614
rect 7944 17610 7972 18022
rect 7932 17604 7984 17610
rect 7932 17546 7984 17552
rect 7380 17536 7432 17542
rect 7380 17478 7432 17484
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 6828 17196 6880 17202
rect 6828 17138 6880 17144
rect 6736 16992 6788 16998
rect 6736 16934 6788 16940
rect 5724 16788 5776 16794
rect 5724 16730 5776 16736
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 5448 16652 5500 16658
rect 5448 16594 5500 16600
rect 5356 16584 5408 16590
rect 5356 16526 5408 16532
rect 5724 16516 5776 16522
rect 5724 16458 5776 16464
rect 5356 16448 5408 16454
rect 5356 16390 5408 16396
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5276 15706 5304 16050
rect 5368 15978 5396 16390
rect 5356 15972 5408 15978
rect 5356 15914 5408 15920
rect 5264 15700 5316 15706
rect 5264 15642 5316 15648
rect 5368 15502 5396 15914
rect 5448 15904 5500 15910
rect 5448 15846 5500 15852
rect 5460 15638 5488 15846
rect 5448 15632 5500 15638
rect 5448 15574 5500 15580
rect 5356 15496 5408 15502
rect 5356 15438 5408 15444
rect 5736 15434 5764 16458
rect 5920 15706 5948 16730
rect 6748 16590 6776 16934
rect 6840 16794 6868 17138
rect 7392 16998 7420 17478
rect 8128 17338 8156 17478
rect 8208 17434 8528 18470
rect 9048 18290 9076 19200
rect 10876 18420 10928 18426
rect 10876 18362 10928 18368
rect 9680 18352 9732 18358
rect 9680 18294 9732 18300
rect 8852 18284 8904 18290
rect 8852 18226 8904 18232
rect 9036 18284 9088 18290
rect 9036 18226 9088 18232
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8208 17382 8214 17434
rect 8266 17382 8278 17434
rect 8330 17382 8342 17434
rect 8394 17382 8406 17434
rect 8458 17382 8470 17434
rect 8522 17382 8528 17434
rect 8116 17332 8168 17338
rect 8116 17274 8168 17280
rect 7932 17128 7984 17134
rect 7932 17070 7984 17076
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 7392 16658 7420 16934
rect 7944 16794 7972 17070
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7196 16652 7248 16658
rect 7196 16594 7248 16600
rect 7380 16652 7432 16658
rect 7380 16594 7432 16600
rect 6736 16584 6788 16590
rect 6736 16526 6788 16532
rect 6000 16448 6052 16454
rect 6000 16390 6052 16396
rect 5908 15700 5960 15706
rect 5908 15642 5960 15648
rect 5724 15428 5776 15434
rect 5724 15370 5776 15376
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5172 15156 5224 15162
rect 5172 15098 5224 15104
rect 4896 14476 4948 14482
rect 4896 14418 4948 14424
rect 4804 14408 4856 14414
rect 4804 14350 4856 14356
rect 4208 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 4528 13626
rect 4068 12912 4120 12918
rect 4068 12854 4120 12860
rect 4208 12538 4528 13574
rect 4908 13394 4936 14418
rect 5540 14340 5592 14346
rect 5644 14328 5672 15302
rect 5592 14300 5672 14328
rect 5540 14282 5592 14288
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 5736 12918 5764 15370
rect 5920 15178 5948 15642
rect 6012 15502 6040 16390
rect 6748 15502 6776 16526
rect 7104 16448 7156 16454
rect 7104 16390 7156 16396
rect 7116 16250 7144 16390
rect 7104 16244 7156 16250
rect 7104 16186 7156 16192
rect 7104 16108 7156 16114
rect 7104 16050 7156 16056
rect 6000 15496 6052 15502
rect 6000 15438 6052 15444
rect 6736 15496 6788 15502
rect 6736 15438 6788 15444
rect 5828 15150 5948 15178
rect 5828 14822 5856 15150
rect 6012 15094 6040 15438
rect 6828 15428 6880 15434
rect 6828 15370 6880 15376
rect 6736 15360 6788 15366
rect 6736 15302 6788 15308
rect 6000 15088 6052 15094
rect 6000 15030 6052 15036
rect 6012 14906 6040 15030
rect 5920 14878 6040 14906
rect 5816 14816 5868 14822
rect 5816 14758 5868 14764
rect 5724 12912 5776 12918
rect 5724 12854 5776 12860
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4208 12486 4214 12538
rect 4266 12518 4278 12538
rect 4330 12518 4342 12538
rect 4394 12518 4406 12538
rect 4458 12518 4470 12538
rect 4276 12486 4278 12518
rect 4458 12486 4460 12518
rect 4522 12486 4528 12538
rect 4208 12462 4220 12486
rect 4276 12462 4300 12486
rect 4356 12462 4380 12486
rect 4436 12462 4460 12486
rect 4516 12462 4528 12486
rect 4208 12438 4528 12462
rect 4208 12382 4220 12438
rect 4276 12382 4300 12438
rect 4356 12382 4380 12438
rect 4436 12382 4460 12438
rect 4516 12382 4528 12438
rect 4208 12358 4528 12382
rect 4208 12302 4220 12358
rect 4276 12302 4300 12358
rect 4356 12302 4380 12358
rect 4436 12302 4460 12358
rect 4516 12302 4528 12358
rect 4208 12278 4528 12302
rect 4068 12232 4120 12238
rect 4068 12174 4120 12180
rect 4208 12222 4220 12278
rect 4276 12222 4300 12278
rect 4356 12222 4380 12278
rect 4436 12222 4460 12278
rect 4516 12222 4528 12278
rect 4080 11898 4108 12174
rect 4068 11892 4120 11898
rect 4068 11834 4120 11840
rect 4208 11450 4528 12222
rect 4632 11898 4660 12786
rect 4712 12640 4764 12646
rect 4712 12582 4764 12588
rect 4620 11892 4672 11898
rect 4620 11834 4672 11840
rect 4208 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 4528 11450
rect 4208 10362 4528 11398
rect 4208 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 4528 10362
rect 4208 9274 4528 10310
rect 4632 9926 4660 11834
rect 4724 11354 4752 12582
rect 4896 12436 4948 12442
rect 5736 12434 5764 12854
rect 5828 12646 5856 14758
rect 5920 14074 5948 14878
rect 6000 14816 6052 14822
rect 6000 14758 6052 14764
rect 6012 14346 6040 14758
rect 6000 14340 6052 14346
rect 6000 14282 6052 14288
rect 6748 14278 6776 15302
rect 6736 14272 6788 14278
rect 6736 14214 6788 14220
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 5920 12918 5948 14010
rect 6184 13728 6236 13734
rect 6184 13670 6236 13676
rect 6196 13530 6224 13670
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6748 13394 6776 14214
rect 6840 14006 6868 15370
rect 7116 15026 7144 16050
rect 7208 15570 7236 16594
rect 8024 16516 8076 16522
rect 8024 16458 8076 16464
rect 8036 16046 8064 16458
rect 8128 16250 8156 17274
rect 8208 16518 8528 17382
rect 8588 16794 8616 18022
rect 8760 17740 8812 17746
rect 8760 17682 8812 17688
rect 8772 17338 8800 17682
rect 8760 17332 8812 17338
rect 8760 17274 8812 17280
rect 8576 16788 8628 16794
rect 8628 16748 8708 16776
rect 8576 16730 8628 16736
rect 8208 16462 8220 16518
rect 8276 16462 8300 16518
rect 8356 16462 8380 16518
rect 8436 16462 8460 16518
rect 8516 16462 8528 16518
rect 8208 16438 8528 16462
rect 8208 16382 8220 16438
rect 8276 16382 8300 16438
rect 8356 16382 8380 16438
rect 8436 16382 8460 16438
rect 8516 16382 8528 16438
rect 8576 16448 8628 16454
rect 8576 16390 8628 16396
rect 8208 16358 8528 16382
rect 8208 16346 8220 16358
rect 8276 16346 8300 16358
rect 8356 16346 8380 16358
rect 8436 16346 8460 16358
rect 8516 16346 8528 16358
rect 8208 16294 8214 16346
rect 8276 16302 8278 16346
rect 8458 16302 8460 16346
rect 8266 16294 8278 16302
rect 8330 16294 8342 16302
rect 8394 16294 8406 16302
rect 8458 16294 8470 16302
rect 8522 16294 8528 16346
rect 8208 16278 8528 16294
rect 8116 16244 8168 16250
rect 8116 16186 8168 16192
rect 8208 16222 8220 16278
rect 8276 16222 8300 16278
rect 8356 16222 8380 16278
rect 8436 16222 8460 16278
rect 8516 16222 8528 16278
rect 7932 16040 7984 16046
rect 7932 15982 7984 15988
rect 8024 16040 8076 16046
rect 8024 15982 8076 15988
rect 7944 15706 7972 15982
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7196 15564 7248 15570
rect 7196 15506 7248 15512
rect 7932 15360 7984 15366
rect 7932 15302 7984 15308
rect 7656 15088 7708 15094
rect 7656 15030 7708 15036
rect 7012 15020 7064 15026
rect 7012 14962 7064 14968
rect 7104 15020 7156 15026
rect 7104 14962 7156 14968
rect 7024 14346 7052 14962
rect 7116 14482 7144 14962
rect 7668 14618 7696 15030
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 7852 14618 7880 14894
rect 7656 14612 7708 14618
rect 7656 14554 7708 14560
rect 7840 14612 7892 14618
rect 7840 14554 7892 14560
rect 7944 14482 7972 15302
rect 7104 14476 7156 14482
rect 7104 14418 7156 14424
rect 7932 14476 7984 14482
rect 7932 14418 7984 14424
rect 7012 14340 7064 14346
rect 7012 14282 7064 14288
rect 6920 14272 6972 14278
rect 6920 14214 6972 14220
rect 6932 14074 6960 14214
rect 6920 14068 6972 14074
rect 6920 14010 6972 14016
rect 6828 14000 6880 14006
rect 6828 13942 6880 13948
rect 7116 13938 7144 14418
rect 8036 14346 8064 15982
rect 8208 15258 8528 16222
rect 8588 16114 8616 16390
rect 8576 16108 8628 16114
rect 8576 16050 8628 16056
rect 8576 15564 8628 15570
rect 8576 15506 8628 15512
rect 8208 15206 8214 15258
rect 8266 15206 8278 15258
rect 8330 15206 8342 15258
rect 8394 15206 8406 15258
rect 8458 15206 8470 15258
rect 8522 15206 8528 15258
rect 8024 14340 8076 14346
rect 8024 14282 8076 14288
rect 8116 14340 8168 14346
rect 8116 14282 8168 14288
rect 8128 14074 8156 14282
rect 8208 14170 8528 15206
rect 8588 14414 8616 15506
rect 8680 14618 8708 16748
rect 8864 16522 8892 18226
rect 9312 18080 9364 18086
rect 9312 18022 9364 18028
rect 9128 17876 9180 17882
rect 9128 17818 9180 17824
rect 8944 17128 8996 17134
rect 8944 17070 8996 17076
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 8852 16516 8904 16522
rect 8772 16476 8852 16504
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8576 14408 8628 14414
rect 8576 14350 8628 14356
rect 8208 14118 8214 14170
rect 8266 14118 8278 14170
rect 8330 14118 8342 14170
rect 8394 14118 8406 14170
rect 8458 14118 8470 14170
rect 8522 14118 8528 14170
rect 8116 14068 8168 14074
rect 8116 14010 8168 14016
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 6736 13388 6788 13394
rect 6736 13330 6788 13336
rect 5908 12912 5960 12918
rect 5908 12854 5960 12860
rect 6552 12912 6604 12918
rect 6552 12854 6604 12860
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 6184 12640 6236 12646
rect 6184 12582 6236 12588
rect 5736 12406 6040 12434
rect 4896 12378 4948 12384
rect 4908 11354 4936 12378
rect 5172 12164 5224 12170
rect 5172 12106 5224 12112
rect 5184 11898 5212 12106
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5816 12096 5868 12102
rect 5816 12038 5868 12044
rect 5172 11892 5224 11898
rect 5172 11834 5224 11840
rect 5552 11830 5580 12038
rect 5828 11898 5856 12038
rect 5816 11892 5868 11898
rect 5816 11834 5868 11840
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 6012 11762 6040 12406
rect 6196 12170 6224 12582
rect 6564 12434 6592 12854
rect 7116 12782 7144 13874
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7392 13530 7420 13806
rect 7380 13524 7432 13530
rect 7380 13466 7432 13472
rect 8128 13394 8156 14010
rect 8116 13388 8168 13394
rect 8116 13330 8168 13336
rect 8116 13252 8168 13258
rect 8116 13194 8168 13200
rect 7104 12776 7156 12782
rect 7104 12718 7156 12724
rect 6736 12708 6788 12714
rect 6736 12650 6788 12656
rect 6564 12406 6684 12434
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6656 11898 6684 12406
rect 6644 11892 6696 11898
rect 6644 11834 6696 11840
rect 5632 11756 5684 11762
rect 5632 11698 5684 11704
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 4712 11348 4764 11354
rect 4712 11290 4764 11296
rect 4896 11348 4948 11354
rect 4896 11290 4948 11296
rect 4724 10266 4752 11290
rect 5644 10810 5672 11698
rect 5816 11688 5868 11694
rect 5816 11630 5868 11636
rect 6644 11688 6696 11694
rect 6644 11630 6696 11636
rect 5632 10804 5684 10810
rect 5632 10746 5684 10752
rect 5080 10736 5132 10742
rect 5080 10678 5132 10684
rect 5092 10266 5120 10678
rect 5356 10600 5408 10606
rect 5356 10542 5408 10548
rect 5828 10554 5856 11630
rect 5908 11552 5960 11558
rect 5908 11494 5960 11500
rect 5920 11082 5948 11494
rect 6656 11150 6684 11630
rect 6748 11558 6776 12650
rect 7116 12306 7144 12718
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 7472 12300 7524 12306
rect 7472 12242 7524 12248
rect 6920 12096 6972 12102
rect 6920 12038 6972 12044
rect 6736 11552 6788 11558
rect 6736 11494 6788 11500
rect 6932 11218 6960 12038
rect 7116 11694 7144 12242
rect 7484 11898 7512 12242
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7380 11824 7432 11830
rect 7380 11766 7432 11772
rect 7104 11688 7156 11694
rect 7104 11630 7156 11636
rect 7392 11354 7420 11766
rect 7380 11348 7432 11354
rect 7380 11290 7432 11296
rect 7484 11218 7512 11834
rect 8128 11558 8156 13194
rect 8208 13082 8528 14118
rect 8588 13394 8616 14350
rect 8772 14278 8800 16476
rect 8852 16458 8904 16464
rect 8956 16250 8984 17070
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 8956 15502 8984 16186
rect 9048 15570 9076 17070
rect 9036 15564 9088 15570
rect 9036 15506 9088 15512
rect 8944 15496 8996 15502
rect 8944 15438 8996 15444
rect 8852 15360 8904 15366
rect 8852 15302 8904 15308
rect 8864 15162 8892 15302
rect 8852 15156 8904 15162
rect 8852 15098 8904 15104
rect 9140 14482 9168 17818
rect 9324 17202 9352 18022
rect 9312 17196 9364 17202
rect 9312 17138 9364 17144
rect 9692 16182 9720 18294
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9692 16046 9720 16118
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9312 14612 9364 14618
rect 9312 14554 9364 14560
rect 9128 14476 9180 14482
rect 9128 14418 9180 14424
rect 9220 14340 9272 14346
rect 9220 14282 9272 14288
rect 8760 14272 8812 14278
rect 8760 14214 8812 14220
rect 9036 14272 9088 14278
rect 9036 14214 9088 14220
rect 9048 14006 9076 14214
rect 9232 14074 9260 14282
rect 9220 14068 9272 14074
rect 9220 14010 9272 14016
rect 9036 14000 9088 14006
rect 9036 13942 9088 13948
rect 8944 13932 8996 13938
rect 8944 13874 8996 13880
rect 8760 13728 8812 13734
rect 8760 13670 8812 13676
rect 8576 13388 8628 13394
rect 8628 13348 8708 13376
rect 8576 13330 8628 13336
rect 8208 13030 8214 13082
rect 8266 13030 8278 13082
rect 8330 13030 8342 13082
rect 8394 13030 8406 13082
rect 8458 13030 8470 13082
rect 8522 13030 8528 13082
rect 8208 11994 8528 13030
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8588 12102 8616 12854
rect 8680 12646 8708 13348
rect 8668 12640 8720 12646
rect 8668 12582 8720 12588
rect 8680 12238 8708 12582
rect 8668 12232 8720 12238
rect 8668 12174 8720 12180
rect 8576 12096 8628 12102
rect 8576 12038 8628 12044
rect 8208 11942 8214 11994
rect 8266 11942 8278 11994
rect 8330 11942 8342 11994
rect 8394 11942 8406 11994
rect 8458 11942 8470 11994
rect 8522 11942 8528 11994
rect 7748 11552 7800 11558
rect 7748 11494 7800 11500
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 6920 11212 6972 11218
rect 6920 11154 6972 11160
rect 7472 11212 7524 11218
rect 7472 11154 7524 11160
rect 7760 11150 7788 11494
rect 7840 11280 7892 11286
rect 7840 11222 7892 11228
rect 6644 11144 6696 11150
rect 6644 11086 6696 11092
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 5908 11076 5960 11082
rect 5908 11018 5960 11024
rect 6552 10736 6604 10742
rect 6552 10678 6604 10684
rect 5368 10266 5396 10542
rect 5828 10526 5948 10554
rect 5448 10464 5500 10470
rect 5816 10464 5868 10470
rect 5500 10412 5580 10418
rect 5448 10406 5580 10412
rect 5816 10406 5868 10412
rect 5460 10390 5580 10406
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 5080 10260 5132 10266
rect 5080 10202 5132 10208
rect 5356 10260 5408 10266
rect 5356 10202 5408 10208
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 5448 9920 5500 9926
rect 5448 9862 5500 9868
rect 4988 9648 5040 9654
rect 4988 9590 5040 9596
rect 4208 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 4528 9274
rect 4208 8186 4528 9222
rect 5000 9178 5028 9590
rect 5264 9512 5316 9518
rect 5264 9454 5316 9460
rect 5276 9178 5304 9454
rect 4804 9172 4856 9178
rect 4804 9114 4856 9120
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 5264 9172 5316 9178
rect 5264 9114 5316 9120
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4724 8634 4752 8842
rect 4712 8628 4764 8634
rect 4712 8570 4764 8576
rect 4208 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 4528 8186
rect 4068 7948 4120 7954
rect 4068 7890 4120 7896
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3988 6662 4016 7346
rect 3976 6656 4028 6662
rect 3976 6598 4028 6604
rect 3988 5846 4016 6598
rect 3976 5840 4028 5846
rect 3976 5782 4028 5788
rect 4080 5710 4108 7890
rect 4208 7098 4528 8134
rect 4620 7812 4672 7818
rect 4620 7754 4672 7760
rect 4632 7546 4660 7754
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4724 7410 4752 8570
rect 4712 7404 4764 7410
rect 4712 7346 4764 7352
rect 4816 7274 4844 9114
rect 5368 8906 5396 9114
rect 5460 8974 5488 9862
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5356 8900 5408 8906
rect 5356 8842 5408 8848
rect 5552 8838 5580 10390
rect 5828 10130 5856 10406
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5644 9042 5672 9998
rect 5920 9518 5948 10526
rect 6564 10198 6592 10678
rect 6656 10538 6684 11086
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 7024 10606 7052 10950
rect 7012 10600 7064 10606
rect 7012 10542 7064 10548
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6552 10192 6604 10198
rect 6552 10134 6604 10140
rect 6656 10062 6684 10474
rect 6644 10056 6696 10062
rect 6644 9998 6696 10004
rect 6276 9648 6328 9654
rect 6276 9590 6328 9596
rect 5908 9512 5960 9518
rect 5908 9454 5960 9460
rect 5816 9376 5868 9382
rect 5816 9318 5868 9324
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5828 8974 5856 9318
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 5552 8294 5580 8774
rect 5540 8288 5592 8294
rect 5540 8230 5592 8236
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 5172 7404 5224 7410
rect 5172 7346 5224 7352
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4896 7200 4948 7206
rect 4896 7142 4948 7148
rect 4208 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 4528 7098
rect 4208 6010 4528 7046
rect 4208 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 4528 6010
rect 4068 5704 4120 5710
rect 4068 5646 4120 5652
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3988 4622 4016 5170
rect 4208 4922 4528 5958
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4632 5166 4660 5510
rect 4908 5352 4936 7142
rect 4988 6316 5040 6322
rect 4988 6258 5040 6264
rect 5000 5914 5028 6258
rect 4988 5908 5040 5914
rect 4988 5850 5040 5856
rect 4908 5324 5028 5352
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4620 5160 4672 5166
rect 4804 5160 4856 5166
rect 4672 5120 4752 5148
rect 4620 5102 4672 5108
rect 4208 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 4528 4922
rect 4068 4684 4120 4690
rect 4068 4626 4120 4632
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 4080 4146 4108 4626
rect 4208 4518 4528 4870
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4208 4462 4220 4518
rect 4276 4462 4300 4518
rect 4356 4462 4380 4518
rect 4436 4462 4460 4518
rect 4516 4462 4528 4518
rect 4208 4438 4528 4462
rect 4208 4382 4220 4438
rect 4276 4382 4300 4438
rect 4356 4382 4380 4438
rect 4436 4382 4460 4438
rect 4516 4382 4528 4438
rect 4208 4358 4528 4382
rect 4208 4302 4220 4358
rect 4276 4302 4300 4358
rect 4356 4302 4380 4358
rect 4436 4302 4460 4358
rect 4516 4302 4528 4358
rect 4208 4278 4528 4302
rect 4632 4282 4660 4558
rect 4208 4222 4220 4278
rect 4276 4222 4300 4278
rect 4356 4222 4380 4278
rect 4436 4222 4460 4278
rect 4516 4222 4528 4278
rect 3976 4140 4028 4146
rect 3976 4082 4028 4088
rect 4068 4140 4120 4146
rect 4068 4082 4120 4088
rect 3988 3670 4016 4082
rect 4208 3834 4528 4222
rect 4620 4276 4672 4282
rect 4620 4218 4672 4224
rect 4724 4078 4752 5120
rect 4804 5102 4856 5108
rect 4816 4622 4844 5102
rect 4908 4826 4936 5170
rect 4896 4820 4948 4826
rect 4896 4762 4948 4768
rect 4804 4616 4856 4622
rect 4804 4558 4856 4564
rect 4896 4140 4948 4146
rect 4896 4082 4948 4088
rect 4712 4072 4764 4078
rect 4712 4014 4764 4020
rect 4908 3942 4936 4082
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4208 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 4528 3834
rect 3976 3664 4028 3670
rect 3976 3606 4028 3612
rect 3974 3088 4030 3097
rect 3974 3023 3976 3032
rect 4028 3023 4030 3032
rect 3976 2994 4028 3000
rect 4068 2916 4120 2922
rect 4068 2858 4120 2864
rect 3976 2440 4028 2446
rect 3976 2382 4028 2388
rect 3988 2106 4016 2382
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3884 1828 3936 1834
rect 3884 1770 3936 1776
rect 3608 1760 3660 1766
rect 3608 1702 3660 1708
rect 3620 1358 3648 1702
rect 3896 1426 3924 1770
rect 3884 1420 3936 1426
rect 3884 1362 3936 1368
rect 4080 1358 4108 2858
rect 4208 2746 4528 3782
rect 4804 3460 4856 3466
rect 4804 3402 4856 3408
rect 4712 3392 4764 3398
rect 4712 3334 4764 3340
rect 4724 3108 4752 3334
rect 4816 3210 4844 3402
rect 4908 3210 4936 3878
rect 5000 3369 5028 5324
rect 5092 4298 5120 7346
rect 5184 6186 5212 7346
rect 5356 7200 5408 7206
rect 5356 7142 5408 7148
rect 5368 6322 5396 7142
rect 5552 6746 5580 8230
rect 6288 8090 6316 9590
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6368 9512 6420 9518
rect 6368 9454 6420 9460
rect 6380 8974 6408 9454
rect 6368 8968 6420 8974
rect 6368 8910 6420 8916
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6380 8634 6408 8910
rect 6368 8628 6420 8634
rect 6368 8570 6420 8576
rect 6380 8498 6408 8570
rect 6472 8566 6500 8910
rect 6460 8560 6512 8566
rect 6460 8502 6512 8508
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6276 8084 6328 8090
rect 6276 8026 6328 8032
rect 6472 7750 6500 8298
rect 6564 8294 6592 9522
rect 6656 9450 6684 9998
rect 6920 9988 6972 9994
rect 6920 9930 6972 9936
rect 6932 9722 6960 9930
rect 6920 9716 6972 9722
rect 6920 9658 6972 9664
rect 6644 9444 6696 9450
rect 6644 9386 6696 9392
rect 6656 8634 6684 9386
rect 6920 8832 6972 8838
rect 7024 8820 7052 10542
rect 7852 10470 7880 11222
rect 7932 11212 7984 11218
rect 7932 11154 7984 11160
rect 7944 10742 7972 11154
rect 8116 11008 8168 11014
rect 8116 10950 8168 10956
rect 7932 10736 7984 10742
rect 7932 10678 7984 10684
rect 8128 10674 8156 10950
rect 8208 10906 8528 11942
rect 8772 11286 8800 13670
rect 8956 13258 8984 13874
rect 9232 13274 9260 14010
rect 9324 13734 9352 14554
rect 9692 14278 9720 15982
rect 9864 15020 9916 15026
rect 9864 14962 9916 14968
rect 9772 14408 9824 14414
rect 9772 14350 9824 14356
rect 9680 14272 9732 14278
rect 9680 14214 9732 14220
rect 9692 13870 9720 14214
rect 9680 13864 9732 13870
rect 9680 13806 9732 13812
rect 9312 13728 9364 13734
rect 9312 13670 9364 13676
rect 9496 13728 9548 13734
rect 9496 13670 9548 13676
rect 9324 13530 9352 13670
rect 9312 13524 9364 13530
rect 9312 13466 9364 13472
rect 9232 13258 9352 13274
rect 8944 13252 8996 13258
rect 9232 13252 9364 13258
rect 9232 13246 9312 13252
rect 8944 13194 8996 13200
rect 9312 13194 9364 13200
rect 8956 12646 8984 13194
rect 9128 13184 9180 13190
rect 9128 13126 9180 13132
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8760 11280 8812 11286
rect 8760 11222 8812 11228
rect 8668 11076 8720 11082
rect 8668 11018 8720 11024
rect 8208 10854 8214 10906
rect 8266 10854 8278 10906
rect 8330 10854 8342 10906
rect 8394 10854 8406 10906
rect 8458 10854 8470 10906
rect 8522 10854 8528 10906
rect 8116 10668 8168 10674
rect 8116 10610 8168 10616
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7300 10266 7328 10406
rect 7288 10260 7340 10266
rect 7288 10202 7340 10208
rect 7104 9920 7156 9926
rect 7104 9862 7156 9868
rect 7116 9586 7144 9862
rect 7104 9580 7156 9586
rect 7104 9522 7156 9528
rect 7196 9036 7248 9042
rect 7196 8978 7248 8984
rect 7104 8900 7156 8906
rect 7104 8842 7156 8848
rect 6972 8792 7052 8820
rect 6920 8774 6972 8780
rect 6644 8628 6696 8634
rect 6644 8570 6696 8576
rect 6552 8288 6604 8294
rect 6552 8230 6604 8236
rect 6564 7886 6592 8230
rect 6656 7954 6684 8570
rect 6932 8498 6960 8774
rect 6828 8492 6880 8498
rect 6828 8434 6880 8440
rect 6920 8492 6972 8498
rect 6920 8434 6972 8440
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6644 7948 6696 7954
rect 6644 7890 6696 7896
rect 6552 7880 6604 7886
rect 6552 7822 6604 7828
rect 6460 7744 6512 7750
rect 6460 7686 6512 7692
rect 6564 7478 6592 7822
rect 5816 7472 5868 7478
rect 5816 7414 5868 7420
rect 6552 7472 6604 7478
rect 6552 7414 6604 7420
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 5644 6866 5672 7278
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5552 6718 5672 6746
rect 5540 6656 5592 6662
rect 5540 6598 5592 6604
rect 5356 6316 5408 6322
rect 5356 6258 5408 6264
rect 5172 6180 5224 6186
rect 5172 6122 5224 6128
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 5184 5710 5212 6122
rect 5460 5914 5488 6122
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 5172 5704 5224 5710
rect 5172 5646 5224 5652
rect 5264 5024 5316 5030
rect 5264 4966 5316 4972
rect 5092 4270 5212 4298
rect 5184 4026 5212 4270
rect 5276 4146 5304 4966
rect 5460 4622 5488 5850
rect 5552 5846 5580 6598
rect 5644 6254 5672 6718
rect 5632 6248 5684 6254
rect 5632 6190 5684 6196
rect 5540 5840 5592 5846
rect 5540 5782 5592 5788
rect 5552 5710 5580 5782
rect 5736 5710 5764 7142
rect 5828 6934 5856 7414
rect 6840 7410 6868 8434
rect 6920 8356 6972 8362
rect 6920 8298 6972 8304
rect 5908 7404 5960 7410
rect 5908 7346 5960 7352
rect 6092 7404 6144 7410
rect 6092 7346 6144 7352
rect 6644 7404 6696 7410
rect 6644 7346 6696 7352
rect 6828 7404 6880 7410
rect 6828 7346 6880 7352
rect 5816 6928 5868 6934
rect 5816 6870 5868 6876
rect 5828 6730 5856 6870
rect 5920 6798 5948 7346
rect 6104 7002 6132 7346
rect 6368 7268 6420 7274
rect 6368 7210 6420 7216
rect 6092 6996 6144 7002
rect 6092 6938 6144 6944
rect 6092 6860 6144 6866
rect 6012 6820 6092 6848
rect 5908 6792 5960 6798
rect 5908 6734 5960 6740
rect 5816 6724 5868 6730
rect 5816 6666 5868 6672
rect 6012 6322 6040 6820
rect 6092 6802 6144 6808
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 5908 6248 5960 6254
rect 5908 6190 5960 6196
rect 5920 5710 5948 6190
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5724 5704 5776 5710
rect 5724 5646 5776 5652
rect 5908 5704 5960 5710
rect 5908 5646 5960 5652
rect 5540 5296 5592 5302
rect 5540 5238 5592 5244
rect 5552 4690 5580 5238
rect 5540 4684 5592 4690
rect 5540 4626 5592 4632
rect 5448 4616 5500 4622
rect 5448 4558 5500 4564
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5368 4146 5396 4422
rect 5264 4140 5316 4146
rect 5264 4082 5316 4088
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 6012 4078 6040 6258
rect 6092 6112 6144 6118
rect 6092 6054 6144 6060
rect 6000 4072 6052 4078
rect 5184 3998 5304 4026
rect 6000 4014 6052 4020
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5184 3466 5212 3878
rect 5276 3482 5304 3998
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 5276 3454 5856 3482
rect 4986 3360 5042 3369
rect 4986 3295 5042 3304
rect 4816 3182 5028 3210
rect 4804 3120 4856 3126
rect 4724 3080 4804 3108
rect 4620 2984 4672 2990
rect 4620 2926 4672 2932
rect 4208 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 4528 2746
rect 4208 1658 4528 2694
rect 4208 1606 4214 1658
rect 4266 1606 4278 1658
rect 4330 1606 4342 1658
rect 4394 1606 4406 1658
rect 4458 1606 4470 1658
rect 4522 1606 4528 1658
rect 3608 1352 3660 1358
rect 3608 1294 3660 1300
rect 4068 1352 4120 1358
rect 4068 1294 4120 1300
rect 3976 1284 4028 1290
rect 3976 1226 4028 1232
rect 3608 1216 3660 1222
rect 3528 1164 3608 1170
rect 3988 1170 4016 1226
rect 3660 1164 4016 1170
rect 3528 1142 4016 1164
rect 4208 1040 4528 1606
rect 4632 1426 4660 2926
rect 4620 1420 4672 1426
rect 4620 1362 4672 1368
rect 4724 1306 4752 3080
rect 4804 3062 4856 3068
rect 4894 3088 4950 3097
rect 4894 3023 4896 3032
rect 4948 3023 4950 3032
rect 4896 2994 4948 3000
rect 4804 2984 4856 2990
rect 4804 2926 4856 2932
rect 4816 2689 4844 2926
rect 5000 2774 5028 3182
rect 5276 2774 5304 3454
rect 5540 3392 5592 3398
rect 5540 3334 5592 3340
rect 5446 3224 5502 3233
rect 5446 3159 5502 3168
rect 5460 3126 5488 3159
rect 5448 3120 5500 3126
rect 5448 3062 5500 3068
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5000 2746 5120 2774
rect 4802 2680 4858 2689
rect 4802 2615 4858 2624
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4816 2106 4844 2382
rect 4804 2100 4856 2106
rect 4804 2042 4856 2048
rect 5092 1970 5120 2746
rect 5184 2746 5304 2774
rect 5184 2106 5212 2746
rect 5368 2514 5396 2858
rect 5356 2508 5408 2514
rect 5356 2450 5408 2456
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 5460 2038 5488 3062
rect 5448 2032 5500 2038
rect 5448 1974 5500 1980
rect 5080 1964 5132 1970
rect 5080 1906 5132 1912
rect 5172 1760 5224 1766
rect 5172 1702 5224 1708
rect 5184 1562 5212 1702
rect 5172 1556 5224 1562
rect 5172 1498 5224 1504
rect 5170 1456 5226 1465
rect 5170 1391 5226 1400
rect 5184 1358 5212 1391
rect 4632 1278 4752 1306
rect 4804 1352 4856 1358
rect 4804 1294 4856 1300
rect 5172 1352 5224 1358
rect 5172 1294 5224 1300
rect 4632 1222 4660 1278
rect 4620 1216 4672 1222
rect 4620 1158 4672 1164
rect 4816 882 4844 1294
rect 4804 876 4856 882
rect 4804 818 4856 824
rect 5552 800 5580 3334
rect 5828 3233 5856 3454
rect 6012 3398 6040 4014
rect 6000 3392 6052 3398
rect 6000 3334 6052 3340
rect 5814 3224 5870 3233
rect 5724 3188 5776 3194
rect 5814 3159 5816 3168
rect 5724 3130 5776 3136
rect 5868 3159 5870 3168
rect 5816 3130 5868 3136
rect 5736 2446 5764 3130
rect 6012 3097 6040 3334
rect 5998 3088 6054 3097
rect 5998 3023 6054 3032
rect 5724 2440 5776 2446
rect 5724 2382 5776 2388
rect 5632 1896 5684 1902
rect 5632 1838 5684 1844
rect 5644 1222 5672 1838
rect 6012 1290 6040 3023
rect 6104 1358 6132 6054
rect 6276 5228 6328 5234
rect 6276 5170 6328 5176
rect 6184 5160 6236 5166
rect 6184 5102 6236 5108
rect 6196 4690 6224 5102
rect 6288 4690 6316 5170
rect 6184 4684 6236 4690
rect 6184 4626 6236 4632
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6380 3738 6408 7210
rect 6552 6724 6604 6730
rect 6552 6666 6604 6672
rect 6564 6322 6592 6666
rect 6656 6662 6684 7346
rect 6932 7206 6960 8298
rect 6736 7200 6788 7206
rect 6736 7142 6788 7148
rect 6920 7200 6972 7206
rect 6920 7142 6972 7148
rect 6748 6866 6776 7142
rect 6736 6860 6788 6866
rect 6736 6802 6788 6808
rect 6644 6656 6696 6662
rect 6644 6598 6696 6604
rect 6656 6458 6684 6598
rect 6644 6452 6696 6458
rect 6644 6394 6696 6400
rect 6748 6390 6776 6802
rect 6736 6384 6788 6390
rect 6736 6326 6788 6332
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6748 5710 6776 6326
rect 7024 6322 7052 8434
rect 7116 8090 7144 8842
rect 7208 8430 7236 8978
rect 7300 8566 7328 10202
rect 7564 10124 7616 10130
rect 7564 10066 7616 10072
rect 7472 9716 7524 9722
rect 7472 9658 7524 9664
rect 7484 9586 7512 9658
rect 7472 9580 7524 9586
rect 7472 9522 7524 9528
rect 7380 9376 7432 9382
rect 7380 9318 7432 9324
rect 7392 8906 7420 9318
rect 7484 8974 7512 9522
rect 7576 9518 7604 10066
rect 7944 9994 7972 10406
rect 7932 9988 7984 9994
rect 7932 9930 7984 9936
rect 8208 9818 8528 10854
rect 8576 10668 8628 10674
rect 8576 10610 8628 10616
rect 8588 10266 8616 10610
rect 8576 10260 8628 10266
rect 8576 10202 8628 10208
rect 8208 9766 8214 9818
rect 8266 9766 8278 9818
rect 8330 9766 8342 9818
rect 8394 9766 8406 9818
rect 8458 9766 8470 9818
rect 8522 9766 8528 9818
rect 7564 9512 7616 9518
rect 7564 9454 7616 9460
rect 7840 9512 7892 9518
rect 7840 9454 7892 9460
rect 7472 8968 7524 8974
rect 7472 8910 7524 8916
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7288 8560 7340 8566
rect 7288 8502 7340 8508
rect 7196 8424 7248 8430
rect 7196 8366 7248 8372
rect 7288 8288 7340 8294
rect 7288 8230 7340 8236
rect 7104 8084 7156 8090
rect 7104 8026 7156 8032
rect 7196 8084 7248 8090
rect 7196 8026 7248 8032
rect 7104 7880 7156 7886
rect 7102 7848 7104 7857
rect 7156 7848 7158 7857
rect 7102 7783 7158 7792
rect 7208 6322 7236 8026
rect 7300 8022 7328 8230
rect 7288 8016 7340 8022
rect 7288 7958 7340 7964
rect 7288 7540 7340 7546
rect 7392 7528 7420 8842
rect 7484 8090 7512 8910
rect 7852 8906 7880 9454
rect 8024 9104 8076 9110
rect 8024 9046 8076 9052
rect 8036 8906 8064 9046
rect 7840 8900 7892 8906
rect 7840 8842 7892 8848
rect 8024 8900 8076 8906
rect 8024 8842 8076 8848
rect 7748 8832 7800 8838
rect 7748 8774 7800 8780
rect 7760 8566 7788 8774
rect 7748 8560 7800 8566
rect 7748 8502 7800 8508
rect 7746 8120 7802 8129
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 7564 8084 7616 8090
rect 7746 8055 7802 8064
rect 7564 8026 7616 8032
rect 7340 7500 7420 7528
rect 7288 7482 7340 7488
rect 7576 6458 7604 8026
rect 7760 8022 7788 8055
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7852 7886 7880 8842
rect 7932 7948 7984 7954
rect 7932 7890 7984 7896
rect 7840 7880 7892 7886
rect 7944 7857 7972 7890
rect 7840 7822 7892 7828
rect 7930 7848 7986 7857
rect 7930 7783 7986 7792
rect 7656 7744 7708 7750
rect 7656 7686 7708 7692
rect 7668 7478 7696 7686
rect 7944 7546 7972 7783
rect 7932 7540 7984 7546
rect 7932 7482 7984 7488
rect 7656 7472 7708 7478
rect 7656 7414 7708 7420
rect 8036 7002 8064 8842
rect 8208 8730 8528 9766
rect 8680 9178 8708 11018
rect 8772 9382 8800 11222
rect 8956 10606 8984 12582
rect 9140 11830 9168 13126
rect 9128 11824 9180 11830
rect 9128 11766 9180 11772
rect 9324 10810 9352 13194
rect 9508 12918 9536 13670
rect 9784 12986 9812 14350
rect 9876 14346 9904 14962
rect 9968 14618 9996 17274
rect 10600 17264 10652 17270
rect 10600 17206 10652 17212
rect 10232 17196 10284 17202
rect 10232 17138 10284 17144
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10152 15026 10180 15846
rect 10244 15502 10272 17138
rect 10324 15972 10376 15978
rect 10324 15914 10376 15920
rect 10336 15502 10364 15914
rect 10612 15502 10640 17206
rect 10704 17134 10732 17614
rect 10692 17128 10744 17134
rect 10692 17070 10744 17076
rect 10232 15496 10284 15502
rect 10232 15438 10284 15444
rect 10324 15496 10376 15502
rect 10324 15438 10376 15444
rect 10600 15496 10652 15502
rect 10600 15438 10652 15444
rect 10244 15162 10272 15438
rect 10232 15156 10284 15162
rect 10232 15098 10284 15104
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 9956 14612 10008 14618
rect 9956 14554 10008 14560
rect 9864 14340 9916 14346
rect 9864 14282 9916 14288
rect 10336 13938 10364 15438
rect 10416 15360 10468 15366
rect 10416 15302 10468 15308
rect 10428 14958 10456 15302
rect 10612 15094 10640 15438
rect 10600 15088 10652 15094
rect 10600 15030 10652 15036
rect 10416 14952 10468 14958
rect 10416 14894 10468 14900
rect 10598 14920 10654 14929
rect 10428 14414 10456 14894
rect 10598 14855 10600 14864
rect 10652 14855 10654 14864
rect 10600 14826 10652 14832
rect 10508 14816 10560 14822
rect 10508 14758 10560 14764
rect 10416 14408 10468 14414
rect 10416 14350 10468 14356
rect 10520 13938 10548 14758
rect 10598 14512 10654 14521
rect 10598 14447 10654 14456
rect 10324 13932 10376 13938
rect 10324 13874 10376 13880
rect 10508 13932 10560 13938
rect 10508 13874 10560 13880
rect 10140 13728 10192 13734
rect 10140 13670 10192 13676
rect 9864 13320 9916 13326
rect 9864 13262 9916 13268
rect 9772 12980 9824 12986
rect 9772 12922 9824 12928
rect 9496 12912 9548 12918
rect 9496 12854 9548 12860
rect 9496 12776 9548 12782
rect 9496 12718 9548 12724
rect 9508 12442 9536 12718
rect 9496 12436 9548 12442
rect 9876 12434 9904 13262
rect 9876 12406 10088 12434
rect 9496 12378 9548 12384
rect 9772 12232 9824 12238
rect 9772 12174 9824 12180
rect 9956 12232 10008 12238
rect 9956 12174 10008 12180
rect 9496 12164 9548 12170
rect 9496 12106 9548 12112
rect 9508 11898 9536 12106
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9680 11620 9732 11626
rect 9680 11562 9732 11568
rect 9692 11150 9720 11562
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9404 11076 9456 11082
rect 9404 11018 9456 11024
rect 9128 10804 9180 10810
rect 9128 10746 9180 10752
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 8944 10600 8996 10606
rect 8944 10542 8996 10548
rect 8956 9654 8984 10542
rect 9036 10532 9088 10538
rect 9036 10474 9088 10480
rect 9048 9722 9076 10474
rect 9036 9716 9088 9722
rect 9036 9658 9088 9664
rect 8944 9648 8996 9654
rect 8944 9590 8996 9596
rect 8760 9376 8812 9382
rect 8760 9318 8812 9324
rect 8668 9172 8720 9178
rect 8668 9114 8720 9120
rect 8208 8678 8214 8730
rect 8266 8678 8278 8730
rect 8330 8678 8342 8730
rect 8394 8678 8406 8730
rect 8458 8678 8470 8730
rect 8522 8678 8528 8730
rect 8208 8518 8528 8678
rect 8208 8462 8220 8518
rect 8276 8462 8300 8518
rect 8356 8462 8380 8518
rect 8436 8462 8460 8518
rect 8516 8462 8528 8518
rect 8208 8438 8528 8462
rect 8208 8382 8220 8438
rect 8276 8382 8300 8438
rect 8356 8382 8380 8438
rect 8436 8382 8460 8438
rect 8516 8382 8528 8438
rect 8208 8358 8528 8382
rect 8208 8302 8220 8358
rect 8276 8302 8300 8358
rect 8356 8302 8380 8358
rect 8436 8302 8460 8358
rect 8516 8302 8528 8358
rect 8208 8278 8528 8302
rect 8208 8222 8220 8278
rect 8276 8222 8300 8278
rect 8356 8222 8380 8278
rect 8436 8222 8460 8278
rect 8516 8222 8528 8278
rect 8116 7880 8168 7886
rect 8116 7822 8168 7828
rect 8128 7546 8156 7822
rect 8208 7642 8528 8222
rect 8208 7590 8214 7642
rect 8266 7590 8278 7642
rect 8330 7590 8342 7642
rect 8394 7590 8406 7642
rect 8458 7590 8470 7642
rect 8522 7590 8528 7642
rect 8116 7540 8168 7546
rect 8116 7482 8168 7488
rect 8024 6996 8076 7002
rect 8024 6938 8076 6944
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7564 6452 7616 6458
rect 7564 6394 7616 6400
rect 7852 6390 7880 6734
rect 8116 6656 8168 6662
rect 8116 6598 8168 6604
rect 8128 6458 8156 6598
rect 8208 6554 8528 7590
rect 8680 7478 8708 9114
rect 8760 8832 8812 8838
rect 8760 8774 8812 8780
rect 8772 8566 8800 8774
rect 8760 8560 8812 8566
rect 8760 8502 8812 8508
rect 9048 7886 9076 9658
rect 9140 9654 9168 10746
rect 9220 9988 9272 9994
rect 9220 9930 9272 9936
rect 9312 9988 9364 9994
rect 9312 9930 9364 9936
rect 9128 9648 9180 9654
rect 9128 9590 9180 9596
rect 9232 8634 9260 9930
rect 9324 9178 9352 9930
rect 9312 9172 9364 9178
rect 9312 9114 9364 9120
rect 9416 8974 9444 11018
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9404 8968 9456 8974
rect 9404 8910 9456 8916
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9036 7880 9088 7886
rect 9036 7822 9088 7828
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8576 7200 8628 7206
rect 8576 7142 8628 7148
rect 8668 7200 8720 7206
rect 8668 7142 8720 7148
rect 8208 6502 8214 6554
rect 8266 6502 8278 6554
rect 8330 6502 8342 6554
rect 8394 6502 8406 6554
rect 8458 6502 8470 6554
rect 8522 6502 8528 6554
rect 8116 6452 8168 6458
rect 8116 6394 8168 6400
rect 7840 6384 7892 6390
rect 7840 6326 7892 6332
rect 7012 6316 7064 6322
rect 7196 6316 7248 6322
rect 7012 6258 7064 6264
rect 7116 6276 7196 6304
rect 6736 5704 6788 5710
rect 6736 5646 6788 5652
rect 6460 5636 6512 5642
rect 6460 5578 6512 5584
rect 6472 5302 6500 5578
rect 6460 5296 6512 5302
rect 6460 5238 6512 5244
rect 7012 5228 7064 5234
rect 7116 5216 7144 6276
rect 7196 6258 7248 6264
rect 7564 6112 7616 6118
rect 7564 6054 7616 6060
rect 7380 5568 7432 5574
rect 7380 5510 7432 5516
rect 7392 5370 7420 5510
rect 7288 5364 7340 5370
rect 7288 5306 7340 5312
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 7064 5188 7144 5216
rect 7012 5170 7064 5176
rect 6460 5024 6512 5030
rect 6460 4966 6512 4972
rect 7012 5024 7064 5030
rect 7012 4966 7064 4972
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6184 3460 6236 3466
rect 6184 3402 6236 3408
rect 6196 3194 6224 3402
rect 6274 3360 6330 3369
rect 6274 3295 6330 3304
rect 6184 3188 6236 3194
rect 6184 3130 6236 3136
rect 6288 3126 6316 3295
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6380 2854 6408 3674
rect 6368 2848 6420 2854
rect 6368 2790 6420 2796
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 6368 1352 6420 1358
rect 6368 1294 6420 1300
rect 6000 1284 6052 1290
rect 6000 1226 6052 1232
rect 5632 1216 5684 1222
rect 6380 1193 6408 1294
rect 5632 1158 5684 1164
rect 6366 1184 6422 1193
rect 6366 1119 6422 1128
rect 6472 882 6500 4966
rect 7024 4622 7052 4966
rect 7116 4622 7144 5188
rect 7300 4826 7328 5306
rect 7576 5234 7604 6054
rect 7852 5914 7880 6326
rect 7840 5908 7892 5914
rect 7840 5850 7892 5856
rect 8128 5710 8156 6394
rect 8116 5704 8168 5710
rect 8116 5646 8168 5652
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7852 5234 7880 5578
rect 8208 5466 8528 6502
rect 8588 6458 8616 7142
rect 8576 6452 8628 6458
rect 8576 6394 8628 6400
rect 8576 6112 8628 6118
rect 8576 6054 8628 6060
rect 8588 5846 8616 6054
rect 8576 5840 8628 5846
rect 8576 5782 8628 5788
rect 8208 5414 8214 5466
rect 8266 5414 8278 5466
rect 8330 5414 8342 5466
rect 8394 5414 8406 5466
rect 8458 5414 8470 5466
rect 8522 5414 8528 5466
rect 7932 5364 7984 5370
rect 7932 5306 7984 5312
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7840 5228 7892 5234
rect 7840 5170 7892 5176
rect 7380 5024 7432 5030
rect 7380 4966 7432 4972
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 7196 4684 7248 4690
rect 7196 4626 7248 4632
rect 7012 4616 7064 4622
rect 7012 4558 7064 4564
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6828 4480 6880 4486
rect 6828 4422 6880 4428
rect 6840 4214 6868 4422
rect 7116 4282 7144 4558
rect 7104 4276 7156 4282
rect 7104 4218 7156 4224
rect 6828 4208 6880 4214
rect 6828 4150 6880 4156
rect 7012 4072 7064 4078
rect 7012 4014 7064 4020
rect 6552 3936 6604 3942
rect 6552 3878 6604 3884
rect 6564 3194 6592 3878
rect 7024 3738 7052 4014
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7116 3602 7144 3878
rect 7208 3602 7236 4626
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 6736 3460 6788 3466
rect 6736 3402 6788 3408
rect 6748 3369 6776 3402
rect 6920 3392 6972 3398
rect 6734 3360 6790 3369
rect 6920 3334 6972 3340
rect 6734 3295 6790 3304
rect 6932 3233 6960 3334
rect 6918 3224 6974 3233
rect 6552 3188 6604 3194
rect 6918 3159 6974 3168
rect 6552 3130 6604 3136
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6552 2984 6604 2990
rect 6552 2926 6604 2932
rect 6564 2650 6592 2926
rect 6552 2644 6604 2650
rect 6552 2586 6604 2592
rect 6748 2514 6776 2994
rect 6736 2508 6788 2514
rect 6736 2450 6788 2456
rect 6644 2304 6696 2310
rect 6644 2246 6696 2252
rect 6656 1850 6684 2246
rect 6748 2038 6776 2450
rect 6828 2440 6880 2446
rect 6828 2382 6880 2388
rect 6736 2032 6788 2038
rect 6736 1974 6788 1980
rect 6656 1834 6776 1850
rect 6656 1828 6788 1834
rect 6656 1822 6736 1828
rect 6736 1770 6788 1776
rect 6840 1426 6868 2382
rect 6932 1578 6960 3159
rect 7012 2440 7064 2446
rect 7012 2382 7064 2388
rect 7024 1766 7052 2382
rect 7116 1902 7144 3538
rect 7300 3534 7328 4762
rect 7392 4690 7420 4966
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7380 4208 7432 4214
rect 7380 4150 7432 4156
rect 7392 3738 7420 4150
rect 7472 4072 7524 4078
rect 7472 4014 7524 4020
rect 7484 3942 7512 4014
rect 7472 3936 7524 3942
rect 7472 3878 7524 3884
rect 7470 3768 7526 3777
rect 7380 3732 7432 3738
rect 7470 3703 7526 3712
rect 7380 3674 7432 3680
rect 7288 3528 7340 3534
rect 7288 3470 7340 3476
rect 7288 3052 7340 3058
rect 7288 2994 7340 3000
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7104 1896 7156 1902
rect 7104 1838 7156 1844
rect 7012 1760 7064 1766
rect 7012 1702 7064 1708
rect 7104 1760 7156 1766
rect 7104 1702 7156 1708
rect 7116 1578 7144 1702
rect 6932 1550 7144 1578
rect 7208 1494 7236 2586
rect 7300 1562 7328 2994
rect 7484 2922 7512 3703
rect 7576 3466 7604 5170
rect 7656 4616 7708 4622
rect 7656 4558 7708 4564
rect 7668 4078 7696 4558
rect 7656 4072 7708 4078
rect 7656 4014 7708 4020
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7564 3460 7616 3466
rect 7564 3402 7616 3408
rect 7472 2916 7524 2922
rect 7472 2858 7524 2864
rect 7564 2848 7616 2854
rect 7564 2790 7616 2796
rect 7576 2038 7604 2790
rect 7668 2446 7696 3606
rect 7944 3534 7972 5306
rect 8116 5160 8168 5166
rect 8116 5102 8168 5108
rect 8128 3534 8156 5102
rect 8208 4378 8528 5414
rect 8680 5234 8708 7142
rect 8772 6662 8800 7346
rect 9232 7342 9260 8570
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9496 7744 9548 7750
rect 9496 7686 9548 7692
rect 9508 7478 9536 7686
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9600 7342 9628 7822
rect 9220 7336 9272 7342
rect 9220 7278 9272 7284
rect 9588 7336 9640 7342
rect 9588 7278 9640 7284
rect 8852 6724 8904 6730
rect 8852 6666 8904 6672
rect 8760 6656 8812 6662
rect 8760 6598 8812 6604
rect 8668 5228 8720 5234
rect 8668 5170 8720 5176
rect 8772 4826 8800 6598
rect 8864 5846 8892 6666
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8852 5840 8904 5846
rect 8852 5782 8904 5788
rect 8956 5710 8984 6394
rect 9232 6390 9260 7278
rect 9692 6934 9720 10610
rect 9784 10538 9812 12174
rect 9968 11830 9996 12174
rect 9956 11824 10008 11830
rect 9956 11766 10008 11772
rect 9968 11218 9996 11766
rect 9956 11212 10008 11218
rect 9956 11154 10008 11160
rect 9864 11144 9916 11150
rect 10060 11098 10088 12406
rect 10152 12170 10180 13670
rect 10336 13326 10364 13874
rect 10612 13870 10640 14447
rect 10600 13864 10652 13870
rect 10600 13806 10652 13812
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10336 12918 10364 13262
rect 10612 12986 10640 13806
rect 10704 13258 10732 17070
rect 10888 15502 10916 18362
rect 11520 18216 11572 18222
rect 11520 18158 11572 18164
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 11164 17270 11192 18022
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11532 17184 11560 18158
rect 11624 17746 11652 19200
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 13176 18624 13228 18630
rect 13176 18566 13228 18572
rect 12072 18148 12124 18154
rect 12072 18090 12124 18096
rect 11612 17740 11664 17746
rect 11612 17682 11664 17688
rect 12084 17270 12112 18090
rect 12208 17978 12528 18544
rect 13188 18290 13216 18566
rect 13372 18426 13400 18634
rect 13360 18420 13412 18426
rect 13360 18362 13412 18368
rect 13832 18290 13860 19246
rect 14186 19200 14242 20000
rect 16762 19200 16818 20000
rect 19338 19200 19394 20000
rect 21914 19200 21970 20000
rect 24400 19304 24452 19310
rect 24400 19246 24452 19252
rect 14200 18426 14228 19200
rect 16208 18522 16528 18544
rect 16208 18470 16214 18522
rect 16266 18470 16278 18522
rect 16330 18470 16342 18522
rect 16394 18470 16406 18522
rect 16458 18470 16470 18522
rect 16522 18470 16528 18522
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 12716 18284 12768 18290
rect 12716 18226 12768 18232
rect 13176 18284 13228 18290
rect 13176 18226 13228 18232
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 12208 17926 12214 17978
rect 12266 17926 12278 17978
rect 12330 17926 12342 17978
rect 12394 17926 12406 17978
rect 12458 17926 12470 17978
rect 12522 17926 12528 17978
rect 12072 17264 12124 17270
rect 12072 17206 12124 17212
rect 11612 17196 11664 17202
rect 11532 17156 11612 17184
rect 11612 17138 11664 17144
rect 11624 17066 11652 17138
rect 11612 17060 11664 17066
rect 11612 17002 11664 17008
rect 12208 16890 12528 17926
rect 12728 17678 12756 18226
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 17270 12756 17614
rect 12808 17604 12860 17610
rect 12808 17546 12860 17552
rect 13544 17604 13596 17610
rect 13544 17546 13596 17552
rect 12716 17264 12768 17270
rect 12716 17206 12768 17212
rect 12716 17128 12768 17134
rect 12820 17116 12848 17546
rect 13084 17196 13136 17202
rect 13084 17138 13136 17144
rect 12768 17088 12848 17116
rect 12716 17070 12768 17076
rect 12208 16838 12214 16890
rect 12266 16838 12278 16890
rect 12330 16838 12342 16890
rect 12394 16838 12406 16890
rect 12458 16838 12470 16890
rect 12522 16838 12528 16890
rect 11060 16720 11112 16726
rect 11060 16662 11112 16668
rect 11072 16590 11100 16662
rect 11060 16584 11112 16590
rect 11060 16526 11112 16532
rect 11072 16250 11100 16526
rect 11060 16244 11112 16250
rect 11060 16186 11112 16192
rect 11152 16176 11204 16182
rect 11152 16118 11204 16124
rect 10876 15496 10928 15502
rect 10876 15438 10928 15444
rect 10876 15360 10928 15366
rect 10876 15302 10928 15308
rect 10784 14816 10836 14822
rect 10784 14758 10836 14764
rect 10796 14414 10824 14758
rect 10784 14408 10836 14414
rect 10782 14376 10784 14385
rect 10836 14376 10838 14385
rect 10782 14311 10838 14320
rect 10784 13932 10836 13938
rect 10784 13874 10836 13880
rect 10796 13394 10824 13874
rect 10888 13462 10916 15302
rect 11164 14890 11192 16118
rect 11612 16108 11664 16114
rect 11612 16050 11664 16056
rect 11624 15570 11652 16050
rect 11980 15904 12032 15910
rect 11980 15846 12032 15852
rect 11992 15570 12020 15846
rect 12208 15802 12528 16838
rect 12820 16590 12848 17088
rect 13096 16658 13124 17138
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13372 16998 13400 17070
rect 13556 17066 13584 17546
rect 13544 17060 13596 17066
rect 13544 17002 13596 17008
rect 13360 16992 13412 16998
rect 13360 16934 13412 16940
rect 13556 16726 13584 17002
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12624 16516 12676 16522
rect 12624 16458 12676 16464
rect 12636 16114 12664 16458
rect 12624 16108 12676 16114
rect 12624 16050 12676 16056
rect 12900 15972 12952 15978
rect 12900 15914 12952 15920
rect 12208 15750 12214 15802
rect 12266 15750 12278 15802
rect 12330 15750 12342 15802
rect 12394 15750 12406 15802
rect 12458 15750 12470 15802
rect 12522 15750 12528 15802
rect 11612 15564 11664 15570
rect 11612 15506 11664 15512
rect 11980 15564 12032 15570
rect 11980 15506 12032 15512
rect 11624 15026 11652 15506
rect 11704 15088 11756 15094
rect 11704 15030 11756 15036
rect 11336 15020 11388 15026
rect 11336 14962 11388 14968
rect 11612 15020 11664 15026
rect 11612 14962 11664 14968
rect 11152 14884 11204 14890
rect 11152 14826 11204 14832
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 10980 14550 11008 14758
rect 10968 14544 11020 14550
rect 10968 14486 11020 14492
rect 11164 14396 11192 14826
rect 11244 14408 11296 14414
rect 11164 14368 11244 14396
rect 10968 14068 11020 14074
rect 10968 14010 11020 14016
rect 10980 13870 11008 14010
rect 11060 14000 11112 14006
rect 11060 13942 11112 13948
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10966 13560 11022 13569
rect 10966 13495 11022 13504
rect 10876 13456 10928 13462
rect 10876 13398 10928 13404
rect 10784 13388 10836 13394
rect 10784 13330 10836 13336
rect 10692 13252 10744 13258
rect 10692 13194 10744 13200
rect 10980 13190 11008 13495
rect 10968 13184 11020 13190
rect 10968 13126 11020 13132
rect 10600 12980 10652 12986
rect 10600 12922 10652 12928
rect 10324 12912 10376 12918
rect 10324 12854 10376 12860
rect 10980 12306 11008 13126
rect 10968 12300 11020 12306
rect 10968 12242 11020 12248
rect 10140 12164 10192 12170
rect 10140 12106 10192 12112
rect 10416 12164 10468 12170
rect 10416 12106 10468 12112
rect 10600 12164 10652 12170
rect 10600 12106 10652 12112
rect 10232 12096 10284 12102
rect 10152 12044 10232 12050
rect 10152 12038 10284 12044
rect 10324 12096 10376 12102
rect 10324 12038 10376 12044
rect 10152 12022 10272 12038
rect 10152 11150 10180 12022
rect 10336 11762 10364 12038
rect 10324 11756 10376 11762
rect 10324 11698 10376 11704
rect 10428 11218 10456 12106
rect 10612 11898 10640 12106
rect 10980 12102 11008 12242
rect 11072 12238 11100 13942
rect 11164 13802 11192 14368
rect 11244 14350 11296 14356
rect 11348 14346 11376 14962
rect 11716 14464 11744 15030
rect 11796 15020 11848 15026
rect 11796 14962 11848 14968
rect 11980 15020 12032 15026
rect 11980 14962 12032 14968
rect 11808 14618 11836 14962
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11624 14436 11744 14464
rect 11428 14408 11480 14414
rect 11428 14350 11480 14356
rect 11336 14340 11388 14346
rect 11336 14282 11388 14288
rect 11244 14272 11296 14278
rect 11244 14214 11296 14220
rect 11152 13796 11204 13802
rect 11152 13738 11204 13744
rect 11150 13424 11206 13433
rect 11150 13359 11206 13368
rect 11164 13326 11192 13359
rect 11152 13320 11204 13326
rect 11152 13262 11204 13268
rect 11256 12356 11284 14214
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11348 13308 11376 13738
rect 11440 13433 11468 14350
rect 11624 13938 11652 14436
rect 11796 14408 11848 14414
rect 11702 14376 11758 14385
rect 11796 14350 11848 14356
rect 11702 14311 11758 14320
rect 11612 13932 11664 13938
rect 11612 13874 11664 13880
rect 11426 13424 11482 13433
rect 11426 13359 11482 13368
rect 11348 13280 11468 13308
rect 11336 12776 11388 12782
rect 11336 12718 11388 12724
rect 11164 12328 11284 12356
rect 11060 12232 11112 12238
rect 11060 12174 11112 12180
rect 10968 12096 11020 12102
rect 10968 12038 11020 12044
rect 10600 11892 10652 11898
rect 10600 11834 10652 11840
rect 10416 11212 10468 11218
rect 10416 11154 10468 11160
rect 9864 11086 9916 11092
rect 9876 10742 9904 11086
rect 9968 11070 10088 11098
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9864 10736 9916 10742
rect 9864 10678 9916 10684
rect 9772 10532 9824 10538
rect 9772 10474 9824 10480
rect 9772 9988 9824 9994
rect 9772 9930 9824 9936
rect 9784 9450 9812 9930
rect 9864 9580 9916 9586
rect 9864 9522 9916 9528
rect 9772 9444 9824 9450
rect 9772 9386 9824 9392
rect 9876 8838 9904 9522
rect 9864 8832 9916 8838
rect 9864 8774 9916 8780
rect 9864 7336 9916 7342
rect 9784 7296 9864 7324
rect 9680 6928 9732 6934
rect 9600 6876 9680 6882
rect 9600 6870 9732 6876
rect 9600 6854 9720 6870
rect 9312 6724 9364 6730
rect 9312 6666 9364 6672
rect 9220 6384 9272 6390
rect 9220 6326 9272 6332
rect 9036 6112 9088 6118
rect 9036 6054 9088 6060
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8760 4820 8812 4826
rect 8760 4762 8812 4768
rect 8668 4616 8720 4622
rect 8668 4558 8720 4564
rect 8208 4326 8214 4378
rect 8266 4326 8278 4378
rect 8330 4326 8342 4378
rect 8394 4326 8406 4378
rect 8458 4326 8470 4378
rect 8522 4326 8528 4378
rect 7932 3528 7984 3534
rect 7932 3470 7984 3476
rect 8116 3528 8168 3534
rect 8116 3470 8168 3476
rect 8024 3392 8076 3398
rect 8024 3334 8076 3340
rect 8036 3058 8064 3334
rect 8208 3290 8528 4326
rect 8680 3942 8708 4558
rect 8760 4004 8812 4010
rect 8760 3946 8812 3952
rect 8668 3936 8720 3942
rect 8668 3878 8720 3884
rect 8208 3238 8214 3290
rect 8266 3238 8278 3290
rect 8330 3238 8342 3290
rect 8394 3238 8406 3290
rect 8458 3238 8470 3290
rect 8522 3238 8528 3290
rect 8024 3052 8076 3058
rect 8024 2994 8076 3000
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7760 2582 7788 2790
rect 8114 2680 8170 2689
rect 8114 2615 8170 2624
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7838 2544 7894 2553
rect 8128 2514 8156 2615
rect 7838 2479 7840 2488
rect 7892 2479 7894 2488
rect 8116 2508 8168 2514
rect 7840 2450 7892 2456
rect 8116 2450 8168 2456
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7932 2440 7984 2446
rect 7932 2382 7984 2388
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 7564 2032 7616 2038
rect 7564 1974 7616 1980
rect 7380 1964 7432 1970
rect 7380 1906 7432 1912
rect 7288 1556 7340 1562
rect 7288 1498 7340 1504
rect 7392 1494 7420 1906
rect 7472 1828 7524 1834
rect 7472 1770 7524 1776
rect 7484 1562 7512 1770
rect 7472 1556 7524 1562
rect 7472 1498 7524 1504
rect 7840 1556 7892 1562
rect 7840 1498 7892 1504
rect 7196 1488 7248 1494
rect 7196 1430 7248 1436
rect 7380 1488 7432 1494
rect 7380 1430 7432 1436
rect 6828 1420 6880 1426
rect 6828 1362 6880 1368
rect 7852 1358 7880 1498
rect 7944 1426 7972 2382
rect 8036 1465 8064 2382
rect 8116 2372 8168 2378
rect 8116 2314 8168 2320
rect 8128 1902 8156 2314
rect 8208 2202 8528 3238
rect 8576 2984 8628 2990
rect 8576 2926 8628 2932
rect 8588 2446 8616 2926
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8208 2150 8214 2202
rect 8266 2150 8278 2202
rect 8330 2150 8342 2202
rect 8394 2150 8406 2202
rect 8458 2150 8470 2202
rect 8522 2150 8528 2202
rect 8116 1896 8168 1902
rect 8116 1838 8168 1844
rect 8022 1456 8078 1465
rect 7932 1420 7984 1426
rect 8022 1391 8078 1400
rect 7932 1362 7984 1368
rect 7840 1352 7892 1358
rect 7840 1294 7892 1300
rect 6644 1216 6696 1222
rect 6644 1158 6696 1164
rect 6656 950 6684 1158
rect 8208 1114 8528 2150
rect 8680 1562 8708 3878
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 8772 1290 8800 3946
rect 9048 3777 9076 6054
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 9140 4690 9168 5102
rect 9128 4684 9180 4690
rect 9128 4626 9180 4632
rect 9034 3768 9090 3777
rect 9034 3703 9090 3712
rect 9232 3466 9260 6326
rect 9324 6254 9352 6666
rect 9404 6452 9456 6458
rect 9404 6394 9456 6400
rect 9416 6322 9444 6394
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5914 9352 6190
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9600 5794 9628 6854
rect 9680 6792 9732 6798
rect 9680 6734 9732 6740
rect 9692 6322 9720 6734
rect 9680 6316 9732 6322
rect 9680 6258 9732 6264
rect 9416 5766 9628 5794
rect 9312 4140 9364 4146
rect 9312 4082 9364 4088
rect 9220 3460 9272 3466
rect 9220 3402 9272 3408
rect 9324 2922 9352 4082
rect 9416 3398 9444 5766
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9508 5302 9536 5646
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9496 5296 9548 5302
rect 9496 5238 9548 5244
rect 9600 4214 9628 5510
rect 9692 5166 9720 6258
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9784 4729 9812 7296
rect 9864 7278 9916 7284
rect 9968 5114 9996 11070
rect 10048 11008 10100 11014
rect 10048 10950 10100 10956
rect 10060 10810 10088 10950
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10152 10690 10180 11086
rect 10612 11082 10640 11834
rect 10692 11824 10744 11830
rect 10692 11766 10744 11772
rect 10704 11234 10732 11766
rect 11164 11744 11192 12328
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11072 11716 11192 11744
rect 10784 11688 10836 11694
rect 10784 11630 10836 11636
rect 10796 11354 10824 11630
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10704 11206 10824 11234
rect 10796 11150 10824 11206
rect 10784 11144 10836 11150
rect 10784 11086 10836 11092
rect 10600 11076 10652 11082
rect 10600 11018 10652 11024
rect 10324 11008 10376 11014
rect 10324 10950 10376 10956
rect 10060 10662 10180 10690
rect 10060 8294 10088 10662
rect 10336 10606 10364 10950
rect 10324 10600 10376 10606
rect 10324 10542 10376 10548
rect 10336 10130 10364 10542
rect 10324 10124 10376 10130
rect 10152 10084 10324 10112
rect 10048 8288 10100 8294
rect 10048 8230 10100 8236
rect 9876 5086 9996 5114
rect 9770 4720 9826 4729
rect 9770 4655 9826 4664
rect 9680 4616 9732 4622
rect 9680 4558 9732 4564
rect 9692 4282 9720 4558
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 9588 4208 9640 4214
rect 9588 4150 9640 4156
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9680 4072 9732 4078
rect 9678 4040 9680 4049
rect 9732 4040 9734 4049
rect 9678 3975 9734 3984
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9692 3602 9720 3878
rect 9784 3618 9812 4082
rect 9876 3738 9904 5086
rect 9954 4720 10010 4729
rect 9954 4655 10010 4664
rect 9968 4554 9996 4655
rect 10060 4554 10088 8230
rect 9956 4548 10008 4554
rect 9956 4490 10008 4496
rect 10048 4548 10100 4554
rect 10048 4490 10100 4496
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9968 3738 9996 4082
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 9956 3732 10008 3738
rect 9956 3674 10008 3680
rect 9680 3596 9732 3602
rect 9784 3590 10088 3618
rect 9680 3538 9732 3544
rect 9404 3392 9456 3398
rect 9404 3334 9456 3340
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 9588 2984 9640 2990
rect 9588 2926 9640 2932
rect 9312 2916 9364 2922
rect 9312 2858 9364 2864
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9048 2582 9076 2790
rect 9036 2576 9088 2582
rect 8850 2544 8906 2553
rect 9036 2518 9088 2524
rect 8850 2479 8852 2488
rect 8904 2479 8906 2488
rect 8852 2450 8904 2456
rect 9036 2304 9088 2310
rect 9036 2246 9088 2252
rect 9048 2106 9076 2246
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 9600 1970 9628 2926
rect 9692 2774 9720 2994
rect 9956 2848 10008 2854
rect 9956 2790 10008 2796
rect 9692 2746 9812 2774
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 9692 2038 9720 2246
rect 9680 2032 9732 2038
rect 9680 1974 9732 1980
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9508 1465 9536 1498
rect 9494 1456 9550 1465
rect 9494 1391 9550 1400
rect 9600 1358 9628 1906
rect 9680 1896 9732 1902
rect 9680 1838 9732 1844
rect 9692 1766 9720 1838
rect 9680 1760 9732 1766
rect 9680 1702 9732 1708
rect 9588 1352 9640 1358
rect 9588 1294 9640 1300
rect 8576 1284 8628 1290
rect 8576 1226 8628 1232
rect 8760 1284 8812 1290
rect 8760 1226 8812 1232
rect 8208 1062 8214 1114
rect 8266 1062 8278 1114
rect 8330 1062 8342 1114
rect 8394 1062 8406 1114
rect 8458 1062 8470 1114
rect 8522 1062 8528 1114
rect 8208 1040 8528 1062
rect 6644 944 6696 950
rect 6644 886 6696 892
rect 8588 882 8616 1226
rect 6460 876 6512 882
rect 6460 818 6512 824
rect 7564 876 7616 882
rect 8576 876 8628 882
rect 7616 836 7696 864
rect 7564 818 7616 824
rect 7668 800 7696 836
rect 8576 818 8628 824
rect 9784 800 9812 2746
rect 9862 2544 9918 2553
rect 9862 2479 9864 2488
rect 9916 2479 9918 2488
rect 9864 2450 9916 2456
rect 9968 1766 9996 2790
rect 10060 2281 10088 3590
rect 10046 2272 10102 2281
rect 10046 2207 10102 2216
rect 10060 1970 10088 2207
rect 10152 2106 10180 10084
rect 10324 10066 10376 10072
rect 10232 9920 10284 9926
rect 10232 9862 10284 9868
rect 10244 9722 10272 9862
rect 10232 9716 10284 9722
rect 10232 9658 10284 9664
rect 10244 8566 10272 9658
rect 10324 9580 10376 9586
rect 10324 9522 10376 9528
rect 10336 8906 10364 9522
rect 10416 9512 10468 9518
rect 10416 9454 10468 9460
rect 10428 8906 10456 9454
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9178 10548 9318
rect 10508 9172 10560 9178
rect 10508 9114 10560 9120
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10508 8900 10560 8906
rect 10508 8842 10560 8848
rect 10336 8566 10364 8842
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10324 8560 10376 8566
rect 10324 8502 10376 8508
rect 10428 8498 10456 8842
rect 10520 8498 10548 8842
rect 10796 8498 10824 11086
rect 10876 10804 10928 10810
rect 10876 10746 10928 10752
rect 10888 10130 10916 10746
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 10124 10928 10130
rect 10876 10066 10928 10072
rect 10980 9994 11008 10678
rect 10968 9988 11020 9994
rect 10968 9930 11020 9936
rect 11072 9674 11100 11716
rect 11152 11620 11204 11626
rect 11152 11562 11204 11568
rect 11164 11082 11192 11562
rect 11152 11076 11204 11082
rect 11152 11018 11204 11024
rect 11072 9646 11192 9674
rect 10876 9580 10928 9586
rect 10876 9522 10928 9528
rect 10888 8974 10916 9522
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 11060 8968 11112 8974
rect 11060 8910 11112 8916
rect 10888 8634 10916 8910
rect 10876 8628 10928 8634
rect 10876 8570 10928 8576
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 10520 8090 10548 8434
rect 11072 8430 11100 8910
rect 11060 8424 11112 8430
rect 11060 8366 11112 8372
rect 10508 8084 10560 8090
rect 10508 8026 10560 8032
rect 11060 8084 11112 8090
rect 11060 8026 11112 8032
rect 11072 7886 11100 8026
rect 11164 8022 11192 9646
rect 11256 9518 11284 12174
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11256 9042 11284 9454
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 11152 8016 11204 8022
rect 11152 7958 11204 7964
rect 11348 7954 11376 12718
rect 11440 12306 11468 13280
rect 11716 13258 11744 14311
rect 11808 13920 11836 14350
rect 11900 14090 11928 14486
rect 11992 14278 12020 14962
rect 12208 14714 12528 15750
rect 12912 15502 12940 15914
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 13096 15162 13124 16594
rect 13832 16250 13860 18226
rect 14556 18216 14608 18222
rect 14476 18176 14556 18204
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 14280 18148 14332 18154
rect 14280 18090 14332 18096
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13924 16114 13952 18090
rect 14292 17202 14320 18090
rect 14476 17678 14504 18176
rect 14556 18158 14608 18164
rect 16120 18216 16172 18222
rect 16120 18158 16172 18164
rect 15292 18148 15344 18154
rect 15292 18090 15344 18096
rect 15304 17814 15332 18090
rect 15292 17808 15344 17814
rect 15292 17750 15344 17756
rect 16132 17678 16160 18158
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 16120 17672 16172 17678
rect 16120 17614 16172 17620
rect 14372 17264 14424 17270
rect 14372 17206 14424 17212
rect 14280 17196 14332 17202
rect 14280 17138 14332 17144
rect 14384 16590 14412 17206
rect 14372 16584 14424 16590
rect 14372 16526 14424 16532
rect 13268 16108 13320 16114
rect 13268 16050 13320 16056
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 13912 16108 13964 16114
rect 13912 16050 13964 16056
rect 13084 15156 13136 15162
rect 13084 15098 13136 15104
rect 13280 15026 13308 16050
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13372 15026 13400 15982
rect 13740 15094 13768 16050
rect 13820 15632 13872 15638
rect 13820 15574 13872 15580
rect 13728 15088 13780 15094
rect 13728 15030 13780 15036
rect 13832 15026 13860 15574
rect 12716 15020 12768 15026
rect 12716 14962 12768 14968
rect 12808 15020 12860 15026
rect 12808 14962 12860 14968
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13820 15020 13872 15026
rect 13820 14962 13872 14968
rect 12208 14662 12214 14714
rect 12266 14662 12278 14714
rect 12330 14662 12342 14714
rect 12394 14662 12406 14714
rect 12458 14662 12470 14714
rect 12522 14662 12528 14714
rect 12072 14544 12124 14550
rect 12070 14512 12072 14521
rect 12124 14512 12126 14521
rect 12070 14447 12126 14456
rect 12072 14408 12124 14414
rect 12072 14350 12124 14356
rect 11980 14272 12032 14278
rect 11980 14214 12032 14220
rect 11900 14062 12020 14090
rect 12084 14074 12112 14350
rect 11888 13932 11940 13938
rect 11808 13892 11888 13920
rect 11888 13874 11940 13880
rect 11900 13841 11928 13874
rect 11886 13832 11942 13841
rect 11992 13802 12020 14062
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12084 13938 12112 14010
rect 12072 13932 12124 13938
rect 12072 13874 12124 13880
rect 11886 13767 11942 13776
rect 11980 13796 12032 13802
rect 11980 13738 12032 13744
rect 11796 13728 11848 13734
rect 11796 13670 11848 13676
rect 11888 13728 11940 13734
rect 11888 13670 11940 13676
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11520 13184 11572 13190
rect 11520 13126 11572 13132
rect 11428 12300 11480 12306
rect 11428 12242 11480 12248
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11440 11626 11468 11698
rect 11428 11620 11480 11626
rect 11428 11562 11480 11568
rect 11440 11150 11468 11562
rect 11428 11144 11480 11150
rect 11428 11086 11480 11092
rect 11532 9586 11560 13126
rect 11716 12986 11744 13194
rect 11704 12980 11756 12986
rect 11704 12922 11756 12928
rect 11612 12844 11664 12850
rect 11612 12786 11664 12792
rect 11704 12844 11756 12850
rect 11704 12786 11756 12792
rect 11624 11218 11652 12786
rect 11716 11898 11744 12786
rect 11808 12714 11836 13670
rect 11900 12986 11928 13670
rect 12208 13626 12528 14662
rect 12624 13864 12676 13870
rect 12624 13806 12676 13812
rect 12208 13574 12214 13626
rect 12266 13574 12278 13626
rect 12330 13574 12342 13626
rect 12394 13574 12406 13626
rect 12458 13574 12470 13626
rect 12522 13574 12528 13626
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11888 12980 11940 12986
rect 11888 12922 11940 12928
rect 11992 12918 12020 13466
rect 12072 13184 12124 13190
rect 12072 13126 12124 13132
rect 12084 12986 12112 13126
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 11980 12912 12032 12918
rect 11980 12854 12032 12860
rect 11888 12844 11940 12850
rect 11888 12786 11940 12792
rect 12072 12844 12124 12850
rect 12072 12786 12124 12792
rect 11796 12708 11848 12714
rect 11796 12650 11848 12656
rect 11900 12238 11928 12786
rect 11980 12436 12032 12442
rect 11980 12378 12032 12384
rect 11888 12232 11940 12238
rect 11888 12174 11940 12180
rect 11704 11892 11756 11898
rect 11704 11834 11756 11840
rect 11716 11286 11744 11834
rect 11900 11694 11928 12174
rect 11796 11688 11848 11694
rect 11796 11630 11848 11636
rect 11888 11688 11940 11694
rect 11888 11630 11940 11636
rect 11704 11280 11756 11286
rect 11704 11222 11756 11228
rect 11612 11212 11664 11218
rect 11612 11154 11664 11160
rect 11808 11098 11836 11630
rect 11992 11558 12020 12378
rect 12084 12238 12112 12786
rect 12208 12538 12528 13574
rect 12636 13326 12664 13806
rect 12624 13320 12676 13326
rect 12624 13262 12676 13268
rect 12636 12782 12664 13262
rect 12624 12776 12676 12782
rect 12624 12718 12676 12724
rect 12208 12486 12214 12538
rect 12266 12518 12278 12538
rect 12330 12518 12342 12538
rect 12394 12518 12406 12538
rect 12458 12518 12470 12538
rect 12276 12486 12278 12518
rect 12458 12486 12460 12518
rect 12522 12486 12528 12538
rect 12208 12462 12220 12486
rect 12276 12462 12300 12486
rect 12356 12462 12380 12486
rect 12436 12462 12460 12486
rect 12516 12462 12528 12486
rect 12208 12438 12528 12462
rect 12208 12382 12220 12438
rect 12276 12382 12300 12438
rect 12356 12382 12380 12438
rect 12436 12382 12460 12438
rect 12516 12382 12528 12438
rect 12208 12358 12528 12382
rect 12208 12302 12220 12358
rect 12276 12302 12300 12358
rect 12356 12302 12380 12358
rect 12436 12302 12460 12358
rect 12516 12302 12528 12358
rect 12208 12278 12528 12302
rect 12072 12232 12124 12238
rect 12072 12174 12124 12180
rect 12208 12222 12220 12278
rect 12276 12222 12300 12278
rect 12356 12222 12380 12278
rect 12436 12222 12460 12278
rect 12516 12222 12528 12278
rect 12072 12096 12124 12102
rect 12072 12038 12124 12044
rect 12084 11762 12112 12038
rect 12072 11756 12124 11762
rect 12072 11698 12124 11704
rect 11980 11552 12032 11558
rect 11980 11494 12032 11500
rect 12208 11450 12528 12222
rect 12624 12232 12676 12238
rect 12624 12174 12676 12180
rect 12208 11398 12214 11450
rect 12266 11398 12278 11450
rect 12330 11398 12342 11450
rect 12394 11398 12406 11450
rect 12458 11398 12470 11450
rect 12522 11398 12528 11450
rect 11888 11144 11940 11150
rect 11808 11092 11888 11098
rect 11808 11086 11940 11092
rect 11808 11070 11928 11086
rect 11808 10742 11836 11070
rect 11888 11008 11940 11014
rect 11888 10950 11940 10956
rect 11796 10736 11848 10742
rect 11796 10678 11848 10684
rect 11900 10606 11928 10950
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 11900 8498 11928 10542
rect 12208 10362 12528 11398
rect 12636 11082 12664 12174
rect 12624 11076 12676 11082
rect 12624 11018 12676 11024
rect 12728 10826 12756 14962
rect 12820 14618 12848 14962
rect 13280 14618 13308 14962
rect 12808 14612 12860 14618
rect 12808 14554 12860 14560
rect 13268 14612 13320 14618
rect 13268 14554 13320 14560
rect 12900 14544 12952 14550
rect 12900 14486 12952 14492
rect 12912 14414 12940 14486
rect 13280 14414 13308 14554
rect 12900 14408 12952 14414
rect 12900 14350 12952 14356
rect 13268 14408 13320 14414
rect 13268 14350 13320 14356
rect 12992 14272 13044 14278
rect 12992 14214 13044 14220
rect 12808 13932 12860 13938
rect 12808 13874 12860 13880
rect 12820 12238 12848 13874
rect 13004 13870 13032 14214
rect 13280 14090 13308 14350
rect 13372 14278 13400 14962
rect 13544 14544 13596 14550
rect 13544 14486 13596 14492
rect 13360 14272 13412 14278
rect 13360 14214 13412 14220
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13280 14074 13400 14090
rect 13280 14068 13412 14074
rect 13280 14062 13360 14068
rect 13360 14010 13412 14016
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 12992 13864 13044 13870
rect 12992 13806 13044 13812
rect 13176 13388 13228 13394
rect 13176 13330 13228 13336
rect 12900 13320 12952 13326
rect 12900 13262 12952 13268
rect 12912 12306 12940 13262
rect 12992 13252 13044 13258
rect 12992 13194 13044 13200
rect 13004 12850 13032 13194
rect 12992 12844 13044 12850
rect 12992 12786 13044 12792
rect 13188 12434 13216 13330
rect 13280 12850 13308 13874
rect 13464 13258 13492 14214
rect 13452 13252 13504 13258
rect 13452 13194 13504 13200
rect 13556 13138 13584 14486
rect 14096 14340 14148 14346
rect 14096 14282 14148 14288
rect 13912 14272 13964 14278
rect 13912 14214 13964 14220
rect 13924 13938 13952 14214
rect 14108 14074 14136 14282
rect 14096 14068 14148 14074
rect 14096 14010 14148 14016
rect 14108 13938 14136 14010
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14096 13932 14148 13938
rect 14096 13874 14148 13880
rect 13820 13728 13872 13734
rect 13820 13670 13872 13676
rect 13634 13424 13690 13433
rect 13634 13359 13690 13368
rect 13648 13326 13676 13359
rect 13636 13320 13688 13326
rect 13636 13262 13688 13268
rect 13464 13110 13584 13138
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13188 12406 13400 12434
rect 12900 12300 12952 12306
rect 12900 12242 12952 12248
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 13268 12164 13320 12170
rect 13268 12106 13320 12112
rect 12808 12096 12860 12102
rect 12808 12038 12860 12044
rect 12820 11626 12848 12038
rect 13176 11756 13228 11762
rect 13176 11698 13228 11704
rect 12808 11620 12860 11626
rect 12808 11562 12860 11568
rect 13188 11218 13216 11698
rect 13280 11354 13308 12106
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 13372 11098 13400 12406
rect 13464 12238 13492 13110
rect 13452 12232 13504 12238
rect 13452 12174 13504 12180
rect 13544 12232 13596 12238
rect 13544 12174 13596 12180
rect 13452 11688 13504 11694
rect 13452 11630 13504 11636
rect 13464 11218 13492 11630
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13372 11070 13492 11098
rect 12728 10798 13124 10826
rect 12900 10736 12952 10742
rect 12900 10678 12952 10684
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12208 10310 12214 10362
rect 12266 10310 12278 10362
rect 12330 10310 12342 10362
rect 12394 10310 12406 10362
rect 12458 10310 12470 10362
rect 12522 10310 12528 10362
rect 12072 9580 12124 9586
rect 12072 9522 12124 9528
rect 12084 8974 12112 9522
rect 12208 9274 12528 10310
rect 12636 10266 12664 10610
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12636 10010 12664 10202
rect 12912 10062 12940 10678
rect 12900 10056 12952 10062
rect 12636 9982 12756 10010
rect 12900 9998 12952 10004
rect 12624 9920 12676 9926
rect 12624 9862 12676 9868
rect 12636 9722 12664 9862
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12728 9586 12756 9982
rect 12900 9920 12952 9926
rect 12900 9862 12952 9868
rect 12716 9580 12768 9586
rect 12716 9522 12768 9528
rect 12208 9222 12214 9274
rect 12266 9222 12278 9274
rect 12330 9222 12342 9274
rect 12394 9222 12406 9274
rect 12458 9222 12470 9274
rect 12522 9222 12528 9274
rect 12072 8968 12124 8974
rect 12072 8910 12124 8916
rect 11888 8492 11940 8498
rect 11888 8434 11940 8440
rect 11980 8492 12032 8498
rect 11980 8434 12032 8440
rect 11704 8356 11756 8362
rect 11704 8298 11756 8304
rect 11336 7948 11388 7954
rect 11336 7890 11388 7896
rect 11716 7886 11744 8298
rect 11992 8090 12020 8434
rect 11980 8084 12032 8090
rect 11980 8026 12032 8032
rect 11060 7880 11112 7886
rect 10690 7848 10746 7857
rect 11060 7822 11112 7828
rect 11704 7880 11756 7886
rect 11704 7822 11756 7828
rect 11888 7880 11940 7886
rect 11992 7868 12020 8026
rect 11940 7840 12020 7868
rect 11888 7822 11940 7828
rect 10690 7783 10692 7792
rect 10744 7783 10746 7792
rect 10692 7754 10744 7760
rect 11716 7750 11744 7822
rect 11704 7744 11756 7750
rect 11704 7686 11756 7692
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 10508 7268 10560 7274
rect 10508 7210 10560 7216
rect 10520 7002 10548 7210
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 11152 6860 11204 6866
rect 11152 6802 11204 6808
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10968 6792 11020 6798
rect 10968 6734 11020 6740
rect 10244 6458 10272 6734
rect 10232 6452 10284 6458
rect 10232 6394 10284 6400
rect 10244 5710 10272 6394
rect 10324 5772 10376 5778
rect 10324 5714 10376 5720
rect 10232 5704 10284 5710
rect 10232 5646 10284 5652
rect 10244 5234 10272 5646
rect 10336 5370 10364 5714
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 10232 5228 10284 5234
rect 10232 5170 10284 5176
rect 10230 4856 10286 4865
rect 10230 4791 10286 4800
rect 10244 4049 10272 4791
rect 10336 4622 10364 5306
rect 10428 5234 10456 6734
rect 10600 6724 10652 6730
rect 10600 6666 10652 6672
rect 10612 6361 10640 6666
rect 10598 6352 10654 6361
rect 10980 6322 11008 6734
rect 10598 6287 10600 6296
rect 10652 6287 10654 6296
rect 10968 6316 11020 6322
rect 10600 6258 10652 6264
rect 10968 6258 11020 6264
rect 10876 5704 10928 5710
rect 10876 5646 10928 5652
rect 10600 5636 10652 5642
rect 10600 5578 10652 5584
rect 10416 5228 10468 5234
rect 10416 5170 10468 5176
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10336 4214 10364 4558
rect 10428 4486 10456 5170
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10612 4282 10640 5578
rect 10784 5568 10836 5574
rect 10784 5510 10836 5516
rect 10692 5228 10744 5234
rect 10692 5170 10744 5176
rect 10704 4622 10732 5170
rect 10692 4616 10744 4622
rect 10692 4558 10744 4564
rect 10692 4480 10744 4486
rect 10692 4422 10744 4428
rect 10600 4276 10652 4282
rect 10600 4218 10652 4224
rect 10324 4208 10376 4214
rect 10324 4150 10376 4156
rect 10704 4146 10732 4422
rect 10600 4140 10652 4146
rect 10600 4082 10652 4088
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10230 4040 10286 4049
rect 10230 3975 10286 3984
rect 10416 3732 10468 3738
rect 10416 3674 10468 3680
rect 10428 3058 10456 3674
rect 10612 3194 10640 4082
rect 10704 3670 10732 4082
rect 10796 4078 10824 5510
rect 10888 4826 10916 5646
rect 10968 5568 11020 5574
rect 10968 5510 11020 5516
rect 10876 4820 10928 4826
rect 10876 4762 10928 4768
rect 10980 4622 11008 5510
rect 10968 4616 11020 4622
rect 10968 4558 11020 4564
rect 10876 4548 10928 4554
rect 10876 4490 10928 4496
rect 10888 4214 10916 4490
rect 10876 4208 10928 4214
rect 10876 4150 10928 4156
rect 10784 4072 10836 4078
rect 10784 4014 10836 4020
rect 10692 3664 10744 3670
rect 10692 3606 10744 3612
rect 10600 3188 10652 3194
rect 10600 3130 10652 3136
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10704 2650 10732 3606
rect 10876 3528 10928 3534
rect 10876 3470 10928 3476
rect 10888 3058 10916 3470
rect 10876 3052 10928 3058
rect 10876 2994 10928 3000
rect 10784 2984 10836 2990
rect 10784 2926 10836 2932
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10796 2564 10824 2926
rect 10888 2689 10916 2994
rect 10980 2922 11008 4558
rect 11060 3596 11112 3602
rect 11060 3538 11112 3544
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10874 2680 10930 2689
rect 10874 2615 10930 2624
rect 10796 2536 10916 2564
rect 10692 2440 10744 2446
rect 10414 2408 10470 2417
rect 10692 2382 10744 2388
rect 10414 2343 10470 2352
rect 10428 2310 10456 2343
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 10704 2258 10732 2382
rect 10888 2281 10916 2536
rect 10874 2272 10930 2281
rect 10704 2230 10824 2258
rect 10140 2100 10192 2106
rect 10140 2042 10192 2048
rect 10048 1964 10100 1970
rect 10048 1906 10100 1912
rect 9956 1760 10008 1766
rect 9956 1702 10008 1708
rect 9968 1358 9996 1702
rect 10690 1592 10746 1601
rect 10796 1562 10824 2230
rect 10874 2207 10930 2216
rect 11072 1970 11100 3538
rect 11164 3058 11192 6802
rect 11624 6798 11652 7278
rect 11716 6866 11744 7686
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11704 6860 11756 6866
rect 11704 6802 11756 6808
rect 11612 6792 11664 6798
rect 11532 6752 11612 6780
rect 11426 4720 11482 4729
rect 11426 4655 11482 4664
rect 11440 4622 11468 4655
rect 11428 4616 11480 4622
rect 11428 4558 11480 4564
rect 11244 4480 11296 4486
rect 11244 4422 11296 4428
rect 11256 4282 11284 4422
rect 11244 4276 11296 4282
rect 11244 4218 11296 4224
rect 11428 3460 11480 3466
rect 11428 3402 11480 3408
rect 11152 3052 11204 3058
rect 11152 2994 11204 3000
rect 11336 2916 11388 2922
rect 11336 2858 11388 2864
rect 11152 2440 11204 2446
rect 11152 2382 11204 2388
rect 11164 1970 11192 2382
rect 11348 2378 11376 2858
rect 11440 2825 11468 3402
rect 11426 2816 11482 2825
rect 11426 2751 11482 2760
rect 11532 2650 11560 6752
rect 11612 6734 11664 6740
rect 11796 6792 11848 6798
rect 11796 6734 11848 6740
rect 11702 5944 11758 5953
rect 11702 5879 11758 5888
rect 11716 5846 11744 5879
rect 11704 5840 11756 5846
rect 11704 5782 11756 5788
rect 11612 5704 11664 5710
rect 11612 5646 11664 5652
rect 11624 5302 11652 5646
rect 11704 5568 11756 5574
rect 11704 5510 11756 5516
rect 11612 5296 11664 5302
rect 11612 5238 11664 5244
rect 11624 3738 11652 5238
rect 11716 4758 11744 5510
rect 11704 4752 11756 4758
rect 11704 4694 11756 4700
rect 11716 4622 11744 4694
rect 11704 4616 11756 4622
rect 11704 4558 11756 4564
rect 11704 4480 11756 4486
rect 11704 4422 11756 4428
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11520 2644 11572 2650
rect 11440 2604 11520 2632
rect 11336 2372 11388 2378
rect 11336 2314 11388 2320
rect 11440 2310 11468 2604
rect 11520 2586 11572 2592
rect 11716 2530 11744 4422
rect 11532 2502 11744 2530
rect 11428 2304 11480 2310
rect 11428 2246 11480 2252
rect 11060 1964 11112 1970
rect 11060 1906 11112 1912
rect 11152 1964 11204 1970
rect 11152 1906 11204 1912
rect 10690 1527 10692 1536
rect 10744 1527 10746 1536
rect 10784 1556 10836 1562
rect 10692 1498 10744 1504
rect 10784 1498 10836 1504
rect 10874 1456 10930 1465
rect 10874 1391 10876 1400
rect 10928 1391 10930 1400
rect 10876 1362 10928 1368
rect 11532 1358 11560 2502
rect 11808 2122 11836 6734
rect 11900 5778 11928 7278
rect 11992 5846 12020 7840
rect 12084 6934 12112 8910
rect 12208 8186 12528 9222
rect 12728 8974 12756 9522
rect 12912 9450 12940 9862
rect 12900 9444 12952 9450
rect 12900 9386 12952 9392
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 12808 8492 12860 8498
rect 12808 8434 12860 8440
rect 12208 8134 12214 8186
rect 12266 8134 12278 8186
rect 12330 8134 12342 8186
rect 12394 8134 12406 8186
rect 12458 8134 12470 8186
rect 12522 8134 12528 8186
rect 12208 7098 12528 8134
rect 12636 7886 12664 8434
rect 12820 7954 12848 8434
rect 12912 8090 12940 9386
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 12808 7948 12860 7954
rect 12808 7890 12860 7896
rect 12624 7880 12676 7886
rect 12624 7822 12676 7828
rect 12208 7046 12214 7098
rect 12266 7046 12278 7098
rect 12330 7046 12342 7098
rect 12394 7046 12406 7098
rect 12458 7046 12470 7098
rect 12522 7046 12528 7098
rect 12072 6928 12124 6934
rect 12072 6870 12124 6876
rect 12072 6248 12124 6254
rect 12072 6190 12124 6196
rect 12084 5914 12112 6190
rect 12208 6010 12528 7046
rect 12636 6866 12664 7822
rect 13004 7546 13032 8774
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12992 7540 13044 7546
rect 12992 7482 13044 7488
rect 12728 7342 12756 7482
rect 12716 7336 12768 7342
rect 12716 7278 12768 7284
rect 12624 6860 12676 6866
rect 12624 6802 12676 6808
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12208 5958 12214 6010
rect 12266 5958 12278 6010
rect 12330 5958 12342 6010
rect 12394 5958 12406 6010
rect 12458 5958 12470 6010
rect 12522 5958 12528 6010
rect 12072 5908 12124 5914
rect 12072 5850 12124 5856
rect 11980 5840 12032 5846
rect 11980 5782 12032 5788
rect 11888 5772 11940 5778
rect 11888 5714 11940 5720
rect 11980 5704 12032 5710
rect 11980 5646 12032 5652
rect 11992 5234 12020 5646
rect 11980 5228 12032 5234
rect 12032 5188 12112 5216
rect 11980 5170 12032 5176
rect 11888 5092 11940 5098
rect 11888 5034 11940 5040
rect 11900 4554 11928 5034
rect 11980 5024 12032 5030
rect 11980 4966 12032 4972
rect 11992 4690 12020 4966
rect 11980 4684 12032 4690
rect 11980 4626 12032 4632
rect 11888 4548 11940 4554
rect 11888 4490 11940 4496
rect 11900 4078 11928 4490
rect 11980 4140 12032 4146
rect 11980 4082 12032 4088
rect 11888 4072 11940 4078
rect 11992 4049 12020 4082
rect 12084 4078 12112 5188
rect 12208 4922 12528 5958
rect 12624 5704 12676 5710
rect 12624 5646 12676 5652
rect 12636 5370 12664 5646
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12728 5370 12756 5578
rect 12820 5574 12848 6734
rect 12992 6724 13044 6730
rect 12992 6666 13044 6672
rect 13004 5642 13032 6666
rect 12992 5636 13044 5642
rect 12992 5578 13044 5584
rect 12808 5568 12860 5574
rect 12808 5510 12860 5516
rect 12624 5364 12676 5370
rect 12624 5306 12676 5312
rect 12716 5364 12768 5370
rect 12716 5306 12768 5312
rect 12716 5160 12768 5166
rect 12716 5102 12768 5108
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12208 4870 12214 4922
rect 12266 4870 12278 4922
rect 12330 4870 12342 4922
rect 12394 4870 12406 4922
rect 12458 4870 12470 4922
rect 12522 4870 12528 4922
rect 12208 4518 12528 4870
rect 12728 4826 12756 5102
rect 12820 5030 12848 5102
rect 12808 5024 12860 5030
rect 12808 4966 12860 4972
rect 12820 4865 12848 4966
rect 12806 4856 12862 4865
rect 12716 4820 12768 4826
rect 12806 4791 12862 4800
rect 12716 4762 12768 4768
rect 12624 4752 12676 4758
rect 12624 4694 12676 4700
rect 12208 4462 12220 4518
rect 12276 4462 12300 4518
rect 12356 4462 12380 4518
rect 12436 4462 12460 4518
rect 12516 4462 12528 4518
rect 12208 4438 12528 4462
rect 12208 4382 12220 4438
rect 12276 4382 12300 4438
rect 12356 4382 12380 4438
rect 12436 4382 12460 4438
rect 12516 4382 12528 4438
rect 12208 4358 12528 4382
rect 12208 4302 12220 4358
rect 12276 4302 12300 4358
rect 12356 4302 12380 4358
rect 12436 4302 12460 4358
rect 12516 4302 12528 4358
rect 12208 4278 12528 4302
rect 12208 4222 12220 4278
rect 12276 4222 12300 4278
rect 12356 4222 12380 4278
rect 12436 4222 12460 4278
rect 12516 4222 12528 4278
rect 12072 4072 12124 4078
rect 11888 4014 11940 4020
rect 11978 4040 12034 4049
rect 12072 4014 12124 4020
rect 11978 3975 12034 3984
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 11900 3097 11928 3878
rect 12084 3398 12112 4014
rect 12208 3834 12528 4222
rect 12208 3782 12214 3834
rect 12266 3782 12278 3834
rect 12330 3782 12342 3834
rect 12394 3782 12406 3834
rect 12458 3782 12470 3834
rect 12522 3782 12528 3834
rect 12072 3392 12124 3398
rect 12072 3334 12124 3340
rect 11886 3088 11942 3097
rect 11886 3023 11942 3032
rect 11888 2984 11940 2990
rect 11888 2926 11940 2932
rect 11624 2106 11836 2122
rect 11612 2100 11836 2106
rect 11664 2094 11836 2100
rect 11612 2042 11664 2048
rect 11900 1850 11928 2926
rect 12208 2746 12528 3782
rect 12208 2694 12214 2746
rect 12266 2694 12278 2746
rect 12330 2694 12342 2746
rect 12394 2694 12406 2746
rect 12458 2694 12470 2746
rect 12522 2694 12528 2746
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 2106 12020 2246
rect 11980 2100 12032 2106
rect 11980 2042 12032 2048
rect 12072 1964 12124 1970
rect 11808 1822 11928 1850
rect 11992 1924 12072 1952
rect 11808 1766 11836 1822
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11992 1494 12020 1924
rect 12072 1906 12124 1912
rect 12072 1828 12124 1834
rect 12072 1770 12124 1776
rect 12084 1601 12112 1770
rect 12208 1658 12528 2694
rect 12636 2582 12664 4694
rect 12728 4146 12756 4762
rect 12808 4616 12860 4622
rect 12808 4558 12860 4564
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12820 4078 12848 4558
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 12808 4072 12860 4078
rect 12808 4014 12860 4020
rect 12716 4004 12768 4010
rect 12716 3946 12768 3952
rect 12728 3738 12756 3946
rect 12716 3732 12768 3738
rect 12716 3674 12768 3680
rect 12728 3126 12756 3674
rect 12716 3120 12768 3126
rect 12716 3062 12768 3068
rect 12820 3058 12848 4014
rect 12912 3466 12940 4490
rect 12900 3460 12952 3466
rect 12900 3402 12952 3408
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 12912 2990 12940 3402
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12624 2576 12676 2582
rect 12624 2518 12676 2524
rect 12624 2440 12676 2446
rect 12622 2408 12624 2417
rect 12676 2408 12678 2417
rect 12622 2343 12678 2352
rect 12208 1606 12214 1658
rect 12266 1606 12278 1658
rect 12330 1606 12342 1658
rect 12394 1606 12406 1658
rect 12458 1606 12470 1658
rect 12522 1606 12528 1658
rect 12070 1592 12126 1601
rect 12070 1527 12126 1536
rect 11980 1488 12032 1494
rect 12072 1488 12124 1494
rect 11980 1430 12032 1436
rect 12070 1456 12072 1465
rect 12124 1456 12126 1465
rect 11992 1358 12020 1430
rect 12070 1391 12126 1400
rect 9956 1352 10008 1358
rect 11060 1352 11112 1358
rect 9956 1294 10008 1300
rect 11058 1320 11060 1329
rect 11520 1352 11572 1358
rect 11112 1320 11114 1329
rect 11520 1294 11572 1300
rect 11888 1352 11940 1358
rect 11888 1294 11940 1300
rect 11980 1352 12032 1358
rect 11980 1294 12032 1300
rect 11058 1255 11114 1264
rect 11900 800 11928 1294
rect 12208 1040 12528 1606
rect 12636 1358 12664 2343
rect 12728 1358 12756 2926
rect 12806 2544 12862 2553
rect 12806 2479 12862 2488
rect 12820 2378 12848 2479
rect 13004 2446 13032 5578
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 12808 2372 12860 2378
rect 12808 2314 12860 2320
rect 12624 1352 12676 1358
rect 12624 1294 12676 1300
rect 12716 1352 12768 1358
rect 12716 1294 12768 1300
rect 13096 1018 13124 10798
rect 13268 10668 13320 10674
rect 13268 10610 13320 10616
rect 13280 10266 13308 10610
rect 13360 10464 13412 10470
rect 13360 10406 13412 10412
rect 13268 10260 13320 10266
rect 13268 10202 13320 10208
rect 13280 9722 13308 10202
rect 13372 10130 13400 10406
rect 13360 10124 13412 10130
rect 13360 10066 13412 10072
rect 13464 10010 13492 11070
rect 13556 10198 13584 12174
rect 13728 12096 13780 12102
rect 13728 12038 13780 12044
rect 13636 11144 13688 11150
rect 13636 11086 13688 11092
rect 13544 10192 13596 10198
rect 13544 10134 13596 10140
rect 13648 10130 13676 11086
rect 13740 10674 13768 12038
rect 13832 11898 13860 13670
rect 13924 13326 13952 13874
rect 14004 13864 14056 13870
rect 14002 13832 14004 13841
rect 14056 13832 14058 13841
rect 14002 13767 14058 13776
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13924 12986 13952 13262
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 14016 12374 14044 13767
rect 14476 13530 14504 17614
rect 14648 17196 14700 17202
rect 14648 17138 14700 17144
rect 15568 17196 15620 17202
rect 15568 17138 15620 17144
rect 14660 16590 14688 17138
rect 15200 17128 15252 17134
rect 15200 17070 15252 17076
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 15212 16522 15240 17070
rect 15580 16794 15608 17138
rect 16132 16794 16160 17614
rect 16208 17434 16528 18470
rect 16776 17814 16804 19200
rect 19352 18358 19380 19200
rect 21456 18692 21508 18698
rect 21456 18634 21508 18640
rect 16948 18352 17000 18358
rect 16948 18294 17000 18300
rect 17500 18352 17552 18358
rect 17500 18294 17552 18300
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 16764 17808 16816 17814
rect 16764 17750 16816 17756
rect 16960 17678 16988 18294
rect 17408 18284 17460 18290
rect 17408 18226 17460 18232
rect 17420 17746 17448 18226
rect 17512 17814 17540 18294
rect 18696 18284 18748 18290
rect 18696 18226 18748 18232
rect 17868 18216 17920 18222
rect 17868 18158 17920 18164
rect 18420 18216 18472 18222
rect 18420 18158 18472 18164
rect 17500 17808 17552 17814
rect 17500 17750 17552 17756
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16208 17382 16214 17434
rect 16266 17382 16278 17434
rect 16330 17382 16342 17434
rect 16394 17382 16406 17434
rect 16458 17382 16470 17434
rect 16522 17382 16528 17434
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 16120 16788 16172 16794
rect 16120 16730 16172 16736
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 16028 16584 16080 16590
rect 16028 16526 16080 16532
rect 16120 16584 16172 16590
rect 16120 16526 16172 16532
rect 15200 16516 15252 16522
rect 15200 16458 15252 16464
rect 15304 16153 15332 16526
rect 15660 16516 15712 16522
rect 15660 16458 15712 16464
rect 15290 16144 15346 16153
rect 15108 16108 15160 16114
rect 15290 16079 15346 16088
rect 15476 16108 15528 16114
rect 15108 16050 15160 16056
rect 15476 16050 15528 16056
rect 14832 15700 14884 15706
rect 14832 15642 14884 15648
rect 14844 15609 14872 15642
rect 15016 15632 15068 15638
rect 14830 15600 14886 15609
rect 15016 15574 15068 15580
rect 14830 15535 14886 15544
rect 14924 15496 14976 15502
rect 14646 15464 14702 15473
rect 14924 15438 14976 15444
rect 14646 15399 14648 15408
rect 14700 15399 14702 15408
rect 14740 15428 14792 15434
rect 14648 15370 14700 15376
rect 14740 15370 14792 15376
rect 14752 15094 14780 15370
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14740 15088 14792 15094
rect 14740 15030 14792 15036
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14660 14346 14688 14894
rect 14648 14340 14700 14346
rect 14648 14282 14700 14288
rect 14844 13734 14872 15302
rect 14936 14958 14964 15438
rect 15028 15162 15056 15574
rect 15120 15570 15148 16050
rect 15200 15700 15252 15706
rect 15200 15642 15252 15648
rect 15108 15564 15160 15570
rect 15108 15506 15160 15512
rect 15120 15366 15148 15506
rect 15108 15360 15160 15366
rect 15108 15302 15160 15308
rect 15016 15156 15068 15162
rect 15016 15098 15068 15104
rect 14924 14952 14976 14958
rect 14924 14894 14976 14900
rect 14936 13870 14964 14894
rect 15016 14816 15068 14822
rect 15016 14758 15068 14764
rect 15028 14414 15056 14758
rect 15120 14414 15148 15302
rect 15212 14822 15240 15642
rect 15488 15586 15516 16050
rect 15672 15910 15700 16458
rect 15856 16046 15884 16526
rect 16040 16454 16068 16526
rect 16028 16448 16080 16454
rect 16028 16390 16080 16396
rect 16040 16250 16068 16390
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15568 15904 15620 15910
rect 15568 15846 15620 15852
rect 15660 15904 15712 15910
rect 15660 15846 15712 15852
rect 15304 15558 15516 15586
rect 15580 15586 15608 15846
rect 16132 15706 16160 16526
rect 16208 16518 16528 17382
rect 17684 16788 17736 16794
rect 17684 16730 17736 16736
rect 17696 16590 17724 16730
rect 17684 16584 17736 16590
rect 17684 16526 17736 16532
rect 16208 16462 16220 16518
rect 16276 16462 16300 16518
rect 16356 16462 16380 16518
rect 16436 16462 16460 16518
rect 16516 16462 16528 16518
rect 16208 16438 16528 16462
rect 17880 16454 17908 18158
rect 18328 18148 18380 18154
rect 18328 18090 18380 18096
rect 18340 17338 18368 18090
rect 18328 17332 18380 17338
rect 18328 17274 18380 17280
rect 18236 17196 18288 17202
rect 18236 17138 18288 17144
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17972 16454 18000 16594
rect 18248 16590 18276 17138
rect 18236 16584 18288 16590
rect 18236 16526 18288 16532
rect 18340 16522 18368 17274
rect 18432 16794 18460 18158
rect 18708 17270 18736 18226
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 18800 17678 18828 18022
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18696 17264 18748 17270
rect 18696 17206 18748 17212
rect 19352 16794 19380 18294
rect 19984 18148 20036 18154
rect 19984 18090 20036 18096
rect 19432 18080 19484 18086
rect 19432 18022 19484 18028
rect 19800 18080 19852 18086
rect 19800 18022 19852 18028
rect 18420 16788 18472 16794
rect 18420 16730 18472 16736
rect 18696 16788 18748 16794
rect 18696 16730 18748 16736
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 18708 16590 18736 16730
rect 18696 16584 18748 16590
rect 18696 16526 18748 16532
rect 18328 16516 18380 16522
rect 18328 16458 18380 16464
rect 19444 16454 19472 18022
rect 19616 17060 19668 17066
rect 19616 17002 19668 17008
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 16208 16382 16220 16438
rect 16276 16382 16300 16438
rect 16356 16382 16380 16438
rect 16436 16382 16460 16438
rect 16516 16382 16528 16438
rect 17868 16448 17920 16454
rect 17868 16390 17920 16396
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 19432 16448 19484 16454
rect 19432 16390 19484 16396
rect 16208 16358 16528 16382
rect 16208 16346 16220 16358
rect 16276 16346 16300 16358
rect 16356 16346 16380 16358
rect 16436 16346 16460 16358
rect 16516 16346 16528 16358
rect 16208 16294 16214 16346
rect 16276 16302 16278 16346
rect 16458 16302 16460 16346
rect 16266 16294 16278 16302
rect 16330 16294 16342 16302
rect 16394 16294 16406 16302
rect 16458 16294 16470 16302
rect 16522 16294 16528 16346
rect 16208 16278 16528 16294
rect 16208 16222 16220 16278
rect 16276 16222 16300 16278
rect 16356 16222 16380 16278
rect 16436 16222 16460 16278
rect 16516 16222 16528 16278
rect 16120 15700 16172 15706
rect 16120 15642 16172 15648
rect 15934 15600 15990 15609
rect 15580 15558 15884 15586
rect 15304 15026 15332 15558
rect 15384 15496 15436 15502
rect 15384 15438 15436 15444
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15200 14816 15252 14822
rect 15200 14758 15252 14764
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15108 14408 15160 14414
rect 15108 14350 15160 14356
rect 15016 13932 15068 13938
rect 15016 13874 15068 13880
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 14924 13864 14976 13870
rect 14924 13806 14976 13812
rect 15028 13734 15056 13874
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 15016 13728 15068 13734
rect 15016 13670 15068 13676
rect 14464 13524 14516 13530
rect 14464 13466 14516 13472
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14660 12850 14688 13126
rect 14844 12850 14872 13670
rect 15212 13530 15240 13874
rect 15200 13524 15252 13530
rect 15200 13466 15252 13472
rect 15304 13394 15332 14962
rect 15396 14482 15424 15438
rect 15488 14958 15516 15438
rect 15660 15156 15712 15162
rect 15660 15098 15712 15104
rect 15568 15088 15620 15094
rect 15568 15030 15620 15036
rect 15476 14952 15528 14958
rect 15476 14894 15528 14900
rect 15488 14618 15516 14894
rect 15476 14612 15528 14618
rect 15476 14554 15528 14560
rect 15384 14476 15436 14482
rect 15384 14418 15436 14424
rect 15488 14346 15516 14554
rect 15476 14340 15528 14346
rect 15476 14282 15528 14288
rect 15580 14226 15608 15030
rect 15488 14198 15608 14226
rect 15292 13388 15344 13394
rect 15292 13330 15344 13336
rect 15016 13320 15068 13326
rect 15016 13262 15068 13268
rect 14648 12844 14700 12850
rect 14648 12786 14700 12792
rect 14832 12844 14884 12850
rect 14832 12786 14884 12792
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 14096 12776 14148 12782
rect 14096 12718 14148 12724
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13820 11892 13872 11898
rect 13820 11834 13872 11840
rect 13820 11144 13872 11150
rect 13820 11086 13872 11092
rect 13728 10668 13780 10674
rect 13728 10610 13780 10616
rect 13636 10124 13688 10130
rect 13636 10066 13688 10072
rect 13464 9982 13676 10010
rect 13832 9994 13860 11086
rect 14016 10062 14044 12310
rect 14108 12102 14136 12718
rect 14844 12306 14872 12786
rect 14936 12646 14964 12786
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14832 12300 14884 12306
rect 14832 12242 14884 12248
rect 14648 12232 14700 12238
rect 14648 12174 14700 12180
rect 14096 12096 14148 12102
rect 14096 12038 14148 12044
rect 14660 11830 14688 12174
rect 14844 12170 14872 12242
rect 14936 12238 14964 12582
rect 15028 12238 15056 13262
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 15016 12232 15068 12238
rect 15120 12220 15148 12582
rect 15292 12232 15344 12238
rect 15120 12192 15292 12220
rect 15016 12174 15068 12180
rect 15292 12174 15344 12180
rect 14832 12164 14884 12170
rect 14832 12106 14884 12112
rect 15028 12102 15056 12174
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14464 11688 14516 11694
rect 14464 11630 14516 11636
rect 14648 11688 14700 11694
rect 14648 11630 14700 11636
rect 14004 10056 14056 10062
rect 14004 9998 14056 10004
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13464 9110 13492 9318
rect 13452 9104 13504 9110
rect 13452 9046 13504 9052
rect 13452 8288 13504 8294
rect 13452 8230 13504 8236
rect 13544 8288 13596 8294
rect 13544 8230 13596 8236
rect 13464 7954 13492 8230
rect 13452 7948 13504 7954
rect 13452 7890 13504 7896
rect 13176 7880 13228 7886
rect 13174 7848 13176 7857
rect 13228 7848 13230 7857
rect 13174 7783 13230 7792
rect 13556 7410 13584 8230
rect 13544 7404 13596 7410
rect 13544 7346 13596 7352
rect 13360 6724 13412 6730
rect 13360 6666 13412 6672
rect 13372 6322 13400 6666
rect 13360 6316 13412 6322
rect 13360 6258 13412 6264
rect 13360 6112 13412 6118
rect 13360 6054 13412 6060
rect 13372 5710 13400 6054
rect 13360 5704 13412 5710
rect 13360 5646 13412 5652
rect 13176 5568 13228 5574
rect 13176 5510 13228 5516
rect 13188 2582 13216 5510
rect 13544 5228 13596 5234
rect 13544 5170 13596 5176
rect 13452 5160 13504 5166
rect 13452 5102 13504 5108
rect 13358 4720 13414 4729
rect 13358 4655 13414 4664
rect 13372 4622 13400 4655
rect 13464 4622 13492 5102
rect 13556 4622 13584 5170
rect 13360 4616 13412 4622
rect 13360 4558 13412 4564
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13544 4616 13596 4622
rect 13544 4558 13596 4564
rect 13648 4162 13676 9982
rect 13820 9988 13872 9994
rect 13820 9930 13872 9936
rect 14476 9625 14504 11630
rect 14660 9654 14688 11630
rect 15028 11218 15056 12038
rect 15488 11898 15516 14198
rect 15672 14074 15700 15098
rect 15764 14278 15792 15438
rect 15856 14958 15884 15558
rect 15934 15535 15990 15544
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15856 14657 15884 14894
rect 15842 14648 15898 14657
rect 15842 14583 15898 14592
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15660 14068 15712 14074
rect 15660 14010 15712 14016
rect 15764 13394 15792 14214
rect 15856 13569 15884 14583
rect 15842 13560 15898 13569
rect 15842 13495 15898 13504
rect 15752 13388 15804 13394
rect 15752 13330 15804 13336
rect 15948 13326 15976 15535
rect 16028 15360 16080 15366
rect 16028 15302 16080 15308
rect 16040 15162 16068 15302
rect 16208 15258 16528 16222
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 16762 16144 16818 16153
rect 16580 16108 16632 16114
rect 16762 16079 16818 16088
rect 18236 16108 18288 16114
rect 16580 16050 16632 16056
rect 16592 15706 16620 16050
rect 16580 15700 16632 15706
rect 16580 15642 16632 15648
rect 16776 15638 16804 16079
rect 18236 16050 18288 16056
rect 17040 16040 17092 16046
rect 17040 15982 17092 15988
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 16764 15632 16816 15638
rect 16578 15600 16634 15609
rect 16764 15574 16816 15580
rect 16578 15535 16634 15544
rect 16592 15502 16620 15535
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16948 15428 17000 15434
rect 16948 15370 17000 15376
rect 16208 15206 16214 15258
rect 16266 15206 16278 15258
rect 16330 15206 16342 15258
rect 16394 15206 16406 15258
rect 16458 15206 16470 15258
rect 16522 15206 16528 15258
rect 16028 15156 16080 15162
rect 16028 15098 16080 15104
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16132 13938 16160 14962
rect 16208 14170 16528 15206
rect 16960 15162 16988 15370
rect 16948 15156 17000 15162
rect 16948 15098 17000 15104
rect 17052 15026 17080 15982
rect 17132 15700 17184 15706
rect 17132 15642 17184 15648
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17040 14816 17092 14822
rect 17040 14758 17092 14764
rect 16946 14648 17002 14657
rect 16946 14583 16948 14592
rect 17000 14583 17002 14592
rect 16948 14554 17000 14560
rect 16948 14408 17000 14414
rect 16208 14118 16214 14170
rect 16266 14118 16278 14170
rect 16330 14118 16342 14170
rect 16394 14118 16406 14170
rect 16458 14118 16470 14170
rect 16522 14118 16528 14170
rect 16120 13932 16172 13938
rect 16120 13874 16172 13880
rect 16132 13530 16160 13874
rect 16120 13524 16172 13530
rect 16120 13466 16172 13472
rect 15936 13320 15988 13326
rect 15936 13262 15988 13268
rect 15948 12986 15976 13262
rect 15936 12980 15988 12986
rect 15988 12940 16068 12968
rect 15936 12922 15988 12928
rect 15660 12776 15712 12782
rect 15660 12718 15712 12724
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 15476 11892 15528 11898
rect 15476 11834 15528 11840
rect 15108 11756 15160 11762
rect 15108 11698 15160 11704
rect 15120 11558 15148 11698
rect 15568 11688 15620 11694
rect 15568 11630 15620 11636
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15120 10742 15148 11494
rect 15384 11076 15436 11082
rect 15384 11018 15436 11024
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15200 10532 15252 10538
rect 15200 10474 15252 10480
rect 14648 9648 14700 9654
rect 14462 9616 14518 9625
rect 14004 9580 14056 9586
rect 14648 9590 14700 9596
rect 14462 9551 14464 9560
rect 14004 9522 14056 9528
rect 14516 9551 14518 9560
rect 14464 9522 14516 9528
rect 13728 9376 13780 9382
rect 13728 9318 13780 9324
rect 13740 8022 13768 9318
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13728 8016 13780 8022
rect 13728 7958 13780 7964
rect 13728 7880 13780 7886
rect 13832 7868 13860 8434
rect 13780 7840 13860 7868
rect 13728 7822 13780 7828
rect 13740 7410 13768 7822
rect 13728 7404 13780 7410
rect 13780 7364 13952 7392
rect 13728 7346 13780 7352
rect 13728 6928 13780 6934
rect 13728 6870 13780 6876
rect 13740 5710 13768 6870
rect 13924 6254 13952 7364
rect 13912 6248 13964 6254
rect 13912 6190 13964 6196
rect 14016 6186 14044 9522
rect 15212 9466 15240 10474
rect 15304 10130 15332 10610
rect 15292 10124 15344 10130
rect 15292 10066 15344 10072
rect 15396 10062 15424 11018
rect 15580 10810 15608 11630
rect 15672 11150 15700 12718
rect 15752 12708 15804 12714
rect 15752 12650 15804 12656
rect 15764 12442 15792 12650
rect 15856 12442 15884 12718
rect 15936 12640 15988 12646
rect 15936 12582 15988 12588
rect 15752 12436 15804 12442
rect 15752 12378 15804 12384
rect 15844 12436 15896 12442
rect 15844 12378 15896 12384
rect 15948 12306 15976 12582
rect 15936 12300 15988 12306
rect 15936 12242 15988 12248
rect 15752 12232 15804 12238
rect 15752 12174 15804 12180
rect 15660 11144 15712 11150
rect 15660 11086 15712 11092
rect 15660 11008 15712 11014
rect 15660 10950 15712 10956
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 15672 10198 15700 10950
rect 15660 10192 15712 10198
rect 15660 10134 15712 10140
rect 15384 10056 15436 10062
rect 15384 9998 15436 10004
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9586 15332 9930
rect 15292 9580 15344 9586
rect 15292 9522 15344 9528
rect 15396 9568 15424 9998
rect 15764 9926 15792 12174
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15856 11762 15884 12038
rect 15844 11756 15896 11762
rect 15844 11698 15896 11704
rect 15856 11014 15884 11698
rect 15948 11694 15976 12242
rect 16040 12238 16068 12940
rect 16132 12850 16160 13466
rect 16208 13082 16528 14118
rect 16684 14368 16948 14396
rect 16684 14074 16712 14368
rect 16948 14350 17000 14356
rect 16764 14272 16816 14278
rect 16764 14214 16816 14220
rect 16776 14074 16804 14214
rect 17052 14074 17080 14758
rect 17144 14414 17172 15642
rect 17328 15502 17356 15982
rect 17316 15496 17368 15502
rect 18144 15496 18196 15502
rect 17316 15438 17368 15444
rect 18142 15464 18144 15473
rect 18196 15464 18198 15473
rect 17328 15162 17356 15438
rect 18142 15399 18198 15408
rect 17316 15156 17368 15162
rect 17316 15098 17368 15104
rect 18156 15094 18184 15399
rect 18144 15088 18196 15094
rect 18144 15030 18196 15036
rect 17224 15020 17276 15026
rect 17224 14962 17276 14968
rect 17132 14408 17184 14414
rect 17132 14350 17184 14356
rect 16672 14068 16724 14074
rect 16672 14010 16724 14016
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 17040 14068 17092 14074
rect 17040 14010 17092 14016
rect 17144 13938 17172 14350
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 17132 13932 17184 13938
rect 17132 13874 17184 13880
rect 16672 13864 16724 13870
rect 16672 13806 16724 13812
rect 16684 13394 16712 13806
rect 16960 13530 16988 13874
rect 17144 13802 17172 13874
rect 17132 13796 17184 13802
rect 17132 13738 17184 13744
rect 16948 13524 17000 13530
rect 16948 13466 17000 13472
rect 16672 13388 16724 13394
rect 16672 13330 16724 13336
rect 16208 13030 16214 13082
rect 16266 13030 16278 13082
rect 16330 13030 16342 13082
rect 16394 13030 16406 13082
rect 16458 13030 16470 13082
rect 16522 13030 16528 13082
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16132 12442 16160 12786
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16120 12300 16172 12306
rect 16120 12242 16172 12248
rect 16028 12232 16080 12238
rect 16028 12174 16080 12180
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15936 11552 15988 11558
rect 15936 11494 15988 11500
rect 16028 11552 16080 11558
rect 16028 11494 16080 11500
rect 15844 11008 15896 11014
rect 15844 10950 15896 10956
rect 15948 10606 15976 11494
rect 16040 10810 16068 11494
rect 16028 10804 16080 10810
rect 16028 10746 16080 10752
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15764 9722 15792 9862
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15750 9616 15806 9625
rect 15660 9580 15712 9586
rect 15396 9540 15660 9568
rect 15120 9450 15240 9466
rect 15108 9444 15240 9450
rect 15160 9438 15240 9444
rect 15108 9386 15160 9392
rect 15396 9330 15424 9540
rect 16132 9586 16160 12242
rect 16208 11994 16528 13030
rect 16684 12918 16712 13330
rect 16764 13252 16816 13258
rect 16764 13194 16816 13200
rect 16776 12986 16804 13194
rect 16764 12980 16816 12986
rect 16764 12922 16816 12928
rect 16672 12912 16724 12918
rect 16672 12854 16724 12860
rect 16948 12912 17000 12918
rect 16948 12854 17000 12860
rect 16208 11942 16214 11994
rect 16266 11942 16278 11994
rect 16330 11942 16342 11994
rect 16394 11942 16406 11994
rect 16458 11942 16470 11994
rect 16522 11942 16528 11994
rect 16208 10906 16528 11942
rect 16672 11892 16724 11898
rect 16672 11834 16724 11840
rect 16580 11076 16632 11082
rect 16580 11018 16632 11024
rect 16208 10854 16214 10906
rect 16266 10854 16278 10906
rect 16330 10854 16342 10906
rect 16394 10854 16406 10906
rect 16458 10854 16470 10906
rect 16522 10854 16528 10906
rect 16208 9818 16528 10854
rect 16592 10810 16620 11018
rect 16580 10804 16632 10810
rect 16580 10746 16632 10752
rect 16684 10062 16712 11834
rect 16960 11694 16988 12854
rect 17144 12306 17172 13738
rect 17132 12300 17184 12306
rect 17132 12242 17184 12248
rect 17236 12238 17264 14962
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 18050 14920 18106 14929
rect 17328 14618 17356 14894
rect 17776 14884 17828 14890
rect 18050 14855 18052 14864
rect 17776 14826 17828 14832
rect 18104 14855 18106 14864
rect 18052 14826 18104 14832
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17316 14612 17368 14618
rect 17316 14554 17368 14560
rect 17604 13938 17632 14758
rect 17684 14340 17736 14346
rect 17684 14282 17736 14288
rect 17592 13932 17644 13938
rect 17592 13874 17644 13880
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17328 13433 17356 13806
rect 17314 13424 17370 13433
rect 17314 13359 17370 13368
rect 17498 13424 17554 13433
rect 17498 13359 17500 13368
rect 17552 13359 17554 13368
rect 17500 13330 17552 13336
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17500 12164 17552 12170
rect 17500 12106 17552 12112
rect 16948 11688 17000 11694
rect 16948 11630 17000 11636
rect 16960 11218 16988 11630
rect 16948 11212 17000 11218
rect 16948 11154 17000 11160
rect 16960 10606 16988 11154
rect 16948 10600 17000 10606
rect 16948 10542 17000 10548
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16208 9766 16214 9818
rect 16266 9766 16278 9818
rect 16330 9766 16342 9818
rect 16394 9766 16406 9818
rect 16458 9766 16470 9818
rect 16522 9766 16528 9818
rect 15750 9551 15806 9560
rect 16120 9580 16172 9586
rect 15660 9522 15712 9528
rect 15764 9518 15792 9551
rect 16120 9522 16172 9528
rect 15752 9512 15804 9518
rect 15752 9454 15804 9460
rect 15844 9512 15896 9518
rect 15844 9454 15896 9460
rect 15212 9302 15424 9330
rect 15212 9042 15240 9302
rect 15200 9036 15252 9042
rect 15200 8978 15252 8984
rect 14096 8968 14148 8974
rect 14096 8910 14148 8916
rect 14188 8968 14240 8974
rect 14188 8910 14240 8916
rect 14108 8430 14136 8910
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14108 7886 14136 8366
rect 14200 7886 14228 8910
rect 14372 8900 14424 8906
rect 14372 8842 14424 8848
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 14384 8634 14412 8842
rect 14648 8832 14700 8838
rect 14648 8774 14700 8780
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14372 8628 14424 8634
rect 14372 8570 14424 8576
rect 14660 8430 14688 8774
rect 14752 8498 14780 8774
rect 15212 8634 15240 8842
rect 15856 8634 15884 9454
rect 16208 8730 16528 9766
rect 16580 9376 16632 9382
rect 16580 9318 16632 9324
rect 16592 8906 16620 9318
rect 16960 9042 16988 10542
rect 17328 10266 17356 10542
rect 17316 10260 17368 10266
rect 17316 10202 17368 10208
rect 17512 9994 17540 12106
rect 17604 10266 17632 12378
rect 17696 12306 17724 14282
rect 17788 12782 17816 14826
rect 17960 13320 18012 13326
rect 17958 13288 17960 13297
rect 18012 13288 18014 13297
rect 17958 13223 18014 13232
rect 18052 12912 18104 12918
rect 18052 12854 18104 12860
rect 17776 12776 17828 12782
rect 17776 12718 17828 12724
rect 18064 12374 18092 12854
rect 18248 12434 18276 16050
rect 18432 15094 18460 16186
rect 18972 16176 19024 16182
rect 18972 16118 19024 16124
rect 18604 16108 18656 16114
rect 18604 16050 18656 16056
rect 18616 15638 18644 16050
rect 18788 16040 18840 16046
rect 18788 15982 18840 15988
rect 18696 15972 18748 15978
rect 18696 15914 18748 15920
rect 18708 15638 18736 15914
rect 18800 15706 18828 15982
rect 18788 15700 18840 15706
rect 18788 15642 18840 15648
rect 18604 15632 18656 15638
rect 18604 15574 18656 15580
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18984 15434 19012 16118
rect 19536 16114 19564 16458
rect 19524 16108 19576 16114
rect 19524 16050 19576 16056
rect 19340 16040 19392 16046
rect 19340 15982 19392 15988
rect 19352 15570 19380 15982
rect 19340 15564 19392 15570
rect 19340 15506 19392 15512
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 19248 15428 19300 15434
rect 19248 15370 19300 15376
rect 19260 15162 19288 15370
rect 18788 15156 18840 15162
rect 18788 15098 18840 15104
rect 19248 15156 19300 15162
rect 19248 15098 19300 15104
rect 18420 15088 18472 15094
rect 18420 15030 18472 15036
rect 18512 14340 18564 14346
rect 18512 14282 18564 14288
rect 18328 13932 18380 13938
rect 18328 13874 18380 13880
rect 18340 13394 18368 13874
rect 18418 13424 18474 13433
rect 18328 13388 18380 13394
rect 18418 13359 18420 13368
rect 18328 13330 18380 13336
rect 18472 13359 18474 13368
rect 18420 13330 18472 13336
rect 18524 13258 18552 14282
rect 18512 13252 18564 13258
rect 18512 13194 18564 13200
rect 18248 12406 18368 12434
rect 18052 12368 18104 12374
rect 18052 12310 18104 12316
rect 17684 12300 17736 12306
rect 17684 12242 17736 12248
rect 18340 12238 18368 12406
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17960 12096 18012 12102
rect 17960 12038 18012 12044
rect 17592 10260 17644 10266
rect 17592 10202 17644 10208
rect 17500 9988 17552 9994
rect 17500 9930 17552 9936
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 16948 9036 17000 9042
rect 16948 8978 17000 8984
rect 16580 8900 16632 8906
rect 16580 8842 16632 8848
rect 16208 8678 16214 8730
rect 16266 8678 16278 8730
rect 16330 8678 16342 8730
rect 16394 8678 16406 8730
rect 16458 8678 16470 8730
rect 16522 8678 16528 8730
rect 15200 8628 15252 8634
rect 15200 8570 15252 8576
rect 15844 8628 15896 8634
rect 15844 8570 15896 8576
rect 15476 8560 15528 8566
rect 15476 8502 15528 8508
rect 16208 8518 16528 8678
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 15108 8492 15160 8498
rect 15108 8434 15160 8440
rect 14648 8424 14700 8430
rect 14648 8366 14700 8372
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14924 7948 14976 7954
rect 14924 7890 14976 7896
rect 14096 7880 14148 7886
rect 14096 7822 14148 7828
rect 14188 7880 14240 7886
rect 14188 7822 14240 7828
rect 14200 7154 14228 7822
rect 14740 7812 14792 7818
rect 14740 7754 14792 7760
rect 14462 7576 14518 7585
rect 14752 7546 14780 7754
rect 14462 7511 14518 7520
rect 14740 7540 14792 7546
rect 14476 7478 14504 7511
rect 14740 7482 14792 7488
rect 14936 7478 14964 7890
rect 14280 7472 14332 7478
rect 14278 7440 14280 7449
rect 14464 7472 14516 7478
rect 14332 7440 14334 7449
rect 14924 7472 14976 7478
rect 14464 7414 14516 7420
rect 14922 7440 14924 7449
rect 14976 7440 14978 7449
rect 14278 7375 14334 7384
rect 14922 7375 14978 7384
rect 15028 7206 15056 8230
rect 15120 7585 15148 8434
rect 15488 7954 15516 8502
rect 15752 8492 15804 8498
rect 15752 8434 15804 8440
rect 16208 8462 16220 8518
rect 16276 8462 16300 8518
rect 16356 8462 16380 8518
rect 16436 8462 16460 8518
rect 16516 8462 16528 8518
rect 16672 8560 16724 8566
rect 16672 8502 16724 8508
rect 16208 8438 16528 8462
rect 15476 7948 15528 7954
rect 15476 7890 15528 7896
rect 15764 7818 15792 8434
rect 16120 8424 16172 8430
rect 16120 8366 16172 8372
rect 16208 8382 16220 8438
rect 16276 8382 16300 8438
rect 16356 8382 16380 8438
rect 16436 8382 16460 8438
rect 16516 8382 16528 8438
rect 15936 8356 15988 8362
rect 15936 8298 15988 8304
rect 15948 8090 15976 8298
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15752 7812 15804 7818
rect 15752 7754 15804 7760
rect 15844 7744 15896 7750
rect 15844 7686 15896 7692
rect 15106 7576 15162 7585
rect 15106 7511 15162 7520
rect 15120 7478 15148 7511
rect 15108 7472 15160 7478
rect 15108 7414 15160 7420
rect 15384 7472 15436 7478
rect 15384 7414 15436 7420
rect 15108 7336 15160 7342
rect 15108 7278 15160 7284
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 14108 7126 14228 7154
rect 15016 7200 15068 7206
rect 15016 7142 15068 7148
rect 14108 6798 14136 7126
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 6458 14136 6734
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 14476 6458 14504 6666
rect 14096 6452 14148 6458
rect 14096 6394 14148 6400
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 15120 6322 15148 7278
rect 15200 7200 15252 7206
rect 15200 7142 15252 7148
rect 15212 6730 15240 7142
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14372 6316 14424 6322
rect 15108 6316 15160 6322
rect 14372 6258 14424 6264
rect 15028 6276 15108 6304
rect 14004 6180 14056 6186
rect 14004 6122 14056 6128
rect 14280 6112 14332 6118
rect 14280 6054 14332 6060
rect 14292 5710 14320 6054
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 14280 5704 14332 5710
rect 14280 5646 14332 5652
rect 14384 5302 14412 6258
rect 14832 5568 14884 5574
rect 14832 5510 14884 5516
rect 14844 5302 14872 5510
rect 14372 5296 14424 5302
rect 14372 5238 14424 5244
rect 14832 5296 14884 5302
rect 14832 5238 14884 5244
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13832 4826 13860 5170
rect 13912 5092 13964 5098
rect 13912 5034 13964 5040
rect 13820 4820 13872 4826
rect 13820 4762 13872 4768
rect 13728 4616 13780 4622
rect 13728 4558 13780 4564
rect 13740 4282 13768 4558
rect 13820 4480 13872 4486
rect 13820 4422 13872 4428
rect 13728 4276 13780 4282
rect 13728 4218 13780 4224
rect 13544 4140 13596 4146
rect 13648 4134 13768 4162
rect 13544 4082 13596 4088
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 13464 3641 13492 3878
rect 13450 3632 13506 3641
rect 13556 3602 13584 4082
rect 13636 4004 13688 4010
rect 13636 3946 13688 3952
rect 13648 3602 13676 3946
rect 13450 3567 13506 3576
rect 13544 3596 13596 3602
rect 13544 3538 13596 3544
rect 13636 3596 13688 3602
rect 13636 3538 13688 3544
rect 13360 3188 13412 3194
rect 13360 3130 13412 3136
rect 13268 2984 13320 2990
rect 13268 2926 13320 2932
rect 13176 2576 13228 2582
rect 13176 2518 13228 2524
rect 13280 1834 13308 2926
rect 13372 2446 13400 3130
rect 13452 3120 13504 3126
rect 13452 3062 13504 3068
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13268 1828 13320 1834
rect 13268 1770 13320 1776
rect 13176 1420 13228 1426
rect 13176 1362 13228 1368
rect 13188 1329 13216 1362
rect 13464 1358 13492 3062
rect 13544 2848 13596 2854
rect 13544 2790 13596 2796
rect 13556 2394 13584 2790
rect 13556 2366 13676 2394
rect 13542 2272 13598 2281
rect 13542 2207 13598 2216
rect 13556 1970 13584 2207
rect 13648 1970 13676 2366
rect 13544 1964 13596 1970
rect 13544 1906 13596 1912
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 13648 1834 13676 1906
rect 13636 1828 13688 1834
rect 13636 1770 13688 1776
rect 13452 1352 13504 1358
rect 13174 1320 13230 1329
rect 13452 1294 13504 1300
rect 13174 1255 13230 1264
rect 13084 1012 13136 1018
rect 13084 954 13136 960
rect 13740 950 13768 4134
rect 13832 3602 13860 4422
rect 13924 4282 13952 5034
rect 14280 4752 14332 4758
rect 14280 4694 14332 4700
rect 14292 4622 14320 4694
rect 14384 4622 14412 5238
rect 14740 5160 14792 5166
rect 14740 5102 14792 5108
rect 14462 4720 14518 4729
rect 14462 4655 14464 4664
rect 14516 4655 14518 4664
rect 14464 4626 14516 4632
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14372 4616 14424 4622
rect 14372 4558 14424 4564
rect 14556 4616 14608 4622
rect 14752 4604 14780 5102
rect 14844 4622 14872 5238
rect 15028 5234 15056 6276
rect 15108 6258 15160 6264
rect 15108 5364 15160 5370
rect 15108 5306 15160 5312
rect 15016 5228 15068 5234
rect 15016 5170 15068 5176
rect 15120 4758 15148 5306
rect 15304 5250 15332 7278
rect 15212 5222 15332 5250
rect 15016 4752 15068 4758
rect 15016 4694 15068 4700
rect 15108 4752 15160 4758
rect 15108 4694 15160 4700
rect 15028 4622 15056 4694
rect 14608 4576 14780 4604
rect 14832 4616 14884 4622
rect 14556 4558 14608 4564
rect 14832 4558 14884 4564
rect 14924 4616 14976 4622
rect 14924 4558 14976 4564
rect 15016 4616 15068 4622
rect 15016 4558 15068 4564
rect 14936 4282 14964 4558
rect 13912 4276 13964 4282
rect 13912 4218 13964 4224
rect 14924 4276 14976 4282
rect 14924 4218 14976 4224
rect 14188 3936 14240 3942
rect 14188 3878 14240 3884
rect 13820 3596 13872 3602
rect 13820 3538 13872 3544
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 14004 3052 14056 3058
rect 14004 2994 14056 3000
rect 14016 2582 14044 2994
rect 14004 2576 14056 2582
rect 14004 2518 14056 2524
rect 14108 2106 14136 3470
rect 14200 3058 14228 3878
rect 14280 3528 14332 3534
rect 14280 3470 14332 3476
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14188 3052 14240 3058
rect 14188 2994 14240 3000
rect 14096 2100 14148 2106
rect 14096 2042 14148 2048
rect 14292 1970 14320 3470
rect 14752 2514 14780 3470
rect 14830 3088 14886 3097
rect 14830 3023 14886 3032
rect 14844 2922 14872 3023
rect 14936 2990 14964 4218
rect 15016 4140 15068 4146
rect 15016 4082 15068 4088
rect 14924 2984 14976 2990
rect 14924 2926 14976 2932
rect 14832 2916 14884 2922
rect 14832 2858 14884 2864
rect 15028 2854 15056 4082
rect 15212 4010 15240 5222
rect 15396 5098 15424 7414
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15476 6928 15528 6934
rect 15476 6870 15528 6876
rect 15384 5092 15436 5098
rect 15384 5034 15436 5040
rect 15396 4554 15424 5034
rect 15384 4548 15436 4554
rect 15384 4490 15436 4496
rect 15488 4264 15516 6870
rect 15580 6458 15608 7142
rect 15568 6452 15620 6458
rect 15568 6394 15620 6400
rect 15856 6322 15884 7686
rect 16028 7472 16080 7478
rect 16028 7414 16080 7420
rect 15936 7200 15988 7206
rect 15936 7142 15988 7148
rect 15948 6934 15976 7142
rect 16040 7002 16068 7414
rect 16132 7410 16160 8366
rect 16208 8358 16528 8382
rect 16208 8302 16220 8358
rect 16276 8302 16300 8358
rect 16356 8302 16380 8358
rect 16436 8302 16460 8358
rect 16516 8302 16528 8358
rect 16208 8278 16528 8302
rect 16208 8222 16220 8278
rect 16276 8222 16300 8278
rect 16356 8222 16380 8278
rect 16436 8222 16460 8278
rect 16516 8222 16528 8278
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16208 7642 16528 8222
rect 16592 8090 16620 8230
rect 16580 8084 16632 8090
rect 16580 8026 16632 8032
rect 16208 7590 16214 7642
rect 16266 7590 16278 7642
rect 16330 7590 16342 7642
rect 16394 7590 16406 7642
rect 16458 7590 16470 7642
rect 16522 7590 16528 7642
rect 16120 7404 16172 7410
rect 16120 7346 16172 7352
rect 16028 6996 16080 7002
rect 16028 6938 16080 6944
rect 15936 6928 15988 6934
rect 15936 6870 15988 6876
rect 16040 6780 16068 6938
rect 15948 6752 16068 6780
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15660 5840 15712 5846
rect 15660 5782 15712 5788
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15304 4236 15516 4264
rect 15304 4049 15332 4236
rect 15580 4214 15608 5306
rect 15672 4842 15700 5782
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15764 5166 15792 5714
rect 15752 5160 15804 5166
rect 15752 5102 15804 5108
rect 15672 4814 15792 4842
rect 15660 4684 15712 4690
rect 15660 4626 15712 4632
rect 15568 4208 15620 4214
rect 15396 4156 15568 4162
rect 15396 4150 15620 4156
rect 15396 4134 15608 4150
rect 15672 4146 15700 4626
rect 15290 4040 15346 4049
rect 15200 4004 15252 4010
rect 15290 3975 15346 3984
rect 15200 3946 15252 3952
rect 15304 3618 15332 3975
rect 15120 3590 15332 3618
rect 15120 3058 15148 3590
rect 15292 3528 15344 3534
rect 15292 3470 15344 3476
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15212 3058 15240 3334
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15016 2848 15068 2854
rect 15016 2790 15068 2796
rect 15304 2774 15332 3470
rect 15396 3398 15424 4134
rect 15580 4078 15608 4134
rect 15660 4140 15712 4146
rect 15660 4082 15712 4088
rect 15476 4072 15528 4078
rect 15476 4014 15528 4020
rect 15568 4072 15620 4078
rect 15764 4026 15792 4814
rect 15844 4480 15896 4486
rect 15844 4422 15896 4428
rect 15568 4014 15620 4020
rect 15384 3392 15436 3398
rect 15384 3334 15436 3340
rect 15212 2746 15332 2774
rect 14740 2508 14792 2514
rect 14740 2450 14792 2456
rect 14752 1970 14780 2450
rect 14280 1964 14332 1970
rect 14280 1906 14332 1912
rect 14740 1964 14792 1970
rect 14740 1906 14792 1912
rect 13820 1760 13872 1766
rect 13820 1702 13872 1708
rect 13832 1290 13860 1702
rect 14004 1352 14056 1358
rect 14004 1294 14056 1300
rect 13820 1284 13872 1290
rect 13820 1226 13872 1232
rect 14016 1222 14044 1294
rect 14292 1290 14320 1906
rect 14752 1426 14780 1906
rect 15212 1834 15240 2746
rect 15396 2514 15424 3334
rect 15488 3058 15516 4014
rect 15672 3998 15792 4026
rect 15672 3890 15700 3998
rect 15580 3862 15700 3890
rect 15752 3936 15804 3942
rect 15752 3878 15804 3884
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15384 2508 15436 2514
rect 15384 2450 15436 2456
rect 15488 2310 15516 2790
rect 15476 2304 15528 2310
rect 15476 2246 15528 2252
rect 15488 2038 15516 2246
rect 15476 2032 15528 2038
rect 15476 1974 15528 1980
rect 15580 1970 15608 3862
rect 15764 3534 15792 3878
rect 15856 3670 15884 4422
rect 15948 4282 15976 6752
rect 16208 6554 16528 7590
rect 16208 6502 16214 6554
rect 16266 6502 16278 6554
rect 16330 6502 16342 6554
rect 16394 6502 16406 6554
rect 16458 6502 16470 6554
rect 16522 6502 16528 6554
rect 16208 5466 16528 6502
rect 16684 6118 16712 8502
rect 16960 8430 16988 8978
rect 17236 8566 17264 9318
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16960 7342 16988 8366
rect 17500 7948 17552 7954
rect 17500 7890 17552 7896
rect 17132 7744 17184 7750
rect 17132 7686 17184 7692
rect 17408 7744 17460 7750
rect 17408 7686 17460 7692
rect 16948 7336 17000 7342
rect 16948 7278 17000 7284
rect 16960 6866 16988 7278
rect 16948 6860 17000 6866
rect 16948 6802 17000 6808
rect 17040 6860 17092 6866
rect 17040 6802 17092 6808
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16776 6458 16804 6666
rect 16764 6452 16816 6458
rect 16764 6394 16816 6400
rect 17052 6361 17080 6802
rect 17144 6633 17172 7686
rect 17420 7478 17448 7686
rect 17408 7472 17460 7478
rect 17408 7414 17460 7420
rect 17224 6656 17276 6662
rect 17130 6624 17186 6633
rect 17224 6598 17276 6604
rect 17130 6559 17186 6568
rect 17038 6352 17094 6361
rect 16948 6316 17000 6322
rect 17038 6287 17094 6296
rect 17144 6338 17172 6559
rect 17236 6458 17264 6598
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17144 6310 17264 6338
rect 16948 6258 17000 6264
rect 16856 6180 16908 6186
rect 16856 6122 16908 6128
rect 16672 6112 16724 6118
rect 16672 6054 16724 6060
rect 16578 5808 16634 5817
rect 16578 5743 16634 5752
rect 16592 5710 16620 5743
rect 16580 5704 16632 5710
rect 16684 5681 16712 6054
rect 16580 5646 16632 5652
rect 16670 5672 16726 5681
rect 16670 5607 16672 5616
rect 16724 5607 16726 5616
rect 16672 5578 16724 5584
rect 16208 5414 16214 5466
rect 16266 5414 16278 5466
rect 16330 5414 16342 5466
rect 16394 5414 16406 5466
rect 16458 5414 16470 5466
rect 16522 5414 16528 5466
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16132 4282 16160 5102
rect 16208 4378 16528 5414
rect 16868 5234 16896 6122
rect 16960 6118 16988 6258
rect 16948 6112 17000 6118
rect 17144 6066 17172 6310
rect 16948 6054 17000 6060
rect 17052 6038 17172 6066
rect 17052 5760 17080 6038
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 16960 5732 17080 5760
rect 16960 5642 16988 5732
rect 16948 5636 17000 5642
rect 16948 5578 17000 5584
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 16856 5228 16908 5234
rect 16856 5170 16908 5176
rect 16764 5160 16816 5166
rect 16764 5102 16816 5108
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 16208 4326 16214 4378
rect 16266 4326 16278 4378
rect 16330 4326 16342 4378
rect 16394 4326 16406 4378
rect 16458 4326 16470 4378
rect 16522 4326 16528 4378
rect 15936 4276 15988 4282
rect 15936 4218 15988 4224
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 15844 3664 15896 3670
rect 15844 3606 15896 3612
rect 15752 3528 15804 3534
rect 15804 3488 15884 3516
rect 15752 3470 15804 3476
rect 15752 2984 15804 2990
rect 15752 2926 15804 2932
rect 15764 2446 15792 2926
rect 15752 2440 15804 2446
rect 15752 2382 15804 2388
rect 15856 2394 15884 3488
rect 16028 3460 16080 3466
rect 16028 3402 16080 3408
rect 16040 3194 16068 3402
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 16026 3088 16082 3097
rect 16026 3023 16082 3032
rect 16040 2774 16068 3023
rect 16132 2990 16160 3878
rect 16208 3290 16528 4326
rect 16592 3534 16620 5034
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 16580 3528 16632 3534
rect 16580 3470 16632 3476
rect 16208 3238 16214 3290
rect 16266 3238 16278 3290
rect 16330 3238 16342 3290
rect 16394 3238 16406 3290
rect 16458 3238 16470 3290
rect 16522 3238 16528 3290
rect 16120 2984 16172 2990
rect 16120 2926 16172 2932
rect 16040 2746 16160 2774
rect 15934 2544 15990 2553
rect 15934 2479 15936 2488
rect 15988 2479 15990 2488
rect 15936 2450 15988 2456
rect 16028 2440 16080 2446
rect 15568 1964 15620 1970
rect 15568 1906 15620 1912
rect 15200 1828 15252 1834
rect 15200 1770 15252 1776
rect 15212 1426 15240 1770
rect 14740 1420 14792 1426
rect 14740 1362 14792 1368
rect 15200 1420 15252 1426
rect 15200 1362 15252 1368
rect 15764 1358 15792 2382
rect 15856 2378 15976 2394
rect 16028 2382 16080 2388
rect 15856 2372 15988 2378
rect 15856 2366 15936 2372
rect 15936 2314 15988 2320
rect 15936 1760 15988 1766
rect 15936 1702 15988 1708
rect 15948 1562 15976 1702
rect 15936 1556 15988 1562
rect 15936 1498 15988 1504
rect 16040 1494 16068 2382
rect 16028 1488 16080 1494
rect 16028 1430 16080 1436
rect 15752 1352 15804 1358
rect 15752 1294 15804 1300
rect 14280 1284 14332 1290
rect 14280 1226 14332 1232
rect 14004 1216 14056 1222
rect 14004 1158 14056 1164
rect 13728 944 13780 950
rect 13728 886 13780 892
rect 14016 800 14044 1158
rect 16132 800 16160 2746
rect 16208 2202 16528 3238
rect 16208 2150 16214 2202
rect 16266 2150 16278 2202
rect 16330 2150 16342 2202
rect 16394 2150 16406 2202
rect 16458 2150 16470 2202
rect 16522 2150 16528 2202
rect 16208 1114 16528 2150
rect 16592 2038 16620 3470
rect 16684 2514 16712 4966
rect 16776 4078 16804 5102
rect 17052 4214 17080 5510
rect 17040 4208 17092 4214
rect 17040 4150 17092 4156
rect 16764 4072 16816 4078
rect 16764 4014 16816 4020
rect 17040 4072 17092 4078
rect 17040 4014 17092 4020
rect 16672 2508 16724 2514
rect 16672 2450 16724 2456
rect 16580 2032 16632 2038
rect 16580 1974 16632 1980
rect 16776 1970 16804 4014
rect 17052 3738 17080 4014
rect 17040 3732 17092 3738
rect 17040 3674 17092 3680
rect 16948 3528 17000 3534
rect 16948 3470 17000 3476
rect 16856 3392 16908 3398
rect 16856 3334 16908 3340
rect 16868 3194 16896 3334
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 16856 3052 16908 3058
rect 16856 2994 16908 3000
rect 16868 2514 16896 2994
rect 16856 2508 16908 2514
rect 16856 2450 16908 2456
rect 16854 2408 16910 2417
rect 16854 2343 16910 2352
rect 16764 1964 16816 1970
rect 16764 1906 16816 1912
rect 16868 1290 16896 2343
rect 16960 1290 16988 3470
rect 17144 2961 17172 5850
rect 17236 5574 17264 6310
rect 17512 6254 17540 7890
rect 17604 7886 17632 10202
rect 17696 9926 17724 12038
rect 17972 10742 18000 12038
rect 18052 11144 18104 11150
rect 18052 11086 18104 11092
rect 17960 10736 18012 10742
rect 17960 10678 18012 10684
rect 18064 10266 18092 11086
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 18064 9178 18092 9590
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18052 9172 18104 9178
rect 18052 9114 18104 9120
rect 17684 8084 17736 8090
rect 17684 8026 17736 8032
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17604 6934 17632 7822
rect 17592 6928 17644 6934
rect 17592 6870 17644 6876
rect 17500 6248 17552 6254
rect 17500 6190 17552 6196
rect 17406 5944 17462 5953
rect 17406 5879 17462 5888
rect 17420 5846 17448 5879
rect 17408 5840 17460 5846
rect 17314 5808 17370 5817
rect 17408 5782 17460 5788
rect 17314 5743 17316 5752
rect 17368 5743 17370 5752
rect 17316 5714 17368 5720
rect 17406 5672 17462 5681
rect 17406 5607 17408 5616
rect 17460 5607 17462 5616
rect 17408 5578 17460 5584
rect 17224 5568 17276 5574
rect 17224 5510 17276 5516
rect 17236 3534 17264 5510
rect 17316 5160 17368 5166
rect 17316 5102 17368 5108
rect 17328 4826 17356 5102
rect 17316 4820 17368 4826
rect 17316 4762 17368 4768
rect 17224 3528 17276 3534
rect 17224 3470 17276 3476
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17224 2984 17276 2990
rect 17130 2952 17186 2961
rect 17224 2926 17276 2932
rect 17130 2887 17186 2896
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17052 2038 17080 2450
rect 17040 2032 17092 2038
rect 17040 1974 17092 1980
rect 17144 1562 17172 2887
rect 17236 2514 17264 2926
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 17132 1556 17184 1562
rect 17132 1498 17184 1504
rect 17328 1358 17356 2994
rect 17420 2417 17448 5578
rect 17512 4690 17540 6190
rect 17696 5914 17724 8026
rect 18248 7954 18276 9454
rect 18236 7948 18288 7954
rect 18236 7890 18288 7896
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 18064 7002 18092 7686
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17684 5908 17736 5914
rect 17684 5850 17736 5856
rect 17500 4684 17552 4690
rect 17500 4626 17552 4632
rect 17512 3058 17540 4626
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17604 3126 17632 4422
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17696 3194 17724 4218
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17592 3120 17644 3126
rect 17592 3062 17644 3068
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17604 2514 17632 3062
rect 17684 2848 17736 2854
rect 17684 2790 17736 2796
rect 17592 2508 17644 2514
rect 17592 2450 17644 2456
rect 17696 2446 17724 2790
rect 17788 2650 17816 6190
rect 17776 2644 17828 2650
rect 17776 2586 17828 2592
rect 17776 2508 17828 2514
rect 17776 2450 17828 2456
rect 17684 2440 17736 2446
rect 17406 2408 17462 2417
rect 17684 2382 17736 2388
rect 17406 2343 17462 2352
rect 17592 2372 17644 2378
rect 17592 2314 17644 2320
rect 17500 2032 17552 2038
rect 17420 1992 17500 2020
rect 17420 1562 17448 1992
rect 17500 1974 17552 1980
rect 17604 1562 17632 2314
rect 17408 1556 17460 1562
rect 17408 1498 17460 1504
rect 17592 1556 17644 1562
rect 17592 1498 17644 1504
rect 17408 1420 17460 1426
rect 17408 1362 17460 1368
rect 17316 1352 17368 1358
rect 17316 1294 17368 1300
rect 17420 1306 17448 1362
rect 17684 1352 17736 1358
rect 17420 1300 17684 1306
rect 17420 1294 17736 1300
rect 16856 1284 16908 1290
rect 16856 1226 16908 1232
rect 16948 1284 17000 1290
rect 17420 1278 17724 1294
rect 16948 1226 17000 1232
rect 16208 1062 16214 1114
rect 16266 1062 16278 1114
rect 16330 1062 16342 1114
rect 16394 1062 16406 1114
rect 16458 1062 16470 1114
rect 16522 1062 16528 1114
rect 16208 1040 16528 1062
rect 1306 0 1362 800
rect 3422 0 3478 800
rect 5538 0 5594 800
rect 7654 0 7710 800
rect 9770 0 9826 800
rect 11886 0 11942 800
rect 14002 0 14058 800
rect 16118 0 16174 800
rect 17696 746 17724 1278
rect 17788 1272 17816 2450
rect 17880 2106 17908 6394
rect 18064 6390 18092 6938
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18052 6384 18104 6390
rect 18052 6326 18104 6332
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 17972 5658 18000 6258
rect 18248 5710 18276 6734
rect 18340 5846 18368 12174
rect 18512 11824 18564 11830
rect 18512 11766 18564 11772
rect 18524 10266 18552 11766
rect 18800 10810 18828 15098
rect 19352 15026 19380 15506
rect 19524 15360 19576 15366
rect 19524 15302 19576 15308
rect 19432 15156 19484 15162
rect 19432 15098 19484 15104
rect 19340 15020 19392 15026
rect 19340 14962 19392 14968
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19352 14346 19380 14554
rect 19444 14482 19472 15098
rect 19536 15065 19564 15302
rect 19522 15056 19578 15065
rect 19628 15026 19656 17002
rect 19812 15978 19840 18022
rect 19996 16590 20024 18090
rect 20208 17978 20528 18544
rect 20628 18420 20680 18426
rect 20628 18362 20680 18368
rect 20904 18420 20956 18426
rect 20904 18362 20956 18368
rect 20208 17926 20214 17978
rect 20266 17926 20278 17978
rect 20330 17926 20342 17978
rect 20394 17926 20406 17978
rect 20458 17926 20470 17978
rect 20522 17926 20528 17978
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 20088 17270 20116 17478
rect 20076 17264 20128 17270
rect 20076 17206 20128 17212
rect 20208 16890 20528 17926
rect 20640 17814 20668 18362
rect 20812 18284 20864 18290
rect 20812 18226 20864 18232
rect 20628 17808 20680 17814
rect 20628 17750 20680 17756
rect 20824 17202 20852 18226
rect 20916 18222 20944 18362
rect 20904 18216 20956 18222
rect 20904 18158 20956 18164
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 21364 17128 21416 17134
rect 21364 17070 21416 17076
rect 20904 16992 20956 16998
rect 20904 16934 20956 16940
rect 20208 16838 20214 16890
rect 20266 16838 20278 16890
rect 20330 16838 20342 16890
rect 20394 16838 20406 16890
rect 20458 16838 20470 16890
rect 20522 16838 20528 16890
rect 19984 16584 20036 16590
rect 19984 16526 20036 16532
rect 19892 16040 19944 16046
rect 19892 15982 19944 15988
rect 19800 15972 19852 15978
rect 19800 15914 19852 15920
rect 19904 15586 19932 15982
rect 19984 15904 20036 15910
rect 19984 15846 20036 15852
rect 19812 15558 19932 15586
rect 19708 15156 19760 15162
rect 19708 15098 19760 15104
rect 19522 14991 19578 15000
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19628 14618 19656 14962
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19432 14476 19484 14482
rect 19432 14418 19484 14424
rect 19340 14340 19392 14346
rect 19340 14282 19392 14288
rect 19352 13938 19380 14282
rect 19432 14000 19484 14006
rect 19432 13942 19484 13948
rect 19340 13932 19392 13938
rect 19340 13874 19392 13880
rect 19444 13462 19472 13942
rect 19432 13456 19484 13462
rect 19432 13398 19484 13404
rect 19720 13394 19748 15098
rect 19708 13388 19760 13394
rect 19708 13330 19760 13336
rect 19340 13320 19392 13326
rect 18878 13288 18934 13297
rect 19340 13262 19392 13268
rect 18878 13223 18880 13232
rect 18932 13223 18934 13232
rect 18880 13194 18932 13200
rect 19352 12238 19380 13262
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19352 11762 19380 12174
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19444 11626 19472 12106
rect 19432 11620 19484 11626
rect 19432 11562 19484 11568
rect 19720 11286 19748 13330
rect 19812 12646 19840 15558
rect 19892 15496 19944 15502
rect 19892 15438 19944 15444
rect 19904 15026 19932 15438
rect 19996 15366 20024 15846
rect 20208 15802 20528 16838
rect 20916 16794 20944 16934
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 21180 16584 21232 16590
rect 21180 16526 21232 16532
rect 20208 15750 20214 15802
rect 20266 15750 20278 15802
rect 20330 15750 20342 15802
rect 20394 15750 20406 15802
rect 20458 15750 20470 15802
rect 20522 15750 20528 15802
rect 19984 15360 20036 15366
rect 19984 15302 20036 15308
rect 19892 15020 19944 15026
rect 19892 14962 19944 14968
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19812 12306 19840 12582
rect 19800 12300 19852 12306
rect 19800 12242 19852 12248
rect 19812 11694 19840 12242
rect 19904 12073 19932 14962
rect 19996 13938 20024 15302
rect 20208 14714 20528 15750
rect 20640 15706 20668 16526
rect 20720 16108 20772 16114
rect 20720 16050 20772 16056
rect 20996 16108 21048 16114
rect 20996 16050 21048 16056
rect 20628 15700 20680 15706
rect 20628 15642 20680 15648
rect 20628 15428 20680 15434
rect 20628 15370 20680 15376
rect 20640 15162 20668 15370
rect 20628 15156 20680 15162
rect 20628 15098 20680 15104
rect 20626 15056 20682 15065
rect 20732 15042 20760 16050
rect 21008 15910 21036 16050
rect 20996 15904 21048 15910
rect 20996 15846 21048 15852
rect 20904 15496 20956 15502
rect 20904 15438 20956 15444
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20682 15014 20760 15042
rect 20626 14991 20628 15000
rect 20680 14991 20682 15000
rect 20628 14962 20680 14968
rect 20208 14662 20214 14714
rect 20266 14662 20278 14714
rect 20330 14662 20342 14714
rect 20394 14662 20406 14714
rect 20458 14662 20470 14714
rect 20522 14662 20528 14714
rect 20076 14272 20128 14278
rect 20076 14214 20128 14220
rect 19984 13932 20036 13938
rect 19984 13874 20036 13880
rect 20088 13394 20116 14214
rect 20208 13626 20528 14662
rect 20628 14408 20680 14414
rect 20628 14350 20680 14356
rect 20640 13734 20668 14350
rect 20628 13728 20680 13734
rect 20628 13670 20680 13676
rect 20208 13574 20214 13626
rect 20266 13574 20278 13626
rect 20330 13574 20342 13626
rect 20394 13574 20406 13626
rect 20458 13574 20470 13626
rect 20522 13574 20528 13626
rect 20076 13388 20128 13394
rect 20076 13330 20128 13336
rect 19984 13252 20036 13258
rect 19984 13194 20036 13200
rect 19996 12238 20024 13194
rect 20208 12538 20528 13574
rect 20640 12850 20668 13670
rect 20732 13376 20760 15014
rect 20824 14074 20852 15302
rect 20916 15201 20944 15438
rect 20902 15192 20958 15201
rect 20902 15127 20958 15136
rect 20904 15088 20956 15094
rect 20904 15030 20956 15036
rect 20812 14068 20864 14074
rect 20812 14010 20864 14016
rect 20732 13348 20852 13376
rect 20720 13252 20772 13258
rect 20720 13194 20772 13200
rect 20628 12844 20680 12850
rect 20628 12786 20680 12792
rect 20208 12486 20214 12538
rect 20266 12518 20278 12538
rect 20330 12518 20342 12538
rect 20394 12518 20406 12538
rect 20458 12518 20470 12538
rect 20276 12486 20278 12518
rect 20458 12486 20460 12518
rect 20522 12486 20528 12538
rect 20208 12462 20220 12486
rect 20276 12462 20300 12486
rect 20356 12462 20380 12486
rect 20436 12462 20460 12486
rect 20516 12462 20528 12486
rect 20208 12438 20528 12462
rect 20208 12382 20220 12438
rect 20276 12382 20300 12438
rect 20356 12382 20380 12438
rect 20436 12382 20460 12438
rect 20516 12382 20528 12438
rect 20076 12368 20128 12374
rect 20076 12310 20128 12316
rect 20208 12358 20528 12382
rect 19984 12232 20036 12238
rect 19984 12174 20036 12180
rect 19890 12064 19946 12073
rect 19890 11999 19946 12008
rect 19800 11688 19852 11694
rect 19800 11630 19852 11636
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19904 11150 19932 11999
rect 19996 11898 20024 12174
rect 20088 11898 20116 12310
rect 20208 12302 20220 12358
rect 20276 12302 20300 12358
rect 20356 12302 20380 12358
rect 20436 12302 20460 12358
rect 20516 12302 20528 12358
rect 20208 12278 20528 12302
rect 20208 12222 20220 12278
rect 20276 12222 20300 12278
rect 20356 12222 20380 12278
rect 20436 12222 20460 12278
rect 20516 12222 20528 12278
rect 20640 12238 20668 12786
rect 19984 11892 20036 11898
rect 19984 11834 20036 11840
rect 20076 11892 20128 11898
rect 20076 11834 20128 11840
rect 20082 11688 20134 11694
rect 20074 11656 20082 11665
rect 20130 11630 20134 11636
rect 20074 11591 20130 11600
rect 20208 11450 20528 12222
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 20628 12096 20680 12102
rect 20628 12038 20680 12044
rect 20208 11398 20214 11450
rect 20266 11398 20278 11450
rect 20330 11398 20342 11450
rect 20394 11398 20406 11450
rect 20458 11398 20470 11450
rect 20522 11398 20528 11450
rect 19892 11144 19944 11150
rect 19812 11104 19892 11132
rect 18788 10804 18840 10810
rect 18788 10746 18840 10752
rect 18512 10260 18564 10266
rect 18512 10202 18564 10208
rect 19812 9994 19840 11104
rect 19892 11086 19944 11092
rect 20208 10362 20528 11398
rect 20640 11286 20668 12038
rect 20732 11762 20760 13194
rect 20824 11830 20852 13348
rect 20812 11824 20864 11830
rect 20812 11766 20864 11772
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20824 11665 20852 11766
rect 20810 11656 20866 11665
rect 20810 11591 20866 11600
rect 20628 11280 20680 11286
rect 20628 11222 20680 11228
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20640 10810 20668 11086
rect 20628 10804 20680 10810
rect 20628 10746 20680 10752
rect 20208 10310 20214 10362
rect 20266 10310 20278 10362
rect 20330 10310 20342 10362
rect 20394 10310 20406 10362
rect 20458 10310 20470 10362
rect 20522 10310 20528 10362
rect 19892 10124 19944 10130
rect 19892 10066 19944 10072
rect 19800 9988 19852 9994
rect 19800 9930 19852 9936
rect 19616 9920 19668 9926
rect 19616 9862 19668 9868
rect 18604 9648 18656 9654
rect 18604 9590 18656 9596
rect 18616 8838 18644 9590
rect 18696 9580 18748 9586
rect 18696 9522 18748 9528
rect 18880 9580 18932 9586
rect 18880 9522 18932 9528
rect 19340 9580 19392 9586
rect 19340 9522 19392 9528
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18616 7936 18644 8774
rect 18708 8634 18736 9522
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18696 8628 18748 8634
rect 18696 8570 18748 8576
rect 18800 8566 18828 9318
rect 18892 8906 18920 9522
rect 18972 9376 19024 9382
rect 18972 9318 19024 9324
rect 18984 9178 19012 9318
rect 18972 9172 19024 9178
rect 18972 9114 19024 9120
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18788 8560 18840 8566
rect 18788 8502 18840 8508
rect 18788 8356 18840 8362
rect 18788 8298 18840 8304
rect 18696 7948 18748 7954
rect 18616 7908 18696 7936
rect 18696 7890 18748 7896
rect 18708 7818 18736 7890
rect 18696 7812 18748 7818
rect 18696 7754 18748 7760
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18524 7410 18552 7686
rect 18512 7404 18564 7410
rect 18512 7346 18564 7352
rect 18420 6656 18472 6662
rect 18418 6624 18420 6633
rect 18472 6624 18474 6633
rect 18418 6559 18474 6568
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18236 5704 18288 5710
rect 18234 5672 18236 5681
rect 18288 5672 18290 5681
rect 17972 5630 18092 5658
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17972 5302 18000 5510
rect 17960 5296 18012 5302
rect 17960 5238 18012 5244
rect 18064 3097 18092 5630
rect 18234 5607 18290 5616
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 18248 3466 18276 3878
rect 18524 3738 18552 6258
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18708 4622 18736 5306
rect 18696 4616 18748 4622
rect 18696 4558 18748 4564
rect 18512 3732 18564 3738
rect 18512 3674 18564 3680
rect 18800 3466 18828 8298
rect 18892 8294 18920 8842
rect 18880 8288 18932 8294
rect 18880 8230 18932 8236
rect 18892 7818 18920 8230
rect 18984 8090 19012 9114
rect 19352 9042 19380 9522
rect 19628 9042 19656 9862
rect 19812 9178 19840 9930
rect 19800 9172 19852 9178
rect 19800 9114 19852 9120
rect 19340 9036 19392 9042
rect 19340 8978 19392 8984
rect 19616 9036 19668 9042
rect 19616 8978 19668 8984
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19352 8634 19380 8842
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 18972 8084 19024 8090
rect 18972 8026 19024 8032
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 18880 7812 18932 7818
rect 18880 7754 18932 7760
rect 18892 6798 18920 7754
rect 18984 7002 19012 8026
rect 19432 7744 19484 7750
rect 19432 7686 19484 7692
rect 19444 7478 19472 7686
rect 19340 7472 19392 7478
rect 19340 7414 19392 7420
rect 19432 7472 19484 7478
rect 19432 7414 19484 7420
rect 19352 7324 19380 7414
rect 19352 7296 19472 7324
rect 19248 7200 19300 7206
rect 19248 7142 19300 7148
rect 18972 6996 19024 7002
rect 18972 6938 19024 6944
rect 19260 6882 19288 7142
rect 19260 6854 19380 6882
rect 19352 6798 19380 6854
rect 18880 6792 18932 6798
rect 18880 6734 18932 6740
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 18972 6656 19024 6662
rect 18972 6598 19024 6604
rect 18984 6186 19012 6598
rect 19064 6248 19116 6254
rect 19064 6190 19116 6196
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 18972 6180 19024 6186
rect 18972 6122 19024 6128
rect 19076 5370 19104 6190
rect 19352 6118 19380 6190
rect 19340 6112 19392 6118
rect 19340 6054 19392 6060
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 19156 5568 19208 5574
rect 19156 5510 19208 5516
rect 19064 5364 19116 5370
rect 19064 5306 19116 5312
rect 18880 4616 18932 4622
rect 18880 4558 18932 4564
rect 18892 4214 18920 4558
rect 18880 4208 18932 4214
rect 18880 4150 18932 4156
rect 18880 4072 18932 4078
rect 18880 4014 18932 4020
rect 18236 3460 18288 3466
rect 18236 3402 18288 3408
rect 18696 3460 18748 3466
rect 18696 3402 18748 3408
rect 18788 3460 18840 3466
rect 18788 3402 18840 3408
rect 18604 3392 18656 3398
rect 18604 3334 18656 3340
rect 18616 3126 18644 3334
rect 18708 3194 18736 3402
rect 18696 3188 18748 3194
rect 18696 3130 18748 3136
rect 18512 3120 18564 3126
rect 18050 3088 18106 3097
rect 18512 3062 18564 3068
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18050 3023 18106 3032
rect 18236 2848 18288 2854
rect 18236 2790 18288 2796
rect 18142 2680 18198 2689
rect 17960 2644 18012 2650
rect 18142 2615 18198 2624
rect 17960 2586 18012 2592
rect 17972 2553 18000 2586
rect 17958 2544 18014 2553
rect 17958 2479 18014 2488
rect 18156 2446 18184 2615
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 17868 2100 17920 2106
rect 17868 2042 17920 2048
rect 18156 1834 18184 2382
rect 18144 1828 18196 1834
rect 18144 1770 18196 1776
rect 18248 1562 18276 2790
rect 18420 2032 18472 2038
rect 18420 1974 18472 1980
rect 18236 1556 18288 1562
rect 18236 1498 18288 1504
rect 17868 1284 17920 1290
rect 17788 1244 17868 1272
rect 17868 1226 17920 1232
rect 18432 1222 18460 1974
rect 18420 1216 18472 1222
rect 18420 1158 18472 1164
rect 18524 1018 18552 3062
rect 18786 2816 18842 2825
rect 18786 2751 18842 2760
rect 18800 2650 18828 2751
rect 18788 2644 18840 2650
rect 18788 2586 18840 2592
rect 18696 2576 18748 2582
rect 18696 2518 18748 2524
rect 18708 2106 18736 2518
rect 18892 2496 18920 4014
rect 18972 4004 19024 4010
rect 18972 3946 19024 3952
rect 18984 3194 19012 3946
rect 19064 3664 19116 3670
rect 19064 3606 19116 3612
rect 18972 3188 19024 3194
rect 18972 3130 19024 3136
rect 18984 2854 19012 3130
rect 18972 2848 19024 2854
rect 19076 2825 19104 3606
rect 18972 2790 19024 2796
rect 19062 2816 19118 2825
rect 19062 2751 19118 2760
rect 18892 2468 19104 2496
rect 18972 2372 19024 2378
rect 18972 2314 19024 2320
rect 18696 2100 18748 2106
rect 18696 2042 18748 2048
rect 18708 1358 18736 2042
rect 18788 1896 18840 1902
rect 18788 1838 18840 1844
rect 18800 1562 18828 1838
rect 18788 1556 18840 1562
rect 18788 1498 18840 1504
rect 18984 1358 19012 2314
rect 19076 2106 19104 2468
rect 19064 2100 19116 2106
rect 19064 2042 19116 2048
rect 18696 1352 18748 1358
rect 18696 1294 18748 1300
rect 18972 1352 19024 1358
rect 18972 1294 19024 1300
rect 19076 1222 19104 2042
rect 19168 1340 19196 5510
rect 19260 3534 19288 5646
rect 19340 4548 19392 4554
rect 19340 4490 19392 4496
rect 19352 4214 19380 4490
rect 19340 4208 19392 4214
rect 19340 4150 19392 4156
rect 19444 3534 19472 7296
rect 19536 6934 19564 8026
rect 19628 8022 19656 8978
rect 19708 8832 19760 8838
rect 19708 8774 19760 8780
rect 19720 8634 19748 8774
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19708 8424 19760 8430
rect 19708 8366 19760 8372
rect 19616 8016 19668 8022
rect 19616 7958 19668 7964
rect 19628 7002 19656 7958
rect 19720 7954 19748 8366
rect 19812 8242 19840 9114
rect 19904 8430 19932 10066
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19996 9518 20024 9862
rect 19984 9512 20036 9518
rect 19984 9454 20036 9460
rect 20208 9274 20528 10310
rect 20628 10056 20680 10062
rect 20628 9998 20680 10004
rect 20208 9222 20214 9274
rect 20266 9222 20278 9274
rect 20330 9222 20342 9274
rect 20394 9222 20406 9274
rect 20458 9222 20470 9274
rect 20522 9222 20528 9274
rect 20076 8900 20128 8906
rect 20076 8842 20128 8848
rect 20088 8634 20116 8842
rect 20076 8628 20128 8634
rect 20076 8570 20128 8576
rect 19892 8424 19944 8430
rect 19892 8366 19944 8372
rect 19812 8214 19932 8242
rect 19708 7948 19760 7954
rect 19708 7890 19760 7896
rect 19616 6996 19668 7002
rect 19616 6938 19668 6944
rect 19524 6928 19576 6934
rect 19576 6876 19656 6882
rect 19524 6870 19656 6876
rect 19536 6854 19656 6870
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5302 19564 6054
rect 19628 5914 19656 6854
rect 19720 6322 19748 7890
rect 19800 7744 19852 7750
rect 19800 7686 19852 7692
rect 19812 7546 19840 7686
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19904 7426 19932 8214
rect 20208 8186 20528 9222
rect 20640 8838 20668 9998
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20208 8134 20214 8186
rect 20266 8134 20278 8186
rect 20330 8134 20342 8186
rect 20394 8134 20406 8186
rect 20458 8134 20470 8186
rect 20522 8134 20528 8186
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19812 7398 19932 7426
rect 19708 6316 19760 6322
rect 19708 6258 19760 6264
rect 19812 6254 19840 7398
rect 20088 7002 20116 7686
rect 20208 7098 20528 8134
rect 20916 7834 20944 15030
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21008 12986 21036 14962
rect 21100 14618 21128 16526
rect 21192 16454 21220 16526
rect 21272 16516 21324 16522
rect 21272 16458 21324 16464
rect 21180 16448 21232 16454
rect 21180 16390 21232 16396
rect 21192 16114 21220 16390
rect 21284 16250 21312 16458
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 21180 16108 21232 16114
rect 21232 16068 21312 16096
rect 21180 16050 21232 16056
rect 21180 15904 21232 15910
rect 21180 15846 21232 15852
rect 21192 15570 21220 15846
rect 21180 15564 21232 15570
rect 21180 15506 21232 15512
rect 21192 15026 21220 15506
rect 21284 15065 21312 16068
rect 21270 15056 21326 15065
rect 21180 15020 21232 15026
rect 21270 14991 21272 15000
rect 21180 14962 21232 14968
rect 21324 14991 21326 15000
rect 21272 14962 21324 14968
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21100 14074 21128 14350
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20996 12980 21048 12986
rect 20996 12922 21048 12928
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 21100 12238 21128 12786
rect 20996 12232 21048 12238
rect 20996 12174 21048 12180
rect 21088 12232 21140 12238
rect 21088 12174 21140 12180
rect 21008 11898 21036 12174
rect 20996 11892 21048 11898
rect 20996 11834 21048 11840
rect 21100 11694 21128 12174
rect 21088 11688 21140 11694
rect 21088 11630 21140 11636
rect 20996 11144 21048 11150
rect 21100 11132 21128 11630
rect 21192 11286 21220 14962
rect 21284 13190 21312 14962
rect 21376 14618 21404 17070
rect 21468 16114 21496 18634
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21640 18080 21692 18086
rect 21640 18022 21692 18028
rect 21652 17678 21680 18022
rect 21836 17678 21864 18090
rect 21640 17672 21692 17678
rect 21640 17614 21692 17620
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21548 16584 21600 16590
rect 21548 16526 21600 16532
rect 21456 16108 21508 16114
rect 21456 16050 21508 16056
rect 21456 15904 21508 15910
rect 21456 15846 21508 15852
rect 21468 15502 21496 15846
rect 21456 15496 21508 15502
rect 21456 15438 21508 15444
rect 21454 15192 21510 15201
rect 21454 15127 21510 15136
rect 21468 14906 21496 15127
rect 21560 15026 21588 16526
rect 21732 16516 21784 16522
rect 21732 16458 21784 16464
rect 21744 16182 21772 16458
rect 21732 16176 21784 16182
rect 21732 16118 21784 16124
rect 21732 15564 21784 15570
rect 21732 15506 21784 15512
rect 21640 15496 21692 15502
rect 21640 15438 21692 15444
rect 21548 15020 21600 15026
rect 21548 14962 21600 14968
rect 21468 14878 21588 14906
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21560 13802 21588 14878
rect 21548 13796 21600 13802
rect 21548 13738 21600 13744
rect 21456 13728 21508 13734
rect 21456 13670 21508 13676
rect 21468 13394 21496 13670
rect 21456 13388 21508 13394
rect 21456 13330 21508 13336
rect 21272 13184 21324 13190
rect 21272 13126 21324 13132
rect 21560 12986 21588 13738
rect 21548 12980 21600 12986
rect 21548 12922 21600 12928
rect 21456 12912 21508 12918
rect 21456 12854 21508 12860
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 21284 11558 21312 12718
rect 21364 12708 21416 12714
rect 21364 12650 21416 12656
rect 21376 11694 21404 12650
rect 21468 12442 21496 12854
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21468 11762 21496 12174
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21364 11688 21416 11694
rect 21364 11630 21416 11636
rect 21272 11552 21324 11558
rect 21272 11494 21324 11500
rect 21180 11280 21232 11286
rect 21180 11222 21232 11228
rect 21048 11104 21128 11132
rect 20996 11086 21048 11092
rect 21468 10810 21496 11698
rect 21560 11558 21588 12922
rect 21652 12850 21680 15438
rect 21744 15094 21772 15506
rect 21732 15088 21784 15094
rect 21732 15030 21784 15036
rect 21928 14074 21956 19200
rect 24412 19122 24440 19246
rect 24490 19200 24546 20000
rect 24504 19122 24532 19200
rect 24412 19094 24532 19122
rect 23480 18624 23532 18630
rect 23478 18592 23480 18601
rect 23532 18592 23534 18601
rect 23478 18527 23534 18536
rect 24208 18522 24528 18544
rect 24208 18470 24214 18522
rect 24266 18470 24278 18522
rect 24330 18470 24342 18522
rect 24394 18470 24406 18522
rect 24458 18470 24470 18522
rect 24522 18470 24528 18522
rect 23664 18352 23716 18358
rect 23664 18294 23716 18300
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 22468 18216 22520 18222
rect 22468 18158 22520 18164
rect 22480 17882 22508 18158
rect 23204 18080 23256 18086
rect 23204 18022 23256 18028
rect 23388 18080 23440 18086
rect 23388 18022 23440 18028
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 23216 17814 23244 18022
rect 23204 17808 23256 17814
rect 23204 17750 23256 17756
rect 23296 17672 23348 17678
rect 23296 17614 23348 17620
rect 22192 17196 22244 17202
rect 22192 17138 22244 17144
rect 22204 16114 22232 17138
rect 22468 17128 22520 17134
rect 22468 17070 22520 17076
rect 22928 17128 22980 17134
rect 22928 17070 22980 17076
rect 22284 17060 22336 17066
rect 22284 17002 22336 17008
rect 22296 16182 22324 17002
rect 22480 16590 22508 17070
rect 22376 16584 22428 16590
rect 22376 16526 22428 16532
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22284 16176 22336 16182
rect 22284 16118 22336 16124
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22100 15496 22152 15502
rect 22100 15438 22152 15444
rect 22008 15360 22060 15366
rect 22008 15302 22060 15308
rect 22020 15042 22048 15302
rect 22112 15162 22140 15438
rect 22204 15162 22232 16050
rect 22388 15178 22416 16526
rect 22480 15638 22508 16526
rect 22468 15632 22520 15638
rect 22468 15574 22520 15580
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22192 15156 22244 15162
rect 22388 15150 22508 15178
rect 22192 15098 22244 15104
rect 22282 15056 22338 15065
rect 22020 15026 22140 15042
rect 22020 15020 22152 15026
rect 22020 15014 22100 15020
rect 22282 14991 22284 15000
rect 22100 14962 22152 14968
rect 22336 14991 22338 15000
rect 22376 15020 22428 15026
rect 22284 14962 22336 14968
rect 22376 14962 22428 14968
rect 22284 14884 22336 14890
rect 22284 14826 22336 14832
rect 22296 14414 22324 14826
rect 22284 14408 22336 14414
rect 22284 14350 22336 14356
rect 21916 14068 21968 14074
rect 21916 14010 21968 14016
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22192 13932 22244 13938
rect 22192 13874 22244 13880
rect 22112 12850 22140 13874
rect 22204 13462 22232 13874
rect 22192 13456 22244 13462
rect 22192 13398 22244 13404
rect 22192 13184 22244 13190
rect 22192 13126 22244 13132
rect 21640 12844 21692 12850
rect 21640 12786 21692 12792
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22100 12300 22152 12306
rect 22100 12242 22152 12248
rect 21916 12232 21968 12238
rect 21916 12174 21968 12180
rect 21928 12073 21956 12174
rect 21914 12064 21970 12073
rect 21914 11999 21970 12008
rect 22112 11830 22140 12242
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21744 11150 21772 11766
rect 22112 11286 22140 11766
rect 22204 11762 22232 13126
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22204 11626 22232 11698
rect 22192 11620 22244 11626
rect 22192 11562 22244 11568
rect 22008 11280 22060 11286
rect 22008 11222 22060 11228
rect 22100 11280 22152 11286
rect 22100 11222 22152 11228
rect 21732 11144 21784 11150
rect 21732 11086 21784 11092
rect 21456 10804 21508 10810
rect 21456 10746 21508 10752
rect 21548 10600 21600 10606
rect 21548 10542 21600 10548
rect 21560 9994 21588 10542
rect 21916 10464 21968 10470
rect 21916 10406 21968 10412
rect 21928 9994 21956 10406
rect 22020 10010 22048 11222
rect 22204 11014 22232 11562
rect 22192 11008 22244 11014
rect 22192 10950 22244 10956
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21916 9988 21968 9994
rect 22020 9982 22140 10010
rect 21916 9930 21968 9936
rect 21364 9580 21416 9586
rect 21364 9522 21416 9528
rect 21272 8832 21324 8838
rect 21272 8774 21324 8780
rect 20996 8560 21048 8566
rect 20996 8502 21048 8508
rect 21008 8362 21036 8502
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 20996 8356 21048 8362
rect 20996 8298 21048 8304
rect 20812 7812 20864 7818
rect 20916 7806 21036 7834
rect 20812 7754 20864 7760
rect 20824 7546 20852 7754
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 20208 7046 20214 7098
rect 20266 7046 20278 7098
rect 20330 7046 20342 7098
rect 20394 7046 20406 7098
rect 20458 7046 20470 7098
rect 20522 7046 20528 7098
rect 20076 6996 20128 7002
rect 20076 6938 20128 6944
rect 19984 6792 20036 6798
rect 19984 6734 20036 6740
rect 19892 6724 19944 6730
rect 19892 6666 19944 6672
rect 19800 6248 19852 6254
rect 19800 6190 19852 6196
rect 19616 5908 19668 5914
rect 19616 5850 19668 5856
rect 19800 5704 19852 5710
rect 19800 5646 19852 5652
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19708 5296 19760 5302
rect 19708 5238 19760 5244
rect 19720 4826 19748 5238
rect 19708 4820 19760 4826
rect 19708 4762 19760 4768
rect 19614 4720 19670 4729
rect 19812 4706 19840 5646
rect 19614 4655 19616 4664
rect 19668 4655 19670 4664
rect 19720 4678 19840 4706
rect 19616 4626 19668 4632
rect 19616 4548 19668 4554
rect 19616 4490 19668 4496
rect 19628 4282 19656 4490
rect 19616 4276 19668 4282
rect 19616 4218 19668 4224
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19260 2446 19288 3470
rect 19340 3052 19392 3058
rect 19340 2994 19392 3000
rect 19352 2961 19380 2994
rect 19338 2952 19394 2961
rect 19338 2887 19394 2896
rect 19616 2916 19668 2922
rect 19616 2858 19668 2864
rect 19524 2848 19576 2854
rect 19524 2790 19576 2796
rect 19536 2514 19564 2790
rect 19524 2508 19576 2514
rect 19524 2450 19576 2456
rect 19628 2446 19656 2858
rect 19248 2440 19300 2446
rect 19248 2382 19300 2388
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19340 1352 19392 1358
rect 19168 1312 19340 1340
rect 19340 1294 19392 1300
rect 19064 1216 19116 1222
rect 19064 1158 19116 1164
rect 18512 1012 18564 1018
rect 18512 954 18564 960
rect 18236 944 18288 950
rect 18236 886 18288 892
rect 18248 800 18276 886
rect 19352 882 19380 1294
rect 19340 876 19392 882
rect 19340 818 19392 824
rect 17684 740 17736 746
rect 17684 682 17736 688
rect 18234 0 18290 800
rect 19352 746 19380 818
rect 19720 814 19748 4678
rect 19800 4616 19852 4622
rect 19800 4558 19852 4564
rect 19812 3942 19840 4558
rect 19800 3936 19852 3942
rect 19800 3878 19852 3884
rect 19904 3738 19932 6666
rect 19996 5166 20024 6734
rect 20076 6656 20128 6662
rect 20076 6598 20128 6604
rect 20088 5914 20116 6598
rect 20208 6010 20528 7046
rect 20916 7002 20944 7686
rect 20904 6996 20956 7002
rect 20904 6938 20956 6944
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20208 5958 20214 6010
rect 20266 5958 20278 6010
rect 20330 5958 20342 6010
rect 20394 5958 20406 6010
rect 20458 5958 20470 6010
rect 20522 5958 20528 6010
rect 20076 5908 20128 5914
rect 20076 5850 20128 5856
rect 20088 5778 20116 5850
rect 20076 5772 20128 5778
rect 20076 5714 20128 5720
rect 19984 5160 20036 5166
rect 19984 5102 20036 5108
rect 19996 4622 20024 5102
rect 20208 4922 20528 5958
rect 20628 5908 20680 5914
rect 20628 5850 20680 5856
rect 20208 4870 20214 4922
rect 20266 4870 20278 4922
rect 20330 4870 20342 4922
rect 20394 4870 20406 4922
rect 20458 4870 20470 4922
rect 20522 4870 20528 4922
rect 19984 4616 20036 4622
rect 19984 4558 20036 4564
rect 19996 4010 20024 4558
rect 20208 4518 20528 4870
rect 20076 4480 20128 4486
rect 20076 4422 20128 4428
rect 20208 4462 20220 4518
rect 20276 4462 20300 4518
rect 20356 4462 20380 4518
rect 20436 4462 20460 4518
rect 20516 4462 20528 4518
rect 20208 4438 20528 4462
rect 20088 4282 20116 4422
rect 20208 4382 20220 4438
rect 20276 4382 20300 4438
rect 20356 4382 20380 4438
rect 20436 4382 20460 4438
rect 20516 4382 20528 4438
rect 20208 4358 20528 4382
rect 20208 4302 20220 4358
rect 20276 4302 20300 4358
rect 20356 4302 20380 4358
rect 20436 4302 20460 4358
rect 20516 4302 20528 4358
rect 20076 4276 20128 4282
rect 20076 4218 20128 4224
rect 20208 4278 20528 4302
rect 20208 4222 20220 4278
rect 20276 4222 20300 4278
rect 20356 4222 20380 4278
rect 20436 4222 20460 4278
rect 20516 4222 20528 4278
rect 19984 4004 20036 4010
rect 19984 3946 20036 3952
rect 19892 3732 19944 3738
rect 19892 3674 19944 3680
rect 19800 3052 19852 3058
rect 19800 2994 19852 3000
rect 19812 1766 19840 2994
rect 19904 1902 19932 3674
rect 19996 3602 20024 3946
rect 20208 3834 20528 4222
rect 20208 3782 20214 3834
rect 20266 3782 20278 3834
rect 20330 3782 20342 3834
rect 20394 3782 20406 3834
rect 20458 3782 20470 3834
rect 20522 3782 20528 3834
rect 19984 3596 20036 3602
rect 19984 3538 20036 3544
rect 19996 3126 20024 3538
rect 20076 3528 20128 3534
rect 20076 3470 20128 3476
rect 19984 3120 20036 3126
rect 19984 3062 20036 3068
rect 20088 2650 20116 3470
rect 20208 2746 20528 3782
rect 20640 3754 20668 5850
rect 20732 5370 20760 6394
rect 20812 6316 20864 6322
rect 20812 6258 20864 6264
rect 20720 5364 20772 5370
rect 20720 5306 20772 5312
rect 20720 5024 20772 5030
rect 20720 4966 20772 4972
rect 20732 4826 20760 4966
rect 20720 4820 20772 4826
rect 20720 4762 20772 4768
rect 20720 4548 20772 4554
rect 20824 4536 20852 6258
rect 21008 5914 21036 7806
rect 21100 6390 21128 8434
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21192 8090 21220 8230
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 20904 5636 20956 5642
rect 20904 5578 20956 5584
rect 20916 5370 20944 5578
rect 21100 5574 21128 6326
rect 21192 6118 21220 8026
rect 21180 6112 21232 6118
rect 21180 6054 21232 6060
rect 21088 5568 21140 5574
rect 21088 5510 21140 5516
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 20824 4508 20944 4536
rect 20720 4490 20772 4496
rect 20732 3942 20760 4490
rect 20812 4140 20864 4146
rect 20812 4082 20864 4088
rect 20720 3936 20772 3942
rect 20720 3878 20772 3884
rect 20640 3726 20760 3754
rect 20732 3670 20760 3726
rect 20720 3664 20772 3670
rect 20720 3606 20772 3612
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20640 2990 20668 3334
rect 20824 3074 20852 4082
rect 20732 3046 20852 3074
rect 20628 2984 20680 2990
rect 20628 2926 20680 2932
rect 20208 2694 20214 2746
rect 20266 2694 20278 2746
rect 20330 2694 20342 2746
rect 20394 2694 20406 2746
rect 20458 2694 20470 2746
rect 20522 2694 20528 2746
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20076 2304 20128 2310
rect 20076 2246 20128 2252
rect 19892 1896 19944 1902
rect 19892 1838 19944 1844
rect 19984 1896 20036 1902
rect 19984 1838 20036 1844
rect 19800 1760 19852 1766
rect 19800 1702 19852 1708
rect 19812 1426 19840 1702
rect 19800 1420 19852 1426
rect 19800 1362 19852 1368
rect 19996 1222 20024 1838
rect 20088 1562 20116 2246
rect 20208 1658 20528 2694
rect 20628 2440 20680 2446
rect 20628 2382 20680 2388
rect 20208 1606 20214 1658
rect 20266 1606 20278 1658
rect 20330 1606 20342 1658
rect 20394 1606 20406 1658
rect 20458 1606 20470 1658
rect 20522 1606 20528 1658
rect 20076 1556 20128 1562
rect 20076 1498 20128 1504
rect 20076 1284 20128 1290
rect 20076 1226 20128 1232
rect 19984 1216 20036 1222
rect 19984 1158 20036 1164
rect 20088 1018 20116 1226
rect 20208 1040 20528 1606
rect 20076 1012 20128 1018
rect 20076 954 20128 960
rect 20364 870 20484 898
rect 19708 808 19760 814
rect 20364 800 20392 870
rect 19708 750 19760 756
rect 19340 740 19392 746
rect 19340 682 19392 688
rect 20350 0 20406 800
rect 20456 762 20484 870
rect 20640 762 20668 2382
rect 20732 2038 20760 3046
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20720 2032 20772 2038
rect 20720 1974 20772 1980
rect 20824 1766 20852 2926
rect 20916 2582 20944 4508
rect 21008 4282 21036 5170
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 21100 4146 21128 5510
rect 21192 5030 21220 6054
rect 21284 5778 21312 8774
rect 21376 8498 21404 9522
rect 21560 9518 21588 9930
rect 22112 9926 22140 9982
rect 21640 9920 21692 9926
rect 21640 9862 21692 9868
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 21548 9512 21600 9518
rect 21548 9454 21600 9460
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21364 8492 21416 8498
rect 21364 8434 21416 8440
rect 21364 8356 21416 8362
rect 21364 8298 21416 8304
rect 21376 6730 21404 8298
rect 21468 7206 21496 8910
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21456 7200 21508 7206
rect 21456 7142 21508 7148
rect 21364 6724 21416 6730
rect 21364 6666 21416 6672
rect 21272 5772 21324 5778
rect 21272 5714 21324 5720
rect 21364 5568 21416 5574
rect 21364 5510 21416 5516
rect 21376 5302 21404 5510
rect 21364 5296 21416 5302
rect 21364 5238 21416 5244
rect 21364 5160 21416 5166
rect 21364 5102 21416 5108
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21192 4162 21220 4966
rect 21088 4140 21140 4146
rect 21192 4134 21312 4162
rect 21088 4082 21140 4088
rect 21180 4072 21232 4078
rect 21180 4014 21232 4020
rect 21192 3602 21220 4014
rect 21180 3596 21232 3602
rect 21180 3538 21232 3544
rect 20996 3392 21048 3398
rect 20996 3334 21048 3340
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 21008 3194 21036 3334
rect 20996 3188 21048 3194
rect 20996 3130 21048 3136
rect 20904 2576 20956 2582
rect 20904 2518 20956 2524
rect 21100 2378 21128 3334
rect 21192 2854 21220 3538
rect 21284 2990 21312 4134
rect 21376 3738 21404 5102
rect 21364 3732 21416 3738
rect 21364 3674 21416 3680
rect 21364 3596 21416 3602
rect 21364 3538 21416 3544
rect 21376 3466 21404 3538
rect 21364 3460 21416 3466
rect 21364 3402 21416 3408
rect 21272 2984 21324 2990
rect 21272 2926 21324 2932
rect 21180 2848 21232 2854
rect 21180 2790 21232 2796
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 20812 1760 20864 1766
rect 20812 1702 20864 1708
rect 21100 1562 21128 2314
rect 21088 1556 21140 1562
rect 21088 1498 21140 1504
rect 21468 950 21496 7142
rect 21560 6390 21588 8570
rect 21652 8294 21680 9862
rect 22192 9716 22244 9722
rect 22192 9658 22244 9664
rect 22100 9648 22152 9654
rect 22100 9590 22152 9596
rect 21916 9104 21968 9110
rect 21916 9046 21968 9052
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 21732 8560 21784 8566
rect 21732 8502 21784 8508
rect 21640 8288 21692 8294
rect 21640 8230 21692 8236
rect 21744 7478 21772 8502
rect 21836 7750 21864 8910
rect 21928 8022 21956 9046
rect 21916 8016 21968 8022
rect 21916 7958 21968 7964
rect 22112 7954 22140 9590
rect 22204 8566 22232 9658
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 9058 22324 9318
rect 22388 9178 22416 14962
rect 22480 14958 22508 15150
rect 22468 14952 22520 14958
rect 22468 14894 22520 14900
rect 22560 14408 22612 14414
rect 22560 14350 22612 14356
rect 22572 14006 22600 14350
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 22468 13524 22520 13530
rect 22468 13466 22520 13472
rect 22480 12238 22508 13466
rect 22836 13320 22888 13326
rect 22836 13262 22888 13268
rect 22848 12850 22876 13262
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22744 11756 22796 11762
rect 22744 11698 22796 11704
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22468 10124 22520 10130
rect 22468 10066 22520 10072
rect 22480 9722 22508 10066
rect 22572 9722 22600 10542
rect 22652 10532 22704 10538
rect 22652 10474 22704 10480
rect 22664 10266 22692 10474
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22652 9988 22704 9994
rect 22652 9930 22704 9936
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22560 9716 22612 9722
rect 22560 9658 22612 9664
rect 22664 9178 22692 9930
rect 22376 9172 22428 9178
rect 22376 9114 22428 9120
rect 22652 9172 22704 9178
rect 22652 9114 22704 9120
rect 22296 9030 22416 9058
rect 22192 8560 22244 8566
rect 22192 8502 22244 8508
rect 22100 7948 22152 7954
rect 22100 7890 22152 7896
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21732 7472 21784 7478
rect 21732 7414 21784 7420
rect 21548 6384 21600 6390
rect 21548 6326 21600 6332
rect 21560 5370 21588 6326
rect 21640 6112 21692 6118
rect 21640 6054 21692 6060
rect 21548 5364 21600 5370
rect 21548 5306 21600 5312
rect 21560 4690 21588 5306
rect 21548 4684 21600 4690
rect 21548 4626 21600 4632
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21560 3670 21588 4218
rect 21548 3664 21600 3670
rect 21548 3606 21600 3612
rect 21652 3058 21680 6054
rect 21744 5234 21772 7414
rect 21732 5228 21784 5234
rect 21732 5170 21784 5176
rect 21732 4480 21784 4486
rect 21732 4422 21784 4428
rect 21744 4214 21772 4422
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 21744 3602 21772 4150
rect 21732 3596 21784 3602
rect 21732 3538 21784 3544
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 21836 1193 21864 7686
rect 22112 6866 22140 7754
rect 22204 7410 22232 8502
rect 22284 8424 22336 8430
rect 22284 8366 22336 8372
rect 22296 8090 22324 8366
rect 22284 8084 22336 8090
rect 22284 8026 22336 8032
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 22204 7018 22232 7346
rect 22388 7206 22416 9030
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22572 7478 22600 7686
rect 22560 7472 22612 7478
rect 22560 7414 22612 7420
rect 22664 7342 22692 7890
rect 22756 7750 22784 11698
rect 22848 11150 22876 12786
rect 22836 11144 22888 11150
rect 22836 11086 22888 11092
rect 22836 10464 22888 10470
rect 22836 10406 22888 10412
rect 22848 9654 22876 10406
rect 22940 10130 22968 17070
rect 23308 17066 23336 17614
rect 23400 17270 23428 18022
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23308 16726 23336 17002
rect 23296 16720 23348 16726
rect 23296 16662 23348 16668
rect 23308 16574 23336 16662
rect 23124 16546 23336 16574
rect 23124 16114 23152 16546
rect 23492 16182 23520 18226
rect 23572 16516 23624 16522
rect 23572 16458 23624 16464
rect 23480 16176 23532 16182
rect 23480 16118 23532 16124
rect 23112 16108 23164 16114
rect 23112 16050 23164 16056
rect 23204 16108 23256 16114
rect 23204 16050 23256 16056
rect 23020 14816 23072 14822
rect 23020 14758 23072 14764
rect 23032 13258 23060 14758
rect 23124 14550 23152 16050
rect 23216 15502 23244 16050
rect 23296 15904 23348 15910
rect 23296 15846 23348 15852
rect 23204 15496 23256 15502
rect 23204 15438 23256 15444
rect 23112 14544 23164 14550
rect 23112 14486 23164 14492
rect 23020 13252 23072 13258
rect 23020 13194 23072 13200
rect 23112 12776 23164 12782
rect 23112 12718 23164 12724
rect 23020 11756 23072 11762
rect 23020 11698 23072 11704
rect 23032 11218 23060 11698
rect 23124 11354 23152 12718
rect 23308 12434 23336 15846
rect 23388 15564 23440 15570
rect 23388 15506 23440 15512
rect 23400 15094 23428 15506
rect 23492 15502 23520 16118
rect 23584 15502 23612 16458
rect 23676 16250 23704 18294
rect 24124 18284 24176 18290
rect 24124 18226 24176 18232
rect 23756 18080 23808 18086
rect 23756 18022 23808 18028
rect 23664 16244 23716 16250
rect 23664 16186 23716 16192
rect 23480 15496 23532 15502
rect 23480 15438 23532 15444
rect 23572 15496 23624 15502
rect 23572 15438 23624 15444
rect 23584 15094 23612 15438
rect 23768 15178 23796 18022
rect 23940 17536 23992 17542
rect 23940 17478 23992 17484
rect 23952 17202 23980 17478
rect 24136 17338 24164 18226
rect 24208 17434 24528 18470
rect 24208 17382 24214 17434
rect 24266 17382 24278 17434
rect 24330 17382 24342 17434
rect 24394 17382 24406 17434
rect 24458 17382 24470 17434
rect 24522 17382 24528 17434
rect 24124 17332 24176 17338
rect 24124 17274 24176 17280
rect 23940 17196 23992 17202
rect 23940 17138 23992 17144
rect 24208 16518 24528 17382
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24208 16462 24220 16518
rect 24276 16462 24300 16518
rect 24356 16462 24380 16518
rect 24436 16462 24460 16518
rect 24516 16462 24528 16518
rect 24208 16438 24528 16462
rect 24208 16382 24220 16438
rect 24276 16382 24300 16438
rect 24356 16382 24380 16438
rect 24436 16382 24460 16438
rect 24516 16382 24528 16438
rect 24208 16358 24528 16382
rect 24208 16346 24220 16358
rect 24276 16346 24300 16358
rect 24356 16346 24380 16358
rect 24436 16346 24460 16358
rect 24516 16346 24528 16358
rect 24208 16294 24214 16346
rect 24276 16302 24278 16346
rect 24458 16302 24460 16346
rect 24266 16294 24278 16302
rect 24330 16294 24342 16302
rect 24394 16294 24406 16302
rect 24458 16294 24470 16302
rect 24522 16294 24528 16346
rect 24208 16278 24528 16294
rect 24208 16222 24220 16278
rect 24276 16222 24300 16278
rect 24356 16222 24380 16278
rect 24436 16222 24460 16278
rect 24516 16222 24528 16278
rect 23940 15360 23992 15366
rect 23940 15302 23992 15308
rect 23676 15150 23796 15178
rect 23388 15088 23440 15094
rect 23388 15030 23440 15036
rect 23572 15088 23624 15094
rect 23572 15030 23624 15036
rect 23676 14346 23704 15150
rect 23756 15020 23808 15026
rect 23756 14962 23808 14968
rect 23768 14550 23796 14962
rect 23756 14544 23808 14550
rect 23756 14486 23808 14492
rect 23664 14340 23716 14346
rect 23664 14282 23716 14288
rect 23756 14272 23808 14278
rect 23756 14214 23808 14220
rect 23768 14006 23796 14214
rect 23952 14006 23980 15302
rect 24208 15258 24528 16222
rect 24208 15206 24214 15258
rect 24266 15206 24278 15258
rect 24330 15206 24342 15258
rect 24394 15206 24406 15258
rect 24458 15206 24470 15258
rect 24522 15206 24528 15258
rect 24124 15020 24176 15026
rect 24124 14962 24176 14968
rect 23756 14000 23808 14006
rect 23756 13942 23808 13948
rect 23940 14000 23992 14006
rect 23940 13942 23992 13948
rect 24032 13864 24084 13870
rect 24032 13806 24084 13812
rect 23480 13320 23532 13326
rect 23480 13262 23532 13268
rect 23216 12406 23336 12434
rect 23112 11348 23164 11354
rect 23112 11290 23164 11296
rect 23020 11212 23072 11218
rect 23020 11154 23072 11160
rect 23112 11008 23164 11014
rect 23112 10950 23164 10956
rect 23124 10130 23152 10950
rect 22928 10124 22980 10130
rect 22928 10066 22980 10072
rect 23112 10124 23164 10130
rect 23112 10066 23164 10072
rect 22836 9648 22888 9654
rect 22836 9590 22888 9596
rect 23216 9178 23244 12406
rect 23388 11756 23440 11762
rect 23388 11698 23440 11704
rect 23400 11082 23428 11698
rect 23388 11076 23440 11082
rect 23388 11018 23440 11024
rect 23400 10810 23428 11018
rect 23388 10804 23440 10810
rect 23388 10746 23440 10752
rect 23296 10736 23348 10742
rect 23296 10678 23348 10684
rect 23308 10266 23336 10678
rect 23388 10668 23440 10674
rect 23388 10610 23440 10616
rect 23296 10260 23348 10266
rect 23296 10202 23348 10208
rect 23400 9518 23428 10610
rect 23492 10606 23520 13262
rect 23664 13252 23716 13258
rect 23664 13194 23716 13200
rect 23676 12374 23704 13194
rect 23664 12368 23716 12374
rect 23664 12310 23716 12316
rect 23676 11150 23704 12310
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23860 11830 23888 12174
rect 23848 11824 23900 11830
rect 23848 11766 23900 11772
rect 23664 11144 23716 11150
rect 23664 11086 23716 11092
rect 23572 11076 23624 11082
rect 23572 11018 23624 11024
rect 23584 10810 23612 11018
rect 23664 11008 23716 11014
rect 23664 10950 23716 10956
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23480 10600 23532 10606
rect 23480 10542 23532 10548
rect 23572 10056 23624 10062
rect 23572 9998 23624 10004
rect 23480 9648 23532 9654
rect 23480 9590 23532 9596
rect 23388 9512 23440 9518
rect 23388 9454 23440 9460
rect 23204 9172 23256 9178
rect 23204 9114 23256 9120
rect 23296 8356 23348 8362
rect 23296 8298 23348 8304
rect 23308 7886 23336 8298
rect 23400 7954 23428 9454
rect 23492 9178 23520 9590
rect 23480 9172 23532 9178
rect 23480 9114 23532 9120
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 23020 7812 23072 7818
rect 23020 7754 23072 7760
rect 22744 7744 22796 7750
rect 22744 7686 22796 7692
rect 22940 7342 22968 7754
rect 22652 7336 22704 7342
rect 22652 7278 22704 7284
rect 22928 7336 22980 7342
rect 22928 7278 22980 7284
rect 22376 7200 22428 7206
rect 22376 7142 22428 7148
rect 22204 6990 22416 7018
rect 22100 6860 22152 6866
rect 22100 6802 22152 6808
rect 22284 6860 22336 6866
rect 22284 6802 22336 6808
rect 22008 6656 22060 6662
rect 22008 6598 22060 6604
rect 22020 5846 22048 6598
rect 22296 6474 22324 6802
rect 22112 6458 22324 6474
rect 22100 6452 22324 6458
rect 22152 6446 22324 6452
rect 22100 6394 22152 6400
rect 22008 5840 22060 5846
rect 22008 5782 22060 5788
rect 21916 5772 21968 5778
rect 21916 5714 21968 5720
rect 21928 4010 21956 5714
rect 22112 4706 22140 6394
rect 22388 6254 22416 6990
rect 22664 6254 22692 7278
rect 23032 6866 23060 7754
rect 23296 7200 23348 7206
rect 23348 7148 23428 7154
rect 23296 7142 23428 7148
rect 23308 7126 23428 7142
rect 23020 6860 23072 6866
rect 23020 6802 23072 6808
rect 23032 6746 23060 6802
rect 23032 6718 23244 6746
rect 23020 6656 23072 6662
rect 23020 6598 23072 6604
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 22376 6248 22428 6254
rect 22376 6190 22428 6196
rect 22652 6248 22704 6254
rect 22652 6190 22704 6196
rect 22284 6112 22336 6118
rect 22284 6054 22336 6060
rect 22296 5710 22324 6054
rect 22388 5778 22416 6190
rect 23032 5778 23060 6598
rect 23124 6458 23152 6598
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 22376 5772 22428 5778
rect 22376 5714 22428 5720
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22020 4678 22140 4706
rect 22020 4078 22048 4678
rect 22100 4548 22152 4554
rect 22100 4490 22152 4496
rect 22008 4072 22060 4078
rect 22008 4014 22060 4020
rect 21916 4004 21968 4010
rect 21916 3946 21968 3952
rect 21916 3732 21968 3738
rect 21916 3674 21968 3680
rect 21928 1562 21956 3674
rect 22112 3534 22140 4490
rect 22100 3528 22152 3534
rect 22100 3470 22152 3476
rect 22192 3528 22244 3534
rect 22192 3470 22244 3476
rect 22100 3120 22152 3126
rect 22100 3062 22152 3068
rect 22112 1902 22140 3062
rect 22204 2446 22232 3470
rect 22296 3369 22324 5646
rect 22652 5636 22704 5642
rect 22652 5578 22704 5584
rect 22664 5370 22692 5578
rect 23032 5370 23060 5714
rect 22652 5364 22704 5370
rect 22652 5306 22704 5312
rect 23020 5364 23072 5370
rect 23020 5306 23072 5312
rect 23216 5250 23244 6718
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23308 6118 23336 6598
rect 23400 6186 23428 7126
rect 23388 6180 23440 6186
rect 23388 6122 23440 6128
rect 23296 6112 23348 6118
rect 23296 6054 23348 6060
rect 23308 5370 23336 6054
rect 23478 5536 23534 5545
rect 23478 5471 23534 5480
rect 23296 5364 23348 5370
rect 23296 5306 23348 5312
rect 23216 5222 23428 5250
rect 22744 5024 22796 5030
rect 22744 4966 22796 4972
rect 22376 4820 22428 4826
rect 22376 4762 22428 4768
rect 22388 4729 22416 4762
rect 22374 4720 22430 4729
rect 22374 4655 22430 4664
rect 22560 4072 22612 4078
rect 22560 4014 22612 4020
rect 22572 3738 22600 4014
rect 22560 3732 22612 3738
rect 22560 3674 22612 3680
rect 22376 3460 22428 3466
rect 22376 3402 22428 3408
rect 22282 3360 22338 3369
rect 22282 3295 22338 3304
rect 22388 3126 22416 3402
rect 22560 3188 22612 3194
rect 22560 3130 22612 3136
rect 22376 3120 22428 3126
rect 22376 3062 22428 3068
rect 22468 2644 22520 2650
rect 22468 2586 22520 2592
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 22100 1896 22152 1902
rect 22100 1838 22152 1844
rect 22008 1760 22060 1766
rect 22008 1702 22060 1708
rect 22020 1562 22048 1702
rect 21916 1556 21968 1562
rect 21916 1498 21968 1504
rect 22008 1556 22060 1562
rect 22008 1498 22060 1504
rect 22100 1352 22152 1358
rect 22100 1294 22152 1300
rect 21822 1184 21878 1193
rect 21822 1119 21878 1128
rect 22112 950 22140 1294
rect 21456 944 21508 950
rect 21456 886 21508 892
rect 22100 944 22152 950
rect 22100 886 22152 892
rect 22480 800 22508 2586
rect 22572 2514 22600 3130
rect 22560 2508 22612 2514
rect 22560 2450 22612 2456
rect 22756 1358 22784 4966
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23032 2446 23060 4762
rect 23216 4690 23244 5222
rect 23400 5166 23428 5222
rect 23388 5160 23440 5166
rect 23388 5102 23440 5108
rect 23204 4684 23256 4690
rect 23204 4626 23256 4632
rect 23216 4570 23244 4626
rect 23124 4542 23244 4570
rect 23124 3602 23152 4542
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23388 4480 23440 4486
rect 23388 4422 23440 4428
rect 23204 4072 23256 4078
rect 23308 4060 23336 4422
rect 23256 4032 23336 4060
rect 23204 4014 23256 4020
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 23124 2514 23152 3538
rect 23308 3534 23336 4032
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23400 3194 23428 4422
rect 23492 4282 23520 5471
rect 23480 4276 23532 4282
rect 23480 4218 23532 4224
rect 23584 4162 23612 9998
rect 23676 9178 23704 10950
rect 23860 10674 23888 11766
rect 23848 10668 23900 10674
rect 23848 10610 23900 10616
rect 24044 10266 24072 13806
rect 24136 13190 24164 14962
rect 24208 14170 24528 15206
rect 24596 14249 24624 17274
rect 25042 16416 25098 16425
rect 25042 16351 25098 16360
rect 24676 16108 24728 16114
rect 24676 16050 24728 16056
rect 24582 14240 24638 14249
rect 24582 14175 24638 14184
rect 24208 14118 24214 14170
rect 24266 14118 24278 14170
rect 24330 14118 24342 14170
rect 24394 14118 24406 14170
rect 24458 14118 24470 14170
rect 24522 14118 24528 14170
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24136 12073 24164 13126
rect 24208 13082 24528 14118
rect 24208 13030 24214 13082
rect 24266 13030 24278 13082
rect 24330 13030 24342 13082
rect 24394 13030 24406 13082
rect 24458 13030 24470 13082
rect 24522 13030 24528 13082
rect 24122 12064 24178 12073
rect 24122 11999 24178 12008
rect 24208 11994 24528 13030
rect 24208 11942 24214 11994
rect 24266 11942 24278 11994
rect 24330 11942 24342 11994
rect 24394 11942 24406 11994
rect 24458 11942 24470 11994
rect 24522 11942 24528 11994
rect 24208 10906 24528 11942
rect 24208 10854 24214 10906
rect 24266 10854 24278 10906
rect 24330 10854 24342 10906
rect 24394 10854 24406 10906
rect 24458 10854 24470 10906
rect 24522 10854 24528 10906
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 24122 9888 24178 9897
rect 24122 9823 24178 9832
rect 23756 9716 23808 9722
rect 23756 9658 23808 9664
rect 23664 9172 23716 9178
rect 23664 9114 23716 9120
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23676 7886 23704 8230
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23768 6866 23796 9658
rect 24136 8974 24164 9823
rect 24208 9818 24528 10854
rect 24208 9766 24214 9818
rect 24266 9766 24278 9818
rect 24330 9766 24342 9818
rect 24394 9766 24406 9818
rect 24458 9766 24470 9818
rect 24522 9766 24528 9818
rect 24124 8968 24176 8974
rect 24044 8928 24124 8956
rect 23848 8288 23900 8294
rect 23848 8230 23900 8236
rect 23860 8022 23888 8230
rect 23848 8016 23900 8022
rect 23848 7958 23900 7964
rect 24044 7562 24072 8928
rect 24124 8910 24176 8916
rect 24208 8730 24528 9766
rect 24688 8906 24716 16050
rect 25056 14890 25084 16351
rect 25044 14884 25096 14890
rect 25044 14826 25096 14832
rect 24676 8900 24728 8906
rect 24676 8842 24728 8848
rect 24208 8678 24214 8730
rect 24266 8678 24278 8730
rect 24330 8678 24342 8730
rect 24394 8678 24406 8730
rect 24458 8678 24470 8730
rect 24522 8678 24528 8730
rect 24208 8518 24528 8678
rect 24208 8462 24220 8518
rect 24276 8462 24300 8518
rect 24356 8462 24380 8518
rect 24436 8462 24460 8518
rect 24516 8462 24528 8518
rect 24676 8560 24728 8566
rect 24676 8502 24728 8508
rect 24208 8438 24528 8462
rect 24208 8382 24220 8438
rect 24276 8382 24300 8438
rect 24356 8382 24380 8438
rect 24436 8382 24460 8438
rect 24516 8382 24528 8438
rect 24208 8358 24528 8382
rect 24208 8302 24220 8358
rect 24276 8302 24300 8358
rect 24356 8302 24380 8358
rect 24436 8302 24460 8358
rect 24516 8302 24528 8358
rect 24208 8278 24528 8302
rect 24208 8222 24220 8278
rect 24276 8222 24300 8278
rect 24356 8222 24380 8278
rect 24436 8222 24460 8278
rect 24516 8222 24528 8278
rect 24124 7880 24176 7886
rect 24124 7822 24176 7828
rect 24136 7721 24164 7822
rect 24122 7712 24178 7721
rect 24122 7647 24178 7656
rect 24208 7642 24528 8222
rect 24208 7590 24214 7642
rect 24266 7590 24278 7642
rect 24330 7590 24342 7642
rect 24394 7590 24406 7642
rect 24458 7590 24470 7642
rect 24522 7590 24528 7642
rect 24044 7534 24164 7562
rect 24032 7472 24084 7478
rect 24032 7414 24084 7420
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23664 5636 23716 5642
rect 23664 5578 23716 5584
rect 23492 4134 23612 4162
rect 23492 3670 23520 4134
rect 23480 3664 23532 3670
rect 23480 3606 23532 3612
rect 23572 3528 23624 3534
rect 23572 3470 23624 3476
rect 23584 3398 23612 3470
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23112 2508 23164 2514
rect 23112 2450 23164 2456
rect 23020 2440 23072 2446
rect 23020 2382 23072 2388
rect 23676 2106 23704 5578
rect 23768 4826 23796 6802
rect 24044 6458 24072 7414
rect 24032 6452 24084 6458
rect 24032 6394 24084 6400
rect 23940 6384 23992 6390
rect 23940 6326 23992 6332
rect 23952 5370 23980 6326
rect 23940 5364 23992 5370
rect 23940 5306 23992 5312
rect 24136 4826 24164 7534
rect 24208 6554 24528 7590
rect 24584 7200 24636 7206
rect 24584 7142 24636 7148
rect 24208 6502 24214 6554
rect 24266 6502 24278 6554
rect 24330 6502 24342 6554
rect 24394 6502 24406 6554
rect 24458 6502 24470 6554
rect 24522 6502 24528 6554
rect 24208 5466 24528 6502
rect 24596 5545 24624 7142
rect 24688 6390 24716 8502
rect 24676 6384 24728 6390
rect 24676 6326 24728 6332
rect 24688 5574 24716 6326
rect 24676 5568 24728 5574
rect 24582 5536 24638 5545
rect 24676 5510 24728 5516
rect 24582 5471 24638 5480
rect 24208 5414 24214 5466
rect 24266 5414 24278 5466
rect 24330 5414 24342 5466
rect 24394 5414 24406 5466
rect 24458 5414 24470 5466
rect 24522 5414 24528 5466
rect 23756 4820 23808 4826
rect 23756 4762 23808 4768
rect 24124 4820 24176 4826
rect 24124 4762 24176 4768
rect 23940 4480 23992 4486
rect 23940 4422 23992 4428
rect 23848 4004 23900 4010
rect 23848 3946 23900 3952
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3126 23796 3878
rect 23756 3120 23808 3126
rect 23756 3062 23808 3068
rect 23664 2100 23716 2106
rect 23664 2042 23716 2048
rect 23768 1970 23796 3062
rect 23860 2038 23888 3946
rect 23952 2990 23980 4422
rect 24208 4378 24528 5414
rect 24208 4326 24214 4378
rect 24266 4326 24278 4378
rect 24330 4326 24342 4378
rect 24394 4326 24406 4378
rect 24458 4326 24470 4378
rect 24522 4326 24528 4378
rect 24124 4208 24176 4214
rect 24124 4150 24176 4156
rect 24032 3732 24084 3738
rect 24032 3674 24084 3680
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 24044 2854 24072 3674
rect 24136 3670 24164 4150
rect 24124 3664 24176 3670
rect 24124 3606 24176 3612
rect 24208 3290 24528 4326
rect 24584 4140 24636 4146
rect 24584 4082 24636 4088
rect 24596 3534 24624 4082
rect 24584 3528 24636 3534
rect 24584 3470 24636 3476
rect 24208 3238 24214 3290
rect 24266 3238 24278 3290
rect 24330 3238 24342 3290
rect 24394 3238 24406 3290
rect 24458 3238 24470 3290
rect 24522 3238 24528 3290
rect 24032 2848 24084 2854
rect 23952 2796 24032 2802
rect 23952 2790 24084 2796
rect 23952 2774 24072 2790
rect 23848 2032 23900 2038
rect 23848 1974 23900 1980
rect 23756 1964 23808 1970
rect 23756 1906 23808 1912
rect 23768 1426 23796 1906
rect 23952 1766 23980 2774
rect 24208 2202 24528 3238
rect 24208 2150 24214 2202
rect 24266 2150 24278 2202
rect 24330 2150 24342 2202
rect 24394 2150 24406 2202
rect 24458 2150 24470 2202
rect 24522 2150 24528 2202
rect 23940 1760 23992 1766
rect 23940 1702 23992 1708
rect 23756 1420 23808 1426
rect 23756 1362 23808 1368
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 24208 1114 24528 2150
rect 24208 1062 24214 1114
rect 24266 1062 24278 1114
rect 24330 1062 24342 1114
rect 24394 1062 24406 1114
rect 24458 1062 24470 1114
rect 24522 1062 24528 1114
rect 24208 1040 24528 1062
rect 24596 800 24624 3470
rect 24688 3466 24716 5510
rect 24676 3460 24728 3466
rect 24676 3402 24728 3408
rect 24688 2038 24716 3402
rect 24768 3392 24820 3398
rect 24768 3334 24820 3340
rect 24780 2106 24808 3334
rect 24768 2100 24820 2106
rect 24768 2042 24820 2048
rect 24676 2032 24728 2038
rect 24676 1974 24728 1980
rect 20456 734 20668 762
rect 22466 0 22522 800
rect 24582 0 24638 800
<< via2 >>
rect 2962 18536 3018 18592
rect 1490 16108 1546 16144
rect 1490 16088 1492 16108
rect 1492 16088 1544 16108
rect 1544 16088 1546 16108
rect 1398 14184 1454 14240
rect 1306 12008 1362 12064
rect 1306 9832 1362 9888
rect 1398 7656 1454 7712
rect 1398 5480 1454 5536
rect 1674 8084 1730 8120
rect 1674 8064 1676 8084
rect 1676 8064 1728 8084
rect 1728 8064 1730 8084
rect 1490 3304 1546 3360
rect 1858 4700 1860 4720
rect 1860 4700 1912 4720
rect 1912 4700 1914 4720
rect 1858 4664 1914 4700
rect 2962 4684 3018 4720
rect 2962 4664 2964 4684
rect 2964 4664 3016 4684
rect 3016 4664 3018 4684
rect 3698 3168 3754 3224
rect 4220 12486 4266 12518
rect 4266 12486 4276 12518
rect 4300 12486 4330 12518
rect 4330 12486 4342 12518
rect 4342 12486 4356 12518
rect 4380 12486 4394 12518
rect 4394 12486 4406 12518
rect 4406 12486 4436 12518
rect 4460 12486 4470 12518
rect 4470 12486 4516 12518
rect 4220 12462 4276 12486
rect 4300 12462 4356 12486
rect 4380 12462 4436 12486
rect 4460 12462 4516 12486
rect 4220 12382 4276 12438
rect 4300 12382 4356 12438
rect 4380 12382 4436 12438
rect 4460 12382 4516 12438
rect 4220 12302 4276 12358
rect 4300 12302 4356 12358
rect 4380 12302 4436 12358
rect 4460 12302 4516 12358
rect 4220 12222 4276 12278
rect 4300 12222 4356 12278
rect 4380 12222 4436 12278
rect 4460 12222 4516 12278
rect 8220 16462 8276 16518
rect 8300 16462 8356 16518
rect 8380 16462 8436 16518
rect 8460 16462 8516 16518
rect 8220 16382 8276 16438
rect 8300 16382 8356 16438
rect 8380 16382 8436 16438
rect 8460 16382 8516 16438
rect 8220 16346 8276 16358
rect 8300 16346 8356 16358
rect 8380 16346 8436 16358
rect 8460 16346 8516 16358
rect 8220 16302 8266 16346
rect 8266 16302 8276 16346
rect 8300 16302 8330 16346
rect 8330 16302 8342 16346
rect 8342 16302 8356 16346
rect 8380 16302 8394 16346
rect 8394 16302 8406 16346
rect 8406 16302 8436 16346
rect 8460 16302 8470 16346
rect 8470 16302 8516 16346
rect 8220 16222 8276 16278
rect 8300 16222 8356 16278
rect 8380 16222 8436 16278
rect 8460 16222 8516 16278
rect 4220 4462 4276 4518
rect 4300 4462 4356 4518
rect 4380 4462 4436 4518
rect 4460 4462 4516 4518
rect 4220 4382 4276 4438
rect 4300 4382 4356 4438
rect 4380 4382 4436 4438
rect 4460 4382 4516 4438
rect 4220 4302 4276 4358
rect 4300 4302 4356 4358
rect 4380 4302 4436 4358
rect 4460 4302 4516 4358
rect 4220 4222 4276 4278
rect 4300 4222 4356 4278
rect 4380 4222 4436 4278
rect 4460 4222 4516 4278
rect 3974 3052 4030 3088
rect 3974 3032 3976 3052
rect 3976 3032 4028 3052
rect 4028 3032 4030 3052
rect 4986 3304 5042 3360
rect 4894 3052 4950 3088
rect 4894 3032 4896 3052
rect 4896 3032 4948 3052
rect 4948 3032 4950 3052
rect 5446 3168 5502 3224
rect 4802 2624 4858 2680
rect 5170 1400 5226 1456
rect 5814 3188 5870 3224
rect 5814 3168 5816 3188
rect 5816 3168 5868 3188
rect 5868 3168 5870 3188
rect 5998 3032 6054 3088
rect 7102 7828 7104 7848
rect 7104 7828 7156 7848
rect 7156 7828 7158 7848
rect 7102 7792 7158 7828
rect 7746 8064 7802 8120
rect 7930 7792 7986 7848
rect 10598 14884 10654 14920
rect 10598 14864 10600 14884
rect 10600 14864 10652 14884
rect 10652 14864 10654 14884
rect 10598 14456 10654 14512
rect 8220 8462 8276 8518
rect 8300 8462 8356 8518
rect 8380 8462 8436 8518
rect 8460 8462 8516 8518
rect 8220 8382 8276 8438
rect 8300 8382 8356 8438
rect 8380 8382 8436 8438
rect 8460 8382 8516 8438
rect 8220 8302 8276 8358
rect 8300 8302 8356 8358
rect 8380 8302 8436 8358
rect 8460 8302 8516 8358
rect 8220 8222 8276 8278
rect 8300 8222 8356 8278
rect 8380 8222 8436 8278
rect 8460 8222 8516 8278
rect 6274 3304 6330 3360
rect 6366 1128 6422 1184
rect 6734 3304 6790 3360
rect 6918 3168 6974 3224
rect 7470 3712 7526 3768
rect 10782 14356 10784 14376
rect 10784 14356 10836 14376
rect 10836 14356 10838 14376
rect 10782 14320 10838 14356
rect 10966 13504 11022 13560
rect 11150 13368 11206 13424
rect 11702 14320 11758 14376
rect 11426 13368 11482 13424
rect 8114 2624 8170 2680
rect 7838 2508 7894 2544
rect 7838 2488 7840 2508
rect 7840 2488 7892 2508
rect 7892 2488 7894 2508
rect 8022 1400 8078 1456
rect 9034 3712 9090 3768
rect 9770 4664 9826 4720
rect 9678 4020 9680 4040
rect 9680 4020 9732 4040
rect 9732 4020 9734 4040
rect 9678 3984 9734 4020
rect 9954 4664 10010 4720
rect 8850 2508 8906 2544
rect 8850 2488 8852 2508
rect 8852 2488 8904 2508
rect 8904 2488 8906 2508
rect 9494 1400 9550 1456
rect 9862 2508 9918 2544
rect 9862 2488 9864 2508
rect 9864 2488 9916 2508
rect 9916 2488 9918 2508
rect 10046 2216 10102 2272
rect 12070 14492 12072 14512
rect 12072 14492 12124 14512
rect 12124 14492 12126 14512
rect 12070 14456 12126 14492
rect 11886 13776 11942 13832
rect 12220 12486 12266 12518
rect 12266 12486 12276 12518
rect 12300 12486 12330 12518
rect 12330 12486 12342 12518
rect 12342 12486 12356 12518
rect 12380 12486 12394 12518
rect 12394 12486 12406 12518
rect 12406 12486 12436 12518
rect 12460 12486 12470 12518
rect 12470 12486 12516 12518
rect 12220 12462 12276 12486
rect 12300 12462 12356 12486
rect 12380 12462 12436 12486
rect 12460 12462 12516 12486
rect 12220 12382 12276 12438
rect 12300 12382 12356 12438
rect 12380 12382 12436 12438
rect 12460 12382 12516 12438
rect 12220 12302 12276 12358
rect 12300 12302 12356 12358
rect 12380 12302 12436 12358
rect 12460 12302 12516 12358
rect 12220 12222 12276 12278
rect 12300 12222 12356 12278
rect 12380 12222 12436 12278
rect 12460 12222 12516 12278
rect 13634 13368 13690 13424
rect 10690 7812 10746 7848
rect 10690 7792 10692 7812
rect 10692 7792 10744 7812
rect 10744 7792 10746 7812
rect 10230 4800 10286 4856
rect 10598 6316 10654 6352
rect 10598 6296 10600 6316
rect 10600 6296 10652 6316
rect 10652 6296 10654 6316
rect 10230 3984 10286 4040
rect 10874 2624 10930 2680
rect 10414 2352 10470 2408
rect 10690 1556 10746 1592
rect 10874 2216 10930 2272
rect 11426 4664 11482 4720
rect 11426 2760 11482 2816
rect 11702 5888 11758 5944
rect 10690 1536 10692 1556
rect 10692 1536 10744 1556
rect 10744 1536 10746 1556
rect 10874 1420 10930 1456
rect 10874 1400 10876 1420
rect 10876 1400 10928 1420
rect 10928 1400 10930 1420
rect 12806 4800 12862 4856
rect 12220 4462 12276 4518
rect 12300 4462 12356 4518
rect 12380 4462 12436 4518
rect 12460 4462 12516 4518
rect 12220 4382 12276 4438
rect 12300 4382 12356 4438
rect 12380 4382 12436 4438
rect 12460 4382 12516 4438
rect 12220 4302 12276 4358
rect 12300 4302 12356 4358
rect 12380 4302 12436 4358
rect 12460 4302 12516 4358
rect 12220 4222 12276 4278
rect 12300 4222 12356 4278
rect 12380 4222 12436 4278
rect 12460 4222 12516 4278
rect 11978 3984 12034 4040
rect 11886 3032 11942 3088
rect 12622 2388 12624 2408
rect 12624 2388 12676 2408
rect 12676 2388 12678 2408
rect 12622 2352 12678 2388
rect 12070 1536 12126 1592
rect 12070 1436 12072 1456
rect 12072 1436 12124 1456
rect 12124 1436 12126 1456
rect 12070 1400 12126 1436
rect 11058 1300 11060 1320
rect 11060 1300 11112 1320
rect 11112 1300 11114 1320
rect 11058 1264 11114 1300
rect 12806 2488 12862 2544
rect 14002 13812 14004 13832
rect 14004 13812 14056 13832
rect 14056 13812 14058 13832
rect 14002 13776 14058 13812
rect 15290 16088 15346 16144
rect 14830 15544 14886 15600
rect 14646 15428 14702 15464
rect 14646 15408 14648 15428
rect 14648 15408 14700 15428
rect 14700 15408 14702 15428
rect 16220 16462 16276 16518
rect 16300 16462 16356 16518
rect 16380 16462 16436 16518
rect 16460 16462 16516 16518
rect 16220 16382 16276 16438
rect 16300 16382 16356 16438
rect 16380 16382 16436 16438
rect 16460 16382 16516 16438
rect 16220 16346 16276 16358
rect 16300 16346 16356 16358
rect 16380 16346 16436 16358
rect 16460 16346 16516 16358
rect 16220 16302 16266 16346
rect 16266 16302 16276 16346
rect 16300 16302 16330 16346
rect 16330 16302 16342 16346
rect 16342 16302 16356 16346
rect 16380 16302 16394 16346
rect 16394 16302 16406 16346
rect 16406 16302 16436 16346
rect 16460 16302 16470 16346
rect 16470 16302 16516 16346
rect 16220 16222 16276 16278
rect 16300 16222 16356 16278
rect 16380 16222 16436 16278
rect 16460 16222 16516 16278
rect 13174 7828 13176 7848
rect 13176 7828 13228 7848
rect 13228 7828 13230 7848
rect 13174 7792 13230 7828
rect 13358 4664 13414 4720
rect 15934 15544 15990 15600
rect 15842 14592 15898 14648
rect 15842 13504 15898 13560
rect 16762 16088 16818 16144
rect 16578 15544 16634 15600
rect 16946 14612 17002 14648
rect 16946 14592 16948 14612
rect 16948 14592 17000 14612
rect 17000 14592 17002 14612
rect 14462 9580 14518 9616
rect 14462 9560 14464 9580
rect 14464 9560 14516 9580
rect 14516 9560 14518 9580
rect 18142 15444 18144 15464
rect 18144 15444 18196 15464
rect 18196 15444 18198 15464
rect 18142 15408 18198 15444
rect 15750 9560 15806 9616
rect 18050 14884 18106 14920
rect 18050 14864 18052 14884
rect 18052 14864 18104 14884
rect 18104 14864 18106 14884
rect 17314 13368 17370 13424
rect 17498 13388 17554 13424
rect 17498 13368 17500 13388
rect 17500 13368 17552 13388
rect 17552 13368 17554 13388
rect 17958 13268 17960 13288
rect 17960 13268 18012 13288
rect 18012 13268 18014 13288
rect 17958 13232 18014 13268
rect 18418 13388 18474 13424
rect 18418 13368 18420 13388
rect 18420 13368 18472 13388
rect 18472 13368 18474 13388
rect 14462 7520 14518 7576
rect 14278 7420 14280 7440
rect 14280 7420 14332 7440
rect 14332 7420 14334 7440
rect 14278 7384 14334 7420
rect 14922 7420 14924 7440
rect 14924 7420 14976 7440
rect 14976 7420 14978 7440
rect 14922 7384 14978 7420
rect 16220 8462 16276 8518
rect 16300 8462 16356 8518
rect 16380 8462 16436 8518
rect 16460 8462 16516 8518
rect 16220 8382 16276 8438
rect 16300 8382 16356 8438
rect 16380 8382 16436 8438
rect 16460 8382 16516 8438
rect 15106 7520 15162 7576
rect 13450 3576 13506 3632
rect 13542 2216 13598 2272
rect 13174 1264 13230 1320
rect 14462 4684 14518 4720
rect 14462 4664 14464 4684
rect 14464 4664 14516 4684
rect 14516 4664 14518 4684
rect 14830 3032 14886 3088
rect 16220 8302 16276 8358
rect 16300 8302 16356 8358
rect 16380 8302 16436 8358
rect 16460 8302 16516 8358
rect 16220 8222 16276 8278
rect 16300 8222 16356 8278
rect 16380 8222 16436 8278
rect 16460 8222 16516 8278
rect 15290 3984 15346 4040
rect 17130 6568 17186 6624
rect 17038 6296 17094 6352
rect 16578 5752 16634 5808
rect 16670 5636 16726 5672
rect 16670 5616 16672 5636
rect 16672 5616 16724 5636
rect 16724 5616 16726 5636
rect 16026 3032 16082 3088
rect 15934 2508 15990 2544
rect 15934 2488 15936 2508
rect 15936 2488 15988 2508
rect 15988 2488 15990 2508
rect 16854 2352 16910 2408
rect 17406 5888 17462 5944
rect 17314 5772 17370 5808
rect 17314 5752 17316 5772
rect 17316 5752 17368 5772
rect 17368 5752 17370 5772
rect 17406 5636 17462 5672
rect 17406 5616 17408 5636
rect 17408 5616 17460 5636
rect 17460 5616 17462 5636
rect 17130 2896 17186 2952
rect 17406 2352 17462 2408
rect 19522 15000 19578 15056
rect 18878 13252 18934 13288
rect 18878 13232 18880 13252
rect 18880 13232 18932 13252
rect 18932 13232 18934 13252
rect 20626 15020 20682 15056
rect 20626 15000 20628 15020
rect 20628 15000 20680 15020
rect 20680 15000 20682 15020
rect 20902 15136 20958 15192
rect 20220 12486 20266 12518
rect 20266 12486 20276 12518
rect 20300 12486 20330 12518
rect 20330 12486 20342 12518
rect 20342 12486 20356 12518
rect 20380 12486 20394 12518
rect 20394 12486 20406 12518
rect 20406 12486 20436 12518
rect 20460 12486 20470 12518
rect 20470 12486 20516 12518
rect 20220 12462 20276 12486
rect 20300 12462 20356 12486
rect 20380 12462 20436 12486
rect 20460 12462 20516 12486
rect 20220 12382 20276 12438
rect 20300 12382 20356 12438
rect 20380 12382 20436 12438
rect 20460 12382 20516 12438
rect 19890 12008 19946 12064
rect 20220 12302 20276 12358
rect 20300 12302 20356 12358
rect 20380 12302 20436 12358
rect 20460 12302 20516 12358
rect 20220 12222 20276 12278
rect 20300 12222 20356 12278
rect 20380 12222 20436 12278
rect 20460 12222 20516 12278
rect 20074 11636 20082 11656
rect 20082 11636 20130 11656
rect 20074 11600 20130 11636
rect 20810 11600 20866 11656
rect 18418 6604 18420 6624
rect 18420 6604 18472 6624
rect 18472 6604 18474 6624
rect 18418 6568 18474 6604
rect 18234 5652 18236 5672
rect 18236 5652 18288 5672
rect 18288 5652 18290 5672
rect 18234 5616 18290 5652
rect 18050 3032 18106 3088
rect 18142 2624 18198 2680
rect 17958 2488 18014 2544
rect 18786 2760 18842 2816
rect 19062 2760 19118 2816
rect 21270 15020 21326 15056
rect 21270 15000 21272 15020
rect 21272 15000 21324 15020
rect 21324 15000 21326 15020
rect 21454 15136 21510 15192
rect 23478 18572 23480 18592
rect 23480 18572 23532 18592
rect 23532 18572 23534 18592
rect 23478 18536 23534 18572
rect 22282 15020 22338 15056
rect 22282 15000 22284 15020
rect 22284 15000 22336 15020
rect 22336 15000 22338 15020
rect 21914 12008 21970 12064
rect 19614 4684 19670 4720
rect 19614 4664 19616 4684
rect 19616 4664 19668 4684
rect 19668 4664 19670 4684
rect 19338 2896 19394 2952
rect 20220 4462 20276 4518
rect 20300 4462 20356 4518
rect 20380 4462 20436 4518
rect 20460 4462 20516 4518
rect 20220 4382 20276 4438
rect 20300 4382 20356 4438
rect 20380 4382 20436 4438
rect 20460 4382 20516 4438
rect 20220 4302 20276 4358
rect 20300 4302 20356 4358
rect 20380 4302 20436 4358
rect 20460 4302 20516 4358
rect 20220 4222 20276 4278
rect 20300 4222 20356 4278
rect 20380 4222 20436 4278
rect 20460 4222 20516 4278
rect 24220 16462 24276 16518
rect 24300 16462 24356 16518
rect 24380 16462 24436 16518
rect 24460 16462 24516 16518
rect 24220 16382 24276 16438
rect 24300 16382 24356 16438
rect 24380 16382 24436 16438
rect 24460 16382 24516 16438
rect 24220 16346 24276 16358
rect 24300 16346 24356 16358
rect 24380 16346 24436 16358
rect 24460 16346 24516 16358
rect 24220 16302 24266 16346
rect 24266 16302 24276 16346
rect 24300 16302 24330 16346
rect 24330 16302 24342 16346
rect 24342 16302 24356 16346
rect 24380 16302 24394 16346
rect 24394 16302 24406 16346
rect 24406 16302 24436 16346
rect 24460 16302 24470 16346
rect 24470 16302 24516 16346
rect 24220 16222 24276 16278
rect 24300 16222 24356 16278
rect 24380 16222 24436 16278
rect 24460 16222 24516 16278
rect 23478 5480 23534 5536
rect 22374 4664 22430 4720
rect 22282 3304 22338 3360
rect 21822 1128 21878 1184
rect 25042 16360 25098 16416
rect 24582 14184 24638 14240
rect 24122 12008 24178 12064
rect 24122 9832 24178 9888
rect 24220 8462 24276 8518
rect 24300 8462 24356 8518
rect 24380 8462 24436 8518
rect 24460 8462 24516 8518
rect 24220 8382 24276 8438
rect 24300 8382 24356 8438
rect 24380 8382 24436 8438
rect 24460 8382 24516 8438
rect 24220 8302 24276 8358
rect 24300 8302 24356 8358
rect 24380 8302 24436 8358
rect 24460 8302 24516 8358
rect 24220 8222 24276 8278
rect 24300 8222 24356 8278
rect 24380 8222 24436 8278
rect 24460 8222 24516 8278
rect 24122 7656 24178 7712
rect 24582 5480 24638 5536
<< metal3 >>
rect 0 18594 800 18624
rect 2957 18594 3023 18597
rect 0 18592 3023 18594
rect 0 18536 2962 18592
rect 3018 18536 3023 18592
rect 0 18534 3023 18536
rect 0 18504 800 18534
rect 2957 18531 3023 18534
rect 23473 18594 23539 18597
rect 25200 18594 26000 18624
rect 23473 18592 26000 18594
rect 23473 18536 23478 18592
rect 23534 18536 26000 18592
rect 23473 18534 26000 18536
rect 23473 18531 23539 18534
rect 25200 18504 26000 18534
rect 1056 16518 24888 16530
rect 1056 16462 8220 16518
rect 8276 16462 8300 16518
rect 8356 16462 8380 16518
rect 8436 16462 8460 16518
rect 8516 16462 16220 16518
rect 16276 16462 16300 16518
rect 16356 16462 16380 16518
rect 16436 16462 16460 16518
rect 16516 16462 24220 16518
rect 24276 16462 24300 16518
rect 24356 16462 24380 16518
rect 24436 16462 24460 16518
rect 24516 16462 24888 16518
rect 0 16418 800 16448
rect 1056 16438 24888 16462
rect 0 16328 858 16418
rect 798 16146 858 16328
rect 1056 16382 8220 16438
rect 8276 16382 8300 16438
rect 8356 16382 8380 16438
rect 8436 16382 8460 16438
rect 8516 16382 16220 16438
rect 16276 16382 16300 16438
rect 16356 16382 16380 16438
rect 16436 16382 16460 16438
rect 16516 16382 24220 16438
rect 24276 16382 24300 16438
rect 24356 16382 24380 16438
rect 24436 16382 24460 16438
rect 24516 16382 24888 16438
rect 1056 16358 24888 16382
rect 1056 16302 8220 16358
rect 8276 16302 8300 16358
rect 8356 16302 8380 16358
rect 8436 16302 8460 16358
rect 8516 16302 16220 16358
rect 16276 16302 16300 16358
rect 16356 16302 16380 16358
rect 16436 16302 16460 16358
rect 16516 16302 24220 16358
rect 24276 16302 24300 16358
rect 24356 16302 24380 16358
rect 24436 16302 24460 16358
rect 24516 16302 24888 16358
rect 25037 16418 25103 16421
rect 25200 16418 26000 16448
rect 25037 16416 26000 16418
rect 25037 16360 25042 16416
rect 25098 16360 26000 16416
rect 25037 16358 26000 16360
rect 25037 16355 25103 16358
rect 25200 16328 26000 16358
rect 1056 16278 24888 16302
rect 1056 16222 8220 16278
rect 8276 16222 8300 16278
rect 8356 16222 8380 16278
rect 8436 16222 8460 16278
rect 8516 16222 16220 16278
rect 16276 16222 16300 16278
rect 16356 16222 16380 16278
rect 16436 16222 16460 16278
rect 16516 16222 24220 16278
rect 24276 16222 24300 16278
rect 24356 16222 24380 16278
rect 24436 16222 24460 16278
rect 24516 16222 24888 16278
rect 1056 16210 24888 16222
rect 1485 16146 1551 16149
rect 798 16144 1551 16146
rect 798 16088 1490 16144
rect 1546 16088 1551 16144
rect 798 16086 1551 16088
rect 1485 16083 1551 16086
rect 15285 16146 15351 16149
rect 16757 16146 16823 16149
rect 15285 16144 16823 16146
rect 15285 16088 15290 16144
rect 15346 16088 16762 16144
rect 16818 16088 16823 16144
rect 15285 16086 16823 16088
rect 15285 16083 15351 16086
rect 16757 16083 16823 16086
rect 14825 15602 14891 15605
rect 15929 15602 15995 15605
rect 16573 15602 16639 15605
rect 14825 15600 16639 15602
rect 14825 15544 14830 15600
rect 14886 15544 15934 15600
rect 15990 15544 16578 15600
rect 16634 15544 16639 15600
rect 14825 15542 16639 15544
rect 14825 15539 14891 15542
rect 15929 15539 15995 15542
rect 16573 15539 16639 15542
rect 14641 15466 14707 15469
rect 18137 15466 18203 15469
rect 14641 15464 18203 15466
rect 14641 15408 14646 15464
rect 14702 15408 18142 15464
rect 18198 15408 18203 15464
rect 14641 15406 18203 15408
rect 14641 15403 14707 15406
rect 18137 15403 18203 15406
rect 20897 15194 20963 15197
rect 21449 15194 21515 15197
rect 20897 15192 21515 15194
rect 20897 15136 20902 15192
rect 20958 15136 21454 15192
rect 21510 15136 21515 15192
rect 20897 15134 21515 15136
rect 20897 15131 20963 15134
rect 21449 15131 21515 15134
rect 19517 15058 19583 15061
rect 20621 15058 20687 15061
rect 19517 15056 20687 15058
rect 19517 15000 19522 15056
rect 19578 15000 20626 15056
rect 20682 15000 20687 15056
rect 19517 14998 20687 15000
rect 19517 14995 19583 14998
rect 20621 14995 20687 14998
rect 21265 15058 21331 15061
rect 22277 15058 22343 15061
rect 21265 15056 22343 15058
rect 21265 15000 21270 15056
rect 21326 15000 22282 15056
rect 22338 15000 22343 15056
rect 21265 14998 22343 15000
rect 21265 14995 21331 14998
rect 22277 14995 22343 14998
rect 10593 14922 10659 14925
rect 18045 14922 18111 14925
rect 10593 14920 18111 14922
rect 10593 14864 10598 14920
rect 10654 14864 18050 14920
rect 18106 14864 18111 14920
rect 10593 14862 18111 14864
rect 10593 14859 10659 14862
rect 18045 14859 18111 14862
rect 15837 14650 15903 14653
rect 16941 14650 17007 14653
rect 15837 14648 17007 14650
rect 15837 14592 15842 14648
rect 15898 14592 16946 14648
rect 17002 14592 17007 14648
rect 15837 14590 17007 14592
rect 15837 14587 15903 14590
rect 16941 14587 17007 14590
rect 10593 14514 10659 14517
rect 12065 14514 12131 14517
rect 10593 14512 12131 14514
rect 10593 14456 10598 14512
rect 10654 14456 12070 14512
rect 12126 14456 12131 14512
rect 10593 14454 12131 14456
rect 10593 14451 10659 14454
rect 12065 14451 12131 14454
rect 10777 14378 10843 14381
rect 11697 14378 11763 14381
rect 10777 14376 11763 14378
rect 10777 14320 10782 14376
rect 10838 14320 11702 14376
rect 11758 14320 11763 14376
rect 10777 14318 11763 14320
rect 10777 14315 10843 14318
rect 11697 14315 11763 14318
rect 0 14242 800 14272
rect 1393 14242 1459 14245
rect 0 14240 1459 14242
rect 0 14184 1398 14240
rect 1454 14184 1459 14240
rect 0 14182 1459 14184
rect 0 14152 800 14182
rect 1393 14179 1459 14182
rect 24577 14242 24643 14245
rect 25200 14242 26000 14272
rect 24577 14240 26000 14242
rect 24577 14184 24582 14240
rect 24638 14184 26000 14240
rect 24577 14182 26000 14184
rect 24577 14179 24643 14182
rect 25200 14152 26000 14182
rect 11881 13834 11947 13837
rect 13997 13834 14063 13837
rect 11881 13832 14063 13834
rect 11881 13776 11886 13832
rect 11942 13776 14002 13832
rect 14058 13776 14063 13832
rect 11881 13774 14063 13776
rect 11881 13771 11947 13774
rect 13997 13771 14063 13774
rect 10961 13562 11027 13565
rect 15837 13562 15903 13565
rect 10961 13560 15903 13562
rect 10961 13504 10966 13560
rect 11022 13504 15842 13560
rect 15898 13504 15903 13560
rect 10961 13502 15903 13504
rect 10961 13499 11027 13502
rect 15837 13499 15903 13502
rect 11145 13426 11211 13429
rect 11421 13426 11487 13429
rect 13629 13426 13695 13429
rect 17309 13426 17375 13429
rect 11145 13424 17375 13426
rect 11145 13368 11150 13424
rect 11206 13368 11426 13424
rect 11482 13368 13634 13424
rect 13690 13368 17314 13424
rect 17370 13368 17375 13424
rect 11145 13366 17375 13368
rect 11145 13363 11211 13366
rect 11421 13363 11487 13366
rect 13629 13363 13695 13366
rect 17309 13363 17375 13366
rect 17493 13426 17559 13429
rect 18413 13426 18479 13429
rect 17493 13424 18479 13426
rect 17493 13368 17498 13424
rect 17554 13368 18418 13424
rect 18474 13368 18479 13424
rect 17493 13366 18479 13368
rect 17493 13363 17559 13366
rect 18413 13363 18479 13366
rect 17953 13290 18019 13293
rect 18873 13290 18939 13293
rect 17953 13288 18939 13290
rect 17953 13232 17958 13288
rect 18014 13232 18878 13288
rect 18934 13232 18939 13288
rect 17953 13230 18939 13232
rect 17953 13227 18019 13230
rect 18873 13227 18939 13230
rect 1056 12518 24888 12530
rect 1056 12462 4220 12518
rect 4276 12462 4300 12518
rect 4356 12462 4380 12518
rect 4436 12462 4460 12518
rect 4516 12462 12220 12518
rect 12276 12462 12300 12518
rect 12356 12462 12380 12518
rect 12436 12462 12460 12518
rect 12516 12462 20220 12518
rect 20276 12462 20300 12518
rect 20356 12462 20380 12518
rect 20436 12462 20460 12518
rect 20516 12462 24888 12518
rect 1056 12438 24888 12462
rect 1056 12382 4220 12438
rect 4276 12382 4300 12438
rect 4356 12382 4380 12438
rect 4436 12382 4460 12438
rect 4516 12382 12220 12438
rect 12276 12382 12300 12438
rect 12356 12382 12380 12438
rect 12436 12382 12460 12438
rect 12516 12382 20220 12438
rect 20276 12382 20300 12438
rect 20356 12382 20380 12438
rect 20436 12382 20460 12438
rect 20516 12382 24888 12438
rect 1056 12358 24888 12382
rect 1056 12302 4220 12358
rect 4276 12302 4300 12358
rect 4356 12302 4380 12358
rect 4436 12302 4460 12358
rect 4516 12302 12220 12358
rect 12276 12302 12300 12358
rect 12356 12302 12380 12358
rect 12436 12302 12460 12358
rect 12516 12302 20220 12358
rect 20276 12302 20300 12358
rect 20356 12302 20380 12358
rect 20436 12302 20460 12358
rect 20516 12302 24888 12358
rect 1056 12278 24888 12302
rect 1056 12222 4220 12278
rect 4276 12222 4300 12278
rect 4356 12222 4380 12278
rect 4436 12222 4460 12278
rect 4516 12222 12220 12278
rect 12276 12222 12300 12278
rect 12356 12222 12380 12278
rect 12436 12222 12460 12278
rect 12516 12222 20220 12278
rect 20276 12222 20300 12278
rect 20356 12222 20380 12278
rect 20436 12222 20460 12278
rect 20516 12222 24888 12278
rect 1056 12210 24888 12222
rect 0 12066 800 12096
rect 1301 12066 1367 12069
rect 0 12064 1367 12066
rect 0 12008 1306 12064
rect 1362 12008 1367 12064
rect 0 12006 1367 12008
rect 0 11976 800 12006
rect 1301 12003 1367 12006
rect 19885 12066 19951 12069
rect 21909 12066 21975 12069
rect 19885 12064 21975 12066
rect 19885 12008 19890 12064
rect 19946 12008 21914 12064
rect 21970 12008 21975 12064
rect 19885 12006 21975 12008
rect 19885 12003 19951 12006
rect 21909 12003 21975 12006
rect 24117 12066 24183 12069
rect 25200 12066 26000 12096
rect 24117 12064 26000 12066
rect 24117 12008 24122 12064
rect 24178 12008 26000 12064
rect 24117 12006 26000 12008
rect 24117 12003 24183 12006
rect 25200 11976 26000 12006
rect 20069 11658 20135 11661
rect 20805 11658 20871 11661
rect 20069 11656 20871 11658
rect 20069 11600 20074 11656
rect 20130 11600 20810 11656
rect 20866 11600 20871 11656
rect 20069 11598 20871 11600
rect 20069 11595 20135 11598
rect 20805 11595 20871 11598
rect 0 9890 800 9920
rect 1301 9890 1367 9893
rect 0 9888 1367 9890
rect 0 9832 1306 9888
rect 1362 9832 1367 9888
rect 0 9830 1367 9832
rect 0 9800 800 9830
rect 1301 9827 1367 9830
rect 24117 9890 24183 9893
rect 25200 9890 26000 9920
rect 24117 9888 26000 9890
rect 24117 9832 24122 9888
rect 24178 9832 26000 9888
rect 24117 9830 26000 9832
rect 24117 9827 24183 9830
rect 25200 9800 26000 9830
rect 14457 9618 14523 9621
rect 15745 9618 15811 9621
rect 14457 9616 15811 9618
rect 14457 9560 14462 9616
rect 14518 9560 15750 9616
rect 15806 9560 15811 9616
rect 14457 9558 15811 9560
rect 14457 9555 14523 9558
rect 15745 9555 15811 9558
rect 1056 8518 24888 8530
rect 1056 8462 8220 8518
rect 8276 8462 8300 8518
rect 8356 8462 8380 8518
rect 8436 8462 8460 8518
rect 8516 8462 16220 8518
rect 16276 8462 16300 8518
rect 16356 8462 16380 8518
rect 16436 8462 16460 8518
rect 16516 8462 24220 8518
rect 24276 8462 24300 8518
rect 24356 8462 24380 8518
rect 24436 8462 24460 8518
rect 24516 8462 24888 8518
rect 1056 8438 24888 8462
rect 1056 8382 8220 8438
rect 8276 8382 8300 8438
rect 8356 8382 8380 8438
rect 8436 8382 8460 8438
rect 8516 8382 16220 8438
rect 16276 8382 16300 8438
rect 16356 8382 16380 8438
rect 16436 8382 16460 8438
rect 16516 8382 24220 8438
rect 24276 8382 24300 8438
rect 24356 8382 24380 8438
rect 24436 8382 24460 8438
rect 24516 8382 24888 8438
rect 1056 8358 24888 8382
rect 1056 8302 8220 8358
rect 8276 8302 8300 8358
rect 8356 8302 8380 8358
rect 8436 8302 8460 8358
rect 8516 8302 16220 8358
rect 16276 8302 16300 8358
rect 16356 8302 16380 8358
rect 16436 8302 16460 8358
rect 16516 8302 24220 8358
rect 24276 8302 24300 8358
rect 24356 8302 24380 8358
rect 24436 8302 24460 8358
rect 24516 8302 24888 8358
rect 1056 8278 24888 8302
rect 1056 8222 8220 8278
rect 8276 8222 8300 8278
rect 8356 8222 8380 8278
rect 8436 8222 8460 8278
rect 8516 8222 16220 8278
rect 16276 8222 16300 8278
rect 16356 8222 16380 8278
rect 16436 8222 16460 8278
rect 16516 8222 24220 8278
rect 24276 8222 24300 8278
rect 24356 8222 24380 8278
rect 24436 8222 24460 8278
rect 24516 8222 24888 8278
rect 1056 8210 24888 8222
rect 1669 8122 1735 8125
rect 7741 8122 7807 8125
rect 1669 8120 7807 8122
rect 1669 8064 1674 8120
rect 1730 8064 7746 8120
rect 7802 8064 7807 8120
rect 1669 8062 7807 8064
rect 1669 8059 1735 8062
rect 7741 8059 7807 8062
rect 7097 7850 7163 7853
rect 7925 7850 7991 7853
rect 7097 7848 7991 7850
rect 7097 7792 7102 7848
rect 7158 7792 7930 7848
rect 7986 7792 7991 7848
rect 7097 7790 7991 7792
rect 7097 7787 7163 7790
rect 7925 7787 7991 7790
rect 10685 7850 10751 7853
rect 13169 7850 13235 7853
rect 10685 7848 13235 7850
rect 10685 7792 10690 7848
rect 10746 7792 13174 7848
rect 13230 7792 13235 7848
rect 10685 7790 13235 7792
rect 10685 7787 10751 7790
rect 13169 7787 13235 7790
rect 0 7714 800 7744
rect 1393 7714 1459 7717
rect 0 7712 1459 7714
rect 0 7656 1398 7712
rect 1454 7656 1459 7712
rect 0 7654 1459 7656
rect 0 7624 800 7654
rect 1393 7651 1459 7654
rect 24117 7714 24183 7717
rect 25200 7714 26000 7744
rect 24117 7712 26000 7714
rect 24117 7656 24122 7712
rect 24178 7656 26000 7712
rect 24117 7654 26000 7656
rect 24117 7651 24183 7654
rect 25200 7624 26000 7654
rect 14457 7578 14523 7581
rect 15101 7578 15167 7581
rect 14457 7576 15167 7578
rect 14457 7520 14462 7576
rect 14518 7520 15106 7576
rect 15162 7520 15167 7576
rect 14457 7518 15167 7520
rect 14457 7515 14523 7518
rect 15101 7515 15167 7518
rect 14273 7442 14339 7445
rect 14917 7442 14983 7445
rect 14273 7440 14983 7442
rect 14273 7384 14278 7440
rect 14334 7384 14922 7440
rect 14978 7384 14983 7440
rect 14273 7382 14983 7384
rect 14273 7379 14339 7382
rect 14917 7379 14983 7382
rect 17125 6626 17191 6629
rect 18413 6626 18479 6629
rect 17125 6624 18479 6626
rect 17125 6568 17130 6624
rect 17186 6568 18418 6624
rect 18474 6568 18479 6624
rect 17125 6566 18479 6568
rect 17125 6563 17191 6566
rect 18413 6563 18479 6566
rect 10593 6354 10659 6357
rect 17033 6354 17099 6357
rect 10593 6352 17099 6354
rect 10593 6296 10598 6352
rect 10654 6296 17038 6352
rect 17094 6296 17099 6352
rect 10593 6294 17099 6296
rect 10593 6291 10659 6294
rect 17033 6291 17099 6294
rect 11697 5946 11763 5949
rect 17401 5946 17467 5949
rect 11697 5944 17467 5946
rect 11697 5888 11702 5944
rect 11758 5888 17406 5944
rect 17462 5888 17467 5944
rect 11697 5886 17467 5888
rect 11697 5883 11763 5886
rect 17401 5883 17467 5886
rect 16573 5810 16639 5813
rect 17309 5810 17375 5813
rect 16573 5808 17375 5810
rect 16573 5752 16578 5808
rect 16634 5752 17314 5808
rect 17370 5752 17375 5808
rect 16573 5750 17375 5752
rect 16573 5747 16639 5750
rect 17309 5747 17375 5750
rect 16665 5674 16731 5677
rect 17401 5674 17467 5677
rect 18229 5674 18295 5677
rect 16665 5672 18295 5674
rect 16665 5616 16670 5672
rect 16726 5616 17406 5672
rect 17462 5616 18234 5672
rect 18290 5616 18295 5672
rect 16665 5614 18295 5616
rect 16665 5611 16731 5614
rect 17401 5611 17467 5614
rect 18229 5611 18295 5614
rect 0 5538 800 5568
rect 1393 5538 1459 5541
rect 0 5536 1459 5538
rect 0 5480 1398 5536
rect 1454 5480 1459 5536
rect 0 5478 1459 5480
rect 0 5448 800 5478
rect 1393 5475 1459 5478
rect 23473 5538 23539 5541
rect 24577 5538 24643 5541
rect 25200 5538 26000 5568
rect 23473 5536 26000 5538
rect 23473 5480 23478 5536
rect 23534 5480 24582 5536
rect 24638 5480 26000 5536
rect 23473 5478 26000 5480
rect 23473 5475 23539 5478
rect 24577 5475 24643 5478
rect 25200 5448 26000 5478
rect 10225 4858 10291 4861
rect 12801 4858 12867 4861
rect 10225 4856 12867 4858
rect 10225 4800 10230 4856
rect 10286 4800 12806 4856
rect 12862 4800 12867 4856
rect 10225 4798 12867 4800
rect 10225 4795 10291 4798
rect 12801 4795 12867 4798
rect 1853 4722 1919 4725
rect 2957 4722 3023 4725
rect 1853 4720 3023 4722
rect 1853 4664 1858 4720
rect 1914 4664 2962 4720
rect 3018 4664 3023 4720
rect 1853 4662 3023 4664
rect 1853 4659 1919 4662
rect 2957 4659 3023 4662
rect 9765 4722 9831 4725
rect 9949 4722 10015 4725
rect 11421 4722 11487 4725
rect 13353 4722 13419 4725
rect 14457 4722 14523 4725
rect 9765 4720 14523 4722
rect 9765 4664 9770 4720
rect 9826 4664 9954 4720
rect 10010 4664 11426 4720
rect 11482 4664 13358 4720
rect 13414 4664 14462 4720
rect 14518 4664 14523 4720
rect 9765 4662 14523 4664
rect 9765 4659 9831 4662
rect 9949 4659 10015 4662
rect 11421 4659 11487 4662
rect 13353 4659 13419 4662
rect 14457 4659 14523 4662
rect 19609 4722 19675 4725
rect 22369 4722 22435 4725
rect 19609 4720 22435 4722
rect 19609 4664 19614 4720
rect 19670 4664 22374 4720
rect 22430 4664 22435 4720
rect 19609 4662 22435 4664
rect 19609 4659 19675 4662
rect 22369 4659 22435 4662
rect 1056 4518 24888 4530
rect 1056 4462 4220 4518
rect 4276 4462 4300 4518
rect 4356 4462 4380 4518
rect 4436 4462 4460 4518
rect 4516 4462 12220 4518
rect 12276 4462 12300 4518
rect 12356 4462 12380 4518
rect 12436 4462 12460 4518
rect 12516 4462 20220 4518
rect 20276 4462 20300 4518
rect 20356 4462 20380 4518
rect 20436 4462 20460 4518
rect 20516 4462 24888 4518
rect 1056 4438 24888 4462
rect 1056 4382 4220 4438
rect 4276 4382 4300 4438
rect 4356 4382 4380 4438
rect 4436 4382 4460 4438
rect 4516 4382 12220 4438
rect 12276 4382 12300 4438
rect 12356 4382 12380 4438
rect 12436 4382 12460 4438
rect 12516 4382 20220 4438
rect 20276 4382 20300 4438
rect 20356 4382 20380 4438
rect 20436 4382 20460 4438
rect 20516 4382 24888 4438
rect 1056 4358 24888 4382
rect 1056 4302 4220 4358
rect 4276 4302 4300 4358
rect 4356 4302 4380 4358
rect 4436 4302 4460 4358
rect 4516 4302 12220 4358
rect 12276 4302 12300 4358
rect 12356 4302 12380 4358
rect 12436 4302 12460 4358
rect 12516 4302 20220 4358
rect 20276 4302 20300 4358
rect 20356 4302 20380 4358
rect 20436 4302 20460 4358
rect 20516 4302 24888 4358
rect 1056 4278 24888 4302
rect 1056 4222 4220 4278
rect 4276 4222 4300 4278
rect 4356 4222 4380 4278
rect 4436 4222 4460 4278
rect 4516 4222 12220 4278
rect 12276 4222 12300 4278
rect 12356 4222 12380 4278
rect 12436 4222 12460 4278
rect 12516 4222 20220 4278
rect 20276 4222 20300 4278
rect 20356 4222 20380 4278
rect 20436 4222 20460 4278
rect 20516 4222 24888 4278
rect 1056 4210 24888 4222
rect 9673 4042 9739 4045
rect 10225 4042 10291 4045
rect 9673 4040 10291 4042
rect 9673 3984 9678 4040
rect 9734 3984 10230 4040
rect 10286 3984 10291 4040
rect 9673 3982 10291 3984
rect 9673 3979 9739 3982
rect 10225 3979 10291 3982
rect 11973 4042 12039 4045
rect 15285 4042 15351 4045
rect 11973 4040 15351 4042
rect 11973 3984 11978 4040
rect 12034 3984 15290 4040
rect 15346 3984 15351 4040
rect 11973 3982 15351 3984
rect 11973 3979 12039 3982
rect 15285 3979 15351 3982
rect 7465 3770 7531 3773
rect 9029 3770 9095 3773
rect 7465 3768 9095 3770
rect 7465 3712 7470 3768
rect 7526 3712 9034 3768
rect 9090 3712 9095 3768
rect 7465 3710 9095 3712
rect 7465 3707 7531 3710
rect 9029 3707 9095 3710
rect 13445 3634 13511 3637
rect 13445 3632 15210 3634
rect 13445 3576 13450 3632
rect 13506 3576 15210 3632
rect 13445 3574 15210 3576
rect 13445 3571 13511 3574
rect 0 3362 800 3392
rect 1485 3362 1551 3365
rect 4981 3362 5047 3365
rect 0 3360 5047 3362
rect 0 3304 1490 3360
rect 1546 3304 4986 3360
rect 5042 3304 5047 3360
rect 0 3302 5047 3304
rect 0 3272 800 3302
rect 1485 3299 1551 3302
rect 4981 3299 5047 3302
rect 6269 3362 6335 3365
rect 6729 3362 6795 3365
rect 6269 3360 6795 3362
rect 6269 3304 6274 3360
rect 6330 3304 6734 3360
rect 6790 3304 6795 3360
rect 6269 3302 6795 3304
rect 6269 3299 6335 3302
rect 6729 3299 6795 3302
rect 3693 3226 3759 3229
rect 5441 3226 5507 3229
rect 3693 3224 5507 3226
rect 3693 3168 3698 3224
rect 3754 3168 5446 3224
rect 5502 3168 5507 3224
rect 3693 3166 5507 3168
rect 3693 3163 3759 3166
rect 5441 3163 5507 3166
rect 5809 3226 5875 3229
rect 6913 3226 6979 3229
rect 5809 3224 6979 3226
rect 5809 3168 5814 3224
rect 5870 3168 6918 3224
rect 6974 3168 6979 3224
rect 5809 3166 6979 3168
rect 5809 3163 5875 3166
rect 6913 3163 6979 3166
rect 3969 3090 4035 3093
rect 4889 3090 4955 3093
rect 5993 3090 6059 3093
rect 3969 3088 6059 3090
rect 3969 3032 3974 3088
rect 4030 3032 4894 3088
rect 4950 3032 5998 3088
rect 6054 3032 6059 3088
rect 3969 3030 6059 3032
rect 3969 3027 4035 3030
rect 4889 3027 4955 3030
rect 5993 3027 6059 3030
rect 11881 3090 11947 3093
rect 14825 3090 14891 3093
rect 11881 3088 14891 3090
rect 11881 3032 11886 3088
rect 11942 3032 14830 3088
rect 14886 3032 14891 3088
rect 11881 3030 14891 3032
rect 15150 3090 15210 3574
rect 22277 3362 22343 3365
rect 25200 3362 26000 3392
rect 22277 3360 26000 3362
rect 22277 3304 22282 3360
rect 22338 3304 26000 3360
rect 22277 3302 26000 3304
rect 22277 3299 22343 3302
rect 25200 3272 26000 3302
rect 16021 3090 16087 3093
rect 18045 3090 18111 3093
rect 15150 3088 18111 3090
rect 15150 3032 16026 3088
rect 16082 3032 18050 3088
rect 18106 3032 18111 3088
rect 15150 3030 18111 3032
rect 11881 3027 11947 3030
rect 14825 3027 14891 3030
rect 16021 3027 16087 3030
rect 18045 3027 18111 3030
rect 17125 2954 17191 2957
rect 19333 2954 19399 2957
rect 17125 2952 19399 2954
rect 17125 2896 17130 2952
rect 17186 2896 19338 2952
rect 19394 2896 19399 2952
rect 17125 2894 19399 2896
rect 17125 2891 17191 2894
rect 19333 2891 19399 2894
rect 11421 2818 11487 2821
rect 18781 2818 18847 2821
rect 19057 2818 19123 2821
rect 11421 2816 19123 2818
rect 11421 2760 11426 2816
rect 11482 2760 18786 2816
rect 18842 2760 19062 2816
rect 19118 2760 19123 2816
rect 11421 2758 19123 2760
rect 11421 2755 11487 2758
rect 18781 2755 18847 2758
rect 19057 2755 19123 2758
rect 4797 2682 4863 2685
rect 8109 2682 8175 2685
rect 4797 2680 8175 2682
rect 4797 2624 4802 2680
rect 4858 2624 8114 2680
rect 8170 2624 8175 2680
rect 4797 2622 8175 2624
rect 4797 2619 4863 2622
rect 8109 2619 8175 2622
rect 10869 2682 10935 2685
rect 18137 2682 18203 2685
rect 10869 2680 18203 2682
rect 10869 2624 10874 2680
rect 10930 2624 18142 2680
rect 18198 2624 18203 2680
rect 10869 2622 18203 2624
rect 10869 2619 10935 2622
rect 18137 2619 18203 2622
rect 7833 2546 7899 2549
rect 8845 2546 8911 2549
rect 7833 2544 8911 2546
rect 7833 2488 7838 2544
rect 7894 2488 8850 2544
rect 8906 2488 8911 2544
rect 7833 2486 8911 2488
rect 7833 2483 7899 2486
rect 8845 2483 8911 2486
rect 9857 2546 9923 2549
rect 12801 2546 12867 2549
rect 9857 2544 12867 2546
rect 9857 2488 9862 2544
rect 9918 2488 12806 2544
rect 12862 2488 12867 2544
rect 9857 2486 12867 2488
rect 9857 2483 9923 2486
rect 12801 2483 12867 2486
rect 15929 2546 15995 2549
rect 17953 2546 18019 2549
rect 15929 2544 18019 2546
rect 15929 2488 15934 2544
rect 15990 2488 17958 2544
rect 18014 2488 18019 2544
rect 15929 2486 18019 2488
rect 15929 2483 15995 2486
rect 17953 2483 18019 2486
rect 10409 2410 10475 2413
rect 12617 2410 12683 2413
rect 10409 2408 12683 2410
rect 10409 2352 10414 2408
rect 10470 2352 12622 2408
rect 12678 2352 12683 2408
rect 10409 2350 12683 2352
rect 10409 2347 10475 2350
rect 12617 2347 12683 2350
rect 16849 2410 16915 2413
rect 17401 2410 17467 2413
rect 16849 2408 17467 2410
rect 16849 2352 16854 2408
rect 16910 2352 17406 2408
rect 17462 2352 17467 2408
rect 16849 2350 17467 2352
rect 16849 2347 16915 2350
rect 17401 2347 17467 2350
rect 10041 2274 10107 2277
rect 10869 2274 10935 2277
rect 13537 2274 13603 2277
rect 10041 2272 13603 2274
rect 10041 2216 10046 2272
rect 10102 2216 10874 2272
rect 10930 2216 13542 2272
rect 13598 2216 13603 2272
rect 10041 2214 13603 2216
rect 10041 2211 10107 2214
rect 10869 2211 10935 2214
rect 13537 2211 13603 2214
rect 10685 1594 10751 1597
rect 12065 1594 12131 1597
rect 10685 1592 12131 1594
rect 10685 1536 10690 1592
rect 10746 1536 12070 1592
rect 12126 1536 12131 1592
rect 10685 1534 12131 1536
rect 10685 1531 10751 1534
rect 12065 1531 12131 1534
rect 5165 1458 5231 1461
rect 8017 1458 8083 1461
rect 9489 1458 9555 1461
rect 5165 1456 9555 1458
rect 5165 1400 5170 1456
rect 5226 1400 8022 1456
rect 8078 1400 9494 1456
rect 9550 1400 9555 1456
rect 5165 1398 9555 1400
rect 5165 1395 5231 1398
rect 8017 1395 8083 1398
rect 9489 1395 9555 1398
rect 10869 1458 10935 1461
rect 12065 1458 12131 1461
rect 10869 1456 12131 1458
rect 10869 1400 10874 1456
rect 10930 1400 12070 1456
rect 12126 1400 12131 1456
rect 10869 1398 12131 1400
rect 10869 1395 10935 1398
rect 12065 1395 12131 1398
rect 11053 1322 11119 1325
rect 13169 1322 13235 1325
rect 11053 1320 13235 1322
rect 11053 1264 11058 1320
rect 11114 1264 13174 1320
rect 13230 1264 13235 1320
rect 11053 1262 13235 1264
rect 11053 1259 11119 1262
rect 13169 1259 13235 1262
rect 0 1186 800 1216
rect 6361 1186 6427 1189
rect 0 1184 6427 1186
rect 0 1128 6366 1184
rect 6422 1128 6427 1184
rect 0 1126 6427 1128
rect 0 1096 800 1126
rect 6361 1123 6427 1126
rect 21817 1186 21883 1189
rect 25200 1186 26000 1216
rect 21817 1184 26000 1186
rect 21817 1128 21822 1184
rect 21878 1128 26000 1184
rect 21817 1126 26000 1128
rect 21817 1123 21883 1126
rect 25200 1096 26000 1126
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1562557784
transform -1 0 19044 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _364_
timestamp 21601
transform -1 0 16100 0 1 1088
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _365_
timestamp 1562557784
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _366_
timestamp 1562557784
transform -1 0 2208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _367_
timestamp 1562557784
transform -1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _368_
timestamp 1562557784
transform -1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _369_
timestamp 1562557784
transform 1 0 12236 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _370_
timestamp 1562557784
transform 1 0 11040 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _371_
timestamp 1562557784
transform -1 0 13064 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _372_
timestamp 1562557784
transform -1 0 2852 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__inv_12  _373_
timestamp 21601
transform 1 0 22080 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _374_
timestamp 21601
transform -1 0 19044 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _375_
timestamp 21601
transform -1 0 19044 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _376_
timestamp 21601
transform 1 0 21896 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _377_
timestamp 21601
transform 1 0 18032 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_4  _378_
timestamp 21601
transform 1 0 15456 0 1 5440
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_1  _379_
timestamp 21601
transform -1 0 15272 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_2  _380_
timestamp 21601
transform 1 0 14812 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _381_
timestamp 21601
transform -1 0 15916 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_1  _382_
timestamp 21601
transform -1 0 12144 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _383_
timestamp 21601
transform 1 0 12052 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _384_
timestamp 21601
transform -1 0 11776 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _385_
timestamp 21601
transform 1 0 15456 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _386_
timestamp 21601
transform 1 0 14168 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _387_
timestamp 21601
transform 1 0 14260 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _388_
timestamp 21601
transform -1 0 13800 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_2  _389_
timestamp 21601
transform -1 0 13984 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_4  _390_
timestamp 21601
transform 1 0 9016 0 1 6528
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_1  _391_
timestamp 21601
transform -1 0 10672 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21boi_2  _392_
timestamp 21601
transform -1 0 10028 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_1  _393_
timestamp 21601
transform 1 0 9568 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _394_
timestamp 21601
transform 1 0 11224 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _395_
timestamp 21601
transform 1 0 9016 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3b_1  _396_
timestamp 21601
transform 1 0 10580 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _397_
timestamp 21601
transform 1 0 10212 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _398_
timestamp 21601
transform 1 0 11592 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _399_
timestamp 21601
transform 1 0 5704 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _400_
timestamp 21601
transform 1 0 6440 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _401_
timestamp 21601
transform -1 0 6992 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _402_
timestamp 21601
transform 1 0 6440 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _403_
timestamp 21601
transform -1 0 9016 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _404_
timestamp 21601
transform -1 0 8740 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _405_
timestamp 21601
transform -1 0 7912 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _406_
timestamp 21601
transform -1 0 8740 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _407_
timestamp 1562557784
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _408_
timestamp 21601
transform 1 0 2300 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_2  _409_
timestamp 21601
transform 1 0 3864 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _410_
timestamp 21601
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_1  _411_
timestamp 21601
transform -1 0 3956 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_4  _412_
timestamp 21601
transform -1 0 5796 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3b_1  _413_
timestamp 21601
transform -1 0 5520 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _414_
timestamp 21601
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _415_
timestamp 21601
transform 1 0 6348 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _416_
timestamp 21601
transform 1 0 5428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _417_
timestamp 21601
transform -1 0 5152 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o21bai_4  _418_
timestamp 21601
transform 1 0 2852 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__nand3_2  _419_
timestamp 21601
transform 1 0 1932 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o2bb2ai_4  _420_
timestamp 21601
transform -1 0 3496 0 1 5440
box -38 -48 2062 592
use sky130_fd_sc_hd__nand3_4  _421_
timestamp 21601
transform -1 0 3680 0 -1 5440
box -38 -48 1326 592
use sky130_fd_sc_hd__and2b_1  _422_
timestamp 21601
transform 1 0 1656 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _423_
timestamp 21601
transform -1 0 4232 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _424_
timestamp 21601
transform -1 0 4692 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__o211ai_4  _425_
timestamp 21601
transform 1 0 4600 0 -1 5440
box -38 -48 1602 592
use sky130_fd_sc_hd__a32oi_2  _426_
timestamp 21601
transform 1 0 6808 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_4  _427_
timestamp 21601
transform -1 0 8924 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__o22ai_2  _428_
timestamp 21601
transform -1 0 11040 0 -1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o211ai_2  _429_
timestamp 21601
transform -1 0 11040 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _430_
timestamp 21601
transform 1 0 13156 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _431_
timestamp 21601
transform -1 0 16468 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _432_
timestamp 21601
transform -1 0 11868 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _433_
timestamp 21601
transform 1 0 13800 0 -1 4352
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _434_
timestamp 21601
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _435_
timestamp 21601
transform -1 0 19596 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _436_
timestamp 21601
transform -1 0 15640 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_2  _437_
timestamp 21601
transform 1 0 14628 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _438_
timestamp 21601
transform -1 0 14444 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_2  _439_
timestamp 21601
transform -1 0 5428 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nand3b_1  _440_
timestamp 21601
transform -1 0 8740 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _441_
timestamp 21601
transform 1 0 4048 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _442_
timestamp 21601
transform 1 0 4508 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _443_
timestamp 21601
transform -1 0 16468 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _444_
timestamp 21601
transform 1 0 15824 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o2111ai_1  _445_
timestamp 21601
transform -1 0 16192 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _446_
timestamp 21601
transform 1 0 17480 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _447_
timestamp 21601
transform -1 0 17020 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _448_
timestamp 21601
transform -1 0 16100 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _449_
timestamp 21601
transform 1 0 15824 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _450_
timestamp 21601
transform -1 0 15272 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _451_
timestamp 21601
transform 1 0 12328 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _452_
timestamp 21601
transform 1 0 12236 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _453_
timestamp 21601
transform 1 0 9016 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _454_
timestamp 21601
transform 1 0 10488 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _455_
timestamp 21601
transform -1 0 10304 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _456_
timestamp 21601
transform -1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _457_
timestamp 21601
transform 1 0 6808 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _458_
timestamp 21601
transform 1 0 6716 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _459_
timestamp 21601
transform -1 0 5704 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _460_
timestamp 21601
transform -1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _461_
timestamp 21601
transform 1 0 5888 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _462_
timestamp 21601
transform 1 0 5060 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _463_
timestamp 21601
transform 1 0 1840 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o2111ai_1  _464_
timestamp 21601
transform 1 0 2576 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _465_
timestamp 21601
transform -1 0 4876 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _466_
timestamp 21601
transform 1 0 2576 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _467_
timestamp 21601
transform -1 0 3036 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _468_
timestamp 21601
transform 1 0 2116 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _469_
timestamp 21601
transform 1 0 19320 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 21601
transform 1 0 22540 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _471_
timestamp 21601
transform 1 0 20240 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _472_
timestamp 21601
transform 1 0 2668 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _473_
timestamp 21601
transform 1 0 7912 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _474_
timestamp 21601
transform 1 0 4692 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _475_
timestamp 21601
transform 1 0 22080 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _476_
timestamp 21601
transform 1 0 18216 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _477_
timestamp 21601
transform -1 0 22724 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _478_
timestamp 21601
transform 1 0 2392 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _479_
timestamp 21601
transform -1 0 6256 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _480_
timestamp 21601
transform 1 0 2208 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _481_
timestamp 21601
transform 1 0 17572 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _482_
timestamp 21601
transform 1 0 20332 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _483_
timestamp 21601
transform 1 0 19320 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _484_
timestamp 21601
transform 1 0 3864 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _485_
timestamp 21601
transform 1 0 7820 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _486_
timestamp 21601
transform 1 0 4324 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _487_
timestamp 21601
transform 1 0 22816 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _488_
timestamp 21601
transform 1 0 20608 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _489_
timestamp 21601
transform 1 0 22908 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _490_
timestamp 21601
transform 1 0 2392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _491_
timestamp 21601
transform 1 0 5980 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _492_
timestamp 21601
transform 1 0 2300 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _493_
timestamp 21601
transform 1 0 5704 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _494_
timestamp 21601
transform -1 0 8372 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _495_
timestamp 21601
transform -1 0 7728 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _496_
timestamp 21601
transform 1 0 6900 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _497_
timestamp 21601
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _498_
timestamp 21601
transform -1 0 9752 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _499_
timestamp 21601
transform -1 0 7268 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _500_
timestamp 21601
transform -1 0 6808 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _501_
timestamp 21601
transform -1 0 7728 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _502_
timestamp 21601
transform 1 0 6164 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _503_
timestamp 21601
transform 1 0 6440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _504_
timestamp 21601
transform 1 0 5244 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _505_
timestamp 21601
transform 1 0 8188 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _506_
timestamp 21601
transform 1 0 6440 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _507_
timestamp 21601
transform 1 0 5336 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _508_
timestamp 21601
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _509_
timestamp 21601
transform 1 0 6992 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _510_
timestamp 21601
transform 1 0 20516 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _511_
timestamp 21601
transform -1 0 23828 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _512_
timestamp 21601
transform 1 0 21896 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _513_
timestamp 21601
transform 1 0 2484 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _514_
timestamp 21601
transform 1 0 8464 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _515_
timestamp 21601
transform 1 0 4876 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _516_
timestamp 21601
transform 1 0 14628 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _517_
timestamp 21601
transform 1 0 17296 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _518_
timestamp 21601
transform 1 0 16744 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _519_
timestamp 21601
transform 1 0 5336 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _520_
timestamp 21601
transform 1 0 7360 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _521_
timestamp 21601
transform 1 0 2484 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _522_
timestamp 21601
transform 1 0 23092 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _523_
timestamp 21601
transform -1 0 20240 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _524_
timestamp 21601
transform 1 0 23000 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _525_
timestamp 21601
transform 1 0 2484 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _526_
timestamp 21601
transform -1 0 7912 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _527_
timestamp 21601
transform 1 0 2484 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _528_
timestamp 21601
transform 1 0 16744 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _529_
timestamp 21601
transform -1 0 19596 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _530_
timestamp 21601
transform 1 0 17756 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _531_
timestamp 21601
transform 1 0 6900 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _532_
timestamp 21601
transform 1 0 7820 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _533_
timestamp 21601
transform 1 0 3864 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_2  _534_
timestamp 21601
transform -1 0 12696 0 1 1088
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _535_
timestamp 21601
transform -1 0 10488 0 -1 3264
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2_1  _536_
timestamp 21601
transform 1 0 7728 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _537_
timestamp 21601
transform -1 0 14996 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _538_
timestamp 21601
transform -1 0 9476 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _539_
timestamp 21601
transform -1 0 12788 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _540_
timestamp 21601
transform 1 0 10028 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_2  _541_
timestamp 21601
transform -1 0 12512 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o221ai_4  _542_
timestamp 21601
transform 1 0 12696 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_2  _543_
timestamp 21601
transform -1 0 15364 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _544_
timestamp 21601
transform 1 0 10672 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_2  _545_
timestamp 21601
transform 1 0 12236 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__a41oi_4  _546_
timestamp 21601
transform -1 0 13708 0 1 2176
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2b_4  _547_
timestamp 21601
transform 1 0 12880 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__nand4b_4  _548_
timestamp 21601
transform 1 0 9384 0 1 1088
box -38 -48 1786 592
use sky130_fd_sc_hd__nor3_4  _549_
timestamp 21601
transform 1 0 10304 0 1 2176
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _550_
timestamp 21601
transform 1 0 5612 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__nand2b_4  _551_
timestamp 21601
transform -1 0 7912 0 1 1088
box -38 -48 1050 592
use sky130_fd_sc_hd__nand2b_1  _552_
timestamp 21601
transform 1 0 4968 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _553_
timestamp 21601
transform -1 0 6164 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _554_
timestamp 21601
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand4b_4  _555_
timestamp 21601
transform -1 0 7544 0 1 2176
box -38 -48 1786 592
use sky130_fd_sc_hd__nand2b_1  _556_
timestamp 21601
transform -1 0 4324 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _557_
timestamp 21601
transform -1 0 3496 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _558_
timestamp 21601
transform -1 0 4048 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _559_
timestamp 21601
transform -1 0 4784 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _560_
timestamp 21601
transform 1 0 2944 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_4  _561_
timestamp 21601
transform -1 0 7912 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_2  _562_
timestamp 21601
transform 1 0 13156 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2ai_4  _563_
timestamp 21601
transform 1 0 10672 0 1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_8  _564_
timestamp 21601
transform 1 0 15272 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _565_
timestamp 21601
transform -1 0 12328 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _566_
timestamp 21601
transform -1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _567_
timestamp 21601
transform 1 0 10856 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_4  _568_
timestamp 21601
transform -1 0 12420 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _569_
timestamp 21601
transform -1 0 10304 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o211ai_2  _570_
timestamp 21601
transform 1 0 11592 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _571_
timestamp 21601
transform 1 0 9752 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _572_
timestamp 21601
transform 1 0 15640 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _573_
timestamp 1562557784
transform -1 0 14076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _574_
timestamp 21601
transform -1 0 13432 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _575_
timestamp 21601
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _576_
timestamp 21601
transform 1 0 10488 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__nand3_2  _577_
timestamp 21601
transform -1 0 10948 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_2  _578_
timestamp 21601
transform 1 0 9476 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _579_
timestamp 21601
transform -1 0 12052 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__nand3_2  _580_
timestamp 21601
transform 1 0 13156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _581_
timestamp 21601
transform -1 0 15824 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _582_
timestamp 21601
transform 1 0 16284 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _583_
timestamp 21601
transform 1 0 15640 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _584_
timestamp 21601
transform -1 0 15824 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _585_
timestamp 21601
transform 1 0 13064 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _586_
timestamp 21601
transform -1 0 11960 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_4  _587_
timestamp 21601
transform 1 0 11684 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_2  _588_
timestamp 21601
transform 1 0 19688 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _589_
timestamp 21601
transform -1 0 13616 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _590_
timestamp 21601
transform -1 0 13800 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_8  _591_
timestamp 21601
transform 1 0 13248 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_1  _592_
timestamp 21601
transform -1 0 6808 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__nand4b_4  _593_
timestamp 21601
transform -1 0 5612 0 1 2176
box -38 -48 1786 592
use sky130_fd_sc_hd__and4b_1  _594_
timestamp 21601
transform -1 0 11316 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand4b_4  _595_
timestamp 21601
transform -1 0 12972 0 1 9792
box -38 -48 1786 592
use sky130_fd_sc_hd__o31a_1  _596_
timestamp 21601
transform -1 0 15088 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _597_
timestamp 21601
transform 1 0 13800 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _598_
timestamp 21601
transform -1 0 15180 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _599_
timestamp 21601
transform 1 0 14352 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _600_
timestamp 21601
transform -1 0 15456 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _601_
timestamp 21601
transform 1 0 15640 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_1  _602_
timestamp 21601
transform 1 0 16008 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _603_
timestamp 21601
transform -1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _604_
timestamp 21601
transform -1 0 15640 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_1  _605_
timestamp 21601
transform 1 0 14352 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a31oi_1  _606_
timestamp 21601
transform 1 0 16008 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _607_
timestamp 21601
transform -1 0 12144 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_1  _608_
timestamp 21601
transform 1 0 13248 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _609_
timestamp 21601
transform 1 0 12236 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _610_
timestamp 21601
transform -1 0 10672 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _611_
timestamp 21601
transform -1 0 9384 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__or3b_4  _612_
timestamp 21601
transform 1 0 10304 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _613_
timestamp 21601
transform -1 0 10120 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_1  _614_
timestamp 21601
transform -1 0 10672 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _615_
timestamp 21601
transform 1 0 10488 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a41o_1  _616_
timestamp 21601
transform 1 0 9568 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o31ai_1  _617_
timestamp 21601
transform -1 0 9936 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _618_
timestamp 21601
transform 1 0 13432 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _619_
timestamp 21601
transform -1 0 13892 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _620_
timestamp 21601
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _621_
timestamp 21601
transform 1 0 12696 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _622_
timestamp 21601
transform -1 0 14996 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _623_
timestamp 21601
transform 1 0 12604 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _624_
timestamp 21601
transform 1 0 12144 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _625_
timestamp 21601
transform 1 0 14720 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _626_
timestamp 21601
transform -1 0 16100 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _627_
timestamp 21601
transform 1 0 12512 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _628_
timestamp 21601
transform 1 0 16560 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _629_
timestamp 21601
transform 1 0 16744 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _630_
timestamp 21601
transform -1 0 14904 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _631_
timestamp 21601
transform 1 0 11684 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _632_
timestamp 21601
transform 1 0 10672 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a211oi_4  _633_
timestamp 21601
transform -1 0 14352 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__a32o_1  _634_
timestamp 21601
transform -1 0 13248 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _635_
timestamp 21601
transform -1 0 12052 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_4  _636_
timestamp 21601
transform -1 0 10856 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_1  _637_
timestamp 21601
transform 1 0 11592 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _638_
timestamp 21601
transform 1 0 16928 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _639_
timestamp 21601
transform 1 0 16744 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_2  _640_
timestamp 21601
transform -1 0 10488 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_2  _641_
timestamp 21601
transform -1 0 11316 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _642_
timestamp 21601
transform 1 0 14444 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _643_
timestamp 21601
transform -1 0 15456 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__o311a_1  _644_
timestamp 21601
transform -1 0 16008 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_2  _645_
timestamp 21601
transform 1 0 13432 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__o41a_1  _646_
timestamp 21601
transform 1 0 10396 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _647_
timestamp 21601
transform 1 0 10212 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _648_
timestamp 21601
transform -1 0 13524 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _649_
timestamp 21601
transform -1 0 10856 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _650_
timestamp 21601
transform 1 0 9476 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _651_
timestamp 21601
transform 1 0 13524 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _652_
timestamp 21601
transform -1 0 10488 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _653_
timestamp 21601
transform 1 0 15364 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _654_
timestamp 21601
transform 1 0 16008 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _655_
timestamp 21601
transform 1 0 16008 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _656_
timestamp 21601
transform -1 0 21528 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _657_
timestamp 21601
transform 1 0 15088 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_1  _658_
timestamp 21601
transform -1 0 16836 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _659_
timestamp 21601
transform 1 0 15088 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _660_
timestamp 21601
transform 1 0 19596 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _661_
timestamp 21601
transform -1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _662_
timestamp 21601
transform 1 0 19596 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _663_
timestamp 21601
transform -1 0 21528 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _664_
timestamp 21601
transform -1 0 20608 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _665_
timestamp 21601
transform 1 0 20056 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _666_
timestamp 21601
transform 1 0 20884 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_4  _667_
timestamp 21601
transform -1 0 22264 0 1 15232
box -38 -48 1326 592
use sky130_fd_sc_hd__a21o_1  _668_
timestamp 21601
transform 1 0 21712 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _669_
timestamp 21601
transform 1 0 16008 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _670_
timestamp 21601
transform 1 0 19964 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _671_
timestamp 21601
transform -1 0 21160 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _672_
timestamp 21601
transform 1 0 21620 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _673_
timestamp 21601
transform 1 0 21896 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _674_
timestamp 21601
transform -1 0 21528 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _675_
timestamp 21601
transform -1 0 24196 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _676_
timestamp 21601
transform 1 0 20976 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _677_
timestamp 21601
transform 1 0 21896 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _678_
timestamp 21601
transform -1 0 24472 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _679_
timestamp 21601
transform -1 0 15640 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _680_
timestamp 21601
transform 1 0 14260 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _681_
timestamp 21601
transform 1 0 8924 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _682_
timestamp 21601
transform 1 0 9108 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _683_
timestamp 21601
transform 1 0 18124 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _684_
timestamp 21601
transform 1 0 17480 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _685_
timestamp 21601
transform 1 0 16928 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _686_
timestamp 21601
transform 1 0 17572 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _687_
timestamp 21601
transform 1 0 3588 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _688_
timestamp 21601
transform -1 0 9568 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _689_
timestamp 21601
transform -1 0 6900 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _690_
timestamp 21601
transform -1 0 19228 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _691_
timestamp 21601
transform 1 0 19320 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _692_
timestamp 21601
transform -1 0 18676 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _693_
timestamp 21601
transform 1 0 2300 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _694_
timestamp 21601
transform 1 0 6440 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _695_
timestamp 21601
transform 1 0 1840 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _696_
timestamp 21601
transform 1 0 23092 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _697_
timestamp 21601
transform 1 0 17572 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _698_
timestamp 21601
transform -1 0 24472 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _699_
timestamp 21601
transform 1 0 1840 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _700_
timestamp 21601
transform -1 0 9568 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _701_
timestamp 21601
transform 1 0 5704 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _702_
timestamp 21601
transform -1 0 18768 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _703_
timestamp 21601
transform 1 0 17572 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _704_
timestamp 21601
transform 1 0 14904 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _705_
timestamp 21601
transform -1 0 6164 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _706_
timestamp 21601
transform -1 0 8556 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _707_
timestamp 21601
transform 1 0 1840 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _708_
timestamp 21601
transform 1 0 22356 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _709_
timestamp 21601
transform 1 0 21160 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _710_
timestamp 21601
transform 1 0 20976 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _711_
timestamp 21601
transform 1 0 4140 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _712_
timestamp 21601
transform 1 0 4692 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _713_
timestamp 21601
transform 1 0 4600 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _714_
timestamp 21601
transform 1 0 8188 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _715_
timestamp 21601
transform -1 0 13248 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _716_
timestamp 21601
transform 1 0 7544 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _717_
timestamp 21601
transform 1 0 1840 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _718_
timestamp 21601
transform 1 0 5612 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _719_
timestamp 21601
transform 1 0 1748 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _720_
timestamp 21601
transform -1 0 24472 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _721_
timestamp 21601
transform -1 0 22356 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _722_
timestamp 21601
transform -1 0 24472 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _723_
timestamp 21601
transform -1 0 5796 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _724_
timestamp 21601
transform 1 0 7176 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _725_
timestamp 21601
transform -1 0 4140 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _726_
timestamp 21601
transform -1 0 20792 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _727_
timestamp 21601
transform 1 0 19688 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _728_
timestamp 21601
transform -1 0 19044 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _729_
timestamp 21601
transform 1 0 21160 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _730_
timestamp 21601
transform 1 0 22172 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _731_
timestamp 21601
transform 1 0 17940 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _732_
timestamp 21601
transform 1 0 2116 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _733_
timestamp 21601
transform -1 0 6900 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _734_
timestamp 21601
transform 1 0 1656 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _735_
timestamp 21601
transform -1 0 24472 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _736_
timestamp 21601
transform -1 0 19504 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _737_
timestamp 21601
transform -1 0 21436 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _738_
timestamp 21601
transform 1 0 4048 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _739_
timestamp 21601
transform 1 0 8096 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _740_
timestamp 21601
transform 1 0 2024 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _741_
timestamp 21601
transform -1 0 22356 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _742_
timestamp 21601
transform -1 0 24196 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _743_
timestamp 21601
transform -1 0 21620 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _744_
timestamp 21601
transform -1 0 2392 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _745_
timestamp 21601
transform 1 0 1932 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _746_
timestamp 21601
transform 1 0 5612 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _747_
timestamp 21601
transform 1 0 6992 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _748_
timestamp 21601
transform -1 0 15272 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _749_
timestamp 21601
transform -1 0 16008 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _750_
timestamp 21601
transform 1 0 16652 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _751_
timestamp 21601
transform 1 0 16836 0 1 1088
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _752_
timestamp 21601
transform 1 0 4968 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__dfrtp_2  _753_
timestamp 21601
transform 1 0 14168 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _754_
timestamp 21601
transform 1 0 14168 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _755_
timestamp 21601
transform 1 0 9016 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _756_
timestamp 21601
transform 1 0 8188 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _757_
timestamp 21601
transform 1 0 17204 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _758_
timestamp 21601
transform 1 0 16652 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _759_
timestamp 21601
transform 1 0 16744 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _760_
timestamp 21601
transform 1 0 17020 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _761_
timestamp 21601
transform 1 0 2944 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _762_
timestamp 21601
transform 1 0 7084 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _763_
timestamp 21601
transform -1 0 6716 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _764_
timestamp 21601
transform 1 0 16928 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _765_
timestamp 21601
transform 1 0 18952 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _766_
timestamp 21601
transform 1 0 16192 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _767_
timestamp 21601
transform 1 0 1564 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _768_
timestamp 21601
transform -1 0 8280 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _769_
timestamp 21601
transform 1 0 1656 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _770_
timestamp 21601
transform 1 0 22540 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _771_
timestamp 21601
transform 1 0 19780 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _772_
timestamp 21601
transform 1 0 21988 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _773_
timestamp 21601
transform 1 0 1564 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _774_
timestamp 21601
transform 1 0 7084 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _775_
timestamp 21601
transform 1 0 4876 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _776_
timestamp 21601
transform 1 0 16284 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _777_
timestamp 21601
transform 1 0 16928 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _778_
timestamp 21601
transform 1 0 14168 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _779_
timestamp 21601
transform 1 0 4324 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _780_
timestamp 21601
transform -1 0 8740 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _781_
timestamp 21601
transform 1 0 1656 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _782_
timestamp 21601
transform 1 0 21620 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _783_
timestamp 21601
transform -1 0 24380 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _784_
timestamp 21601
transform 1 0 20056 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _785_
timestamp 21601
transform -1 0 5980 0 1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _786_
timestamp 21601
transform -1 0 6164 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _787_
timestamp 21601
transform 1 0 4232 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _788_
timestamp 21601
transform 1 0 7452 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _789_
timestamp 21601
transform 1 0 9200 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _790_
timestamp 21601
transform 1 0 6624 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _791_
timestamp 21601
transform 1 0 1472 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _792_
timestamp 21601
transform 1 0 4968 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _793_
timestamp 21601
transform 1 0 1564 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _794_
timestamp 21601
transform 1 0 21988 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _795_
timestamp 21601
transform 1 0 19780 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _796_
timestamp 21601
transform 1 0 22356 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _797_
timestamp 21601
transform 1 0 3864 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _798_
timestamp 21601
transform 1 0 7084 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _799_
timestamp 21601
transform 1 0 2300 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _800_
timestamp 21601
transform 1 0 19320 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _801_
timestamp 21601
transform 1 0 19964 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _802_
timestamp 21601
transform 1 0 17112 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _803_
timestamp 21601
transform -1 0 23828 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _804_
timestamp 21601
transform -1 0 24196 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _805_
timestamp 21601
transform -1 0 20700 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _806_
timestamp 21601
transform 1 0 1472 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _807_
timestamp 21601
transform -1 0 6164 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _808_
timestamp 21601
transform 1 0 1472 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _809_
timestamp 21601
transform 1 0 22264 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _810_
timestamp 21601
transform -1 0 19044 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _811_
timestamp 21601
transform -1 0 21712 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _812_
timestamp 21601
transform 1 0 3956 0 -1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _813_
timestamp 21601
transform 1 0 7176 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _814_
timestamp 21601
transform 1 0 1472 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _815_
timestamp 21601
transform 1 0 19688 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _816_
timestamp 21601
transform 1 0 22172 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _817_
timestamp 21601
transform 1 0 19136 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _818_
timestamp 21601
transform -1 0 3312 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _819_
timestamp 21601
transform 1 0 1656 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _820_
timestamp 21601
transform 1 0 4876 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _821_
timestamp 21601
transform 1 0 6624 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _822_
timestamp 21601
transform 1 0 9016 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _823_
timestamp 21601
transform 1 0 11776 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _824_
timestamp 21601
transform 1 0 16744 0 -1 4352
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _825_
timestamp 21601
transform 1 0 16744 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _826_
timestamp 21601
transform 1 0 7728 0 -1 2176
box -38 -48 2154 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 21601
transform -1 0 16468 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 21601
transform -1 0 3588 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 21601
transform -1 0 4048 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 21601
transform -1 0 3588 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 21601
transform -1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 21601
transform -1 0 6164 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 21601
transform -1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 21601
transform -1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 21601
transform -1 0 12972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 21601
transform -1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 21601
transform -1 0 6164 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 21601
transform -1 0 4600 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 21601
transform -1 0 7176 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 21601
transform -1 0 9752 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 21601
transform -1 0 17664 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 21601
transform -1 0 19044 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 21601
transform -1 0 21160 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 21601
transform -1 0 14628 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 21601
transform -1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 21601
transform -1 0 17664 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 21601
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 21601
transform -1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 21601
transform -1 0 24196 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 21601
transform -1 0 24196 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 21601
transform -1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 21601
transform -1 0 24472 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 21601
transform -1 0 19044 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 21601
transform -1 0 21712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 21601
transform -1 0 1656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 21601
transform -1 0 3588 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 21601
transform -1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 21601
transform -1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 21601
transform -1 0 1656 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 21601
transform -1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 21601
transform -1 0 3588 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 21601
transform -1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 21601
transform -1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 21601
transform -1 0 16928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_0
timestamp 21601
transform 1 0 9200 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clockp_buffer_1
timestamp 21601
transform 1 0 19320 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__and2_2  clone1
timestamp 21601
transform 1 0 21712 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__inv_6  clone3
timestamp 21601
transform -1 0 7820 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_4  fanout39
timestamp 21601
transform -1 0 16376 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout40
timestamp 21601
transform -1 0 8464 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout41
timestamp 21601
transform -1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout42
timestamp 21601
transform -1 0 11592 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout43
timestamp 21601
transform 1 0 23460 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout44
timestamp 21601
transform 1 0 21988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout45
timestamp 21601
transform 1 0 20424 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout46
timestamp 21601
transform -1 0 16376 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  fanout47
timestamp 21601
transform 1 0 23920 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout48
timestamp 21601
transform -1 0 4508 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  fanout49
timestamp 21601
transform -1 0 10028 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  fanout51
timestamp 21601
transform 1 0 18216 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout52
timestamp 21601
transform -1 0 16468 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  fanout53
timestamp 21601
transform -1 0 20884 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  fanout54
timestamp 21601
transform 1 0 4784 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout55
timestamp 21601
transform -1 0 9936 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout56
timestamp 21601
transform -1 0 7544 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout57
timestamp 21601
transform 1 0 16652 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout58
timestamp 21601
transform -1 0 16836 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout59
timestamp 21601
transform -1 0 19872 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout60
timestamp 21601
transform 1 0 4324 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout61
timestamp 21601
transform -1 0 8740 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  fanout62
timestamp 21601
transform -1 0 8740 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout63
timestamp 21601
transform 1 0 19228 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout64
timestamp 21601
transform -1 0 17388 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout65
timestamp 21601
transform -1 0 19688 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  fanout66
timestamp 21601
transform -1 0 17296 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  fanout67
timestamp 21601
transform 1 0 18216 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3
timestamp 21601
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7
timestamp 21601
transform 1 0 1748 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14
timestamp 21601
transform 1 0 2392 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19
timestamp 21601
transform 1 0 2852 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26
timestamp 21601
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 21601
transform 1 0 3772 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35
timestamp 21601
transform 1 0 4324 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 21601
transform 1 0 4784 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47
timestamp 21601
transform 1 0 5428 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 21601
transform 1 0 6164 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57
timestamp 21601
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61
timestamp 21601
transform 1 0 6716 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_74
timestamp 21601
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 21601
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_85
timestamp 21601
transform 1 0 8924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_88
timestamp 21601
transform 1 0 9200 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 21601
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_113
timestamp 21601
transform 1 0 11500 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_117
timestamp 21601
transform 1 0 11868 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_126
timestamp 21601
transform 1 0 12696 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 21601
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_141
timestamp 21601
transform 1 0 14076 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_152
timestamp 21601
transform 1 0 15088 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_163
timestamp 21601
transform 1 0 16100 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_166
timestamp 21601
transform 1 0 16376 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 21601
transform 1 0 16652 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 21601
transform 1 0 17296 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_181
timestamp 21601
transform 1 0 17756 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_188
timestamp 21601
transform 1 0 18400 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 21601
transform 1 0 19044 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 21601
transform 1 0 19228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_201
timestamp 21601
transform 1 0 19596 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 21601
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_225
timestamp 21601
transform 1 0 21804 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_229
timestamp 21601
transform 1 0 22172 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 21601
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 21601
transform 1 0 24380 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_3
timestamp 21601
transform 1 0 1380 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_24
timestamp 21601
transform 1 0 3312 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_32
timestamp 21601
transform 1 0 4048 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_40
timestamp 21601
transform 1 0 4784 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_47
timestamp 21601
transform 1 0 5428 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 21601
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 21601
transform 1 0 6348 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_62
timestamp 21601
transform 1 0 6808 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_70
timestamp 21601
transform 1 0 7544 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_95
timestamp 21601
transform 1 0 9844 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_102
timestamp 21601
transform 1 0 10488 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 21601
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 21601
transform 1 0 11500 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_116
timestamp 21601
transform 1 0 11776 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_124
timestamp 21601
transform 1 0 12512 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_147
timestamp 21601
transform 1 0 14628 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_154
timestamp 21601
transform 1 0 15272 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_157
timestamp 21601
transform 1 0 15548 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_166
timestamp 21601
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_169
timestamp 21601
transform 1 0 16652 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_191
timestamp 21601
transform 1 0 18676 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_1_213
timestamp 21601
transform 1 0 20700 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_216
timestamp 21601
transform 1 0 20976 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 21601
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_225
timestamp 21601
transform 1 0 21804 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_1_247
timestamp 21601
transform 1 0 23828 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_254
timestamp 21601
transform 1 0 24472 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 21601
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_9
timestamp 21601
transform 1 0 1932 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_18
timestamp 21601
transform 1 0 2760 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 21601
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_29
timestamp 21601
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_49
timestamp 21601
transform 1 0 5612 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_70
timestamp 21601
transform 1 0 7544 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_75
timestamp 21601
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 21601
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_85
timestamp 21601
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_89
timestamp 21601
transform 1 0 9292 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_98
timestamp 21601
transform 1 0 10120 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_113
timestamp 21601
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_137
timestamp 21601
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_141
timestamp 21601
transform 1 0 14076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_155
timestamp 21601
transform 1 0 15364 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_164
timestamp 21601
transform 1 0 16192 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_173
timestamp 21601
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_182
timestamp 21601
transform 1 0 17848 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_187
timestamp 21601
transform 1 0 18308 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 21601
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_197
timestamp 21601
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_208
timestamp 21601
transform 1 0 20240 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_226
timestamp 21601
transform 1 0 21896 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_241
timestamp 21601
transform 1 0 23276 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_2_249
timestamp 21601
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 21601
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_3
timestamp 21601
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_3_6
timestamp 21601
transform 1 0 1656 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_10
timestamp 21601
transform 1 0 2024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_15
timestamp 21601
transform 1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_21
timestamp 21601
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_24
timestamp 21601
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_30
timestamp 21601
transform 1 0 3864 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_35
timestamp 21601
transform 1 0 4324 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_40
timestamp 21601
transform 1 0 4784 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_47
timestamp 21601
transform 1 0 5428 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_54
timestamp 21601
transform 1 0 6072 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_57
timestamp 21601
transform 1 0 6348 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 21601
transform 1 0 7912 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_3_79
timestamp 21601
transform 1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_89
timestamp 21601
transform 1 0 9292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_102
timestamp 21601
transform 1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 21601
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 21601
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_119
timestamp 21601
transform 1 0 12052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_130
timestamp 21601
transform 1 0 13064 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_145
timestamp 21601
transform 1 0 14444 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_155
timestamp 21601
transform 1 0 15364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_163
timestamp 21601
transform 1 0 16100 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 21601
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_169
timestamp 21601
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_177
timestamp 21601
transform 1 0 17388 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_184
timestamp 21601
transform 1 0 18032 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_195
timestamp 21601
transform 1 0 19044 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_201
timestamp 21601
transform 1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 21601
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_225
timestamp 21601
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_231
timestamp 21601
transform 1 0 22356 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_253
timestamp 21601
transform 1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_3
timestamp 21601
transform 1 0 1380 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_7
timestamp 21601
transform 1 0 1748 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_14
timestamp 21601
transform 1 0 2392 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_23
timestamp 21601
transform 1 0 3220 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 21601
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_29
timestamp 21601
transform 1 0 3772 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_34
timestamp 21601
transform 1 0 4232 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_39
timestamp 21601
transform 1 0 4692 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_61
timestamp 21601
transform 1 0 6716 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_4_69
timestamp 21601
transform 1 0 7452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_77
timestamp 21601
transform 1 0 8188 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 21601
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_85
timestamp 21601
transform 1 0 8924 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_106
timestamp 21601
transform 1 0 10856 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_114
timestamp 21601
transform 1 0 11592 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_126
timestamp 21601
transform 1 0 12696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 21601
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_141
timestamp 21601
transform 1 0 14076 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_151
timestamp 21601
transform 1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_158
timestamp 21601
transform 1 0 15640 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_167
timestamp 21601
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_173
timestamp 21601
transform 1 0 17020 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 21601
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_197
timestamp 21601
transform 1 0 19228 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_205
timestamp 21601
transform 1 0 19964 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_4_210
timestamp 21601
transform 1 0 20424 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_221
timestamp 21601
transform 1 0 21436 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_230
timestamp 21601
transform 1 0 22264 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_242
timestamp 21601
transform 1 0 23368 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_245
timestamp 21601
transform 1 0 23644 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 21601
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_253
timestamp 21601
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 21601
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_26
timestamp 21601
transform 1 0 3496 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_34
timestamp 21601
transform 1 0 4232 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_41
timestamp 21601
transform 1 0 4876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_51
timestamp 21601
transform 1 0 5796 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 21601
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_57
timestamp 21601
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_80
timestamp 21601
transform 1 0 8464 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_83
timestamp 21601
transform 1 0 8740 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_91
timestamp 21601
transform 1 0 9476 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_100
timestamp 21601
transform 1 0 10304 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_108
timestamp 21601
transform 1 0 11040 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 21601
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_113
timestamp 21601
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_117
timestamp 21601
transform 1 0 11868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_125
timestamp 21601
transform 1 0 12604 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_129
timestamp 21601
transform 1 0 12972 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_136
timestamp 21601
transform 1 0 13616 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_152
timestamp 21601
transform 1 0 15088 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_161
timestamp 21601
transform 1 0 15916 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 21601
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_169
timestamp 21601
transform 1 0 16652 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_193
timestamp 21601
transform 1 0 18860 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_200
timestamp 21601
transform 1 0 19504 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_207
timestamp 21601
transform 1 0 20148 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_5_218
timestamp 21601
transform 1 0 21160 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 21601
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_5_225
timestamp 21601
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_228
timestamp 21601
transform 1 0 22080 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_249
timestamp 21601
transform 1 0 24012 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_254
timestamp 21601
transform 1 0 24472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_3
timestamp 21601
transform 1 0 1380 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_6
timestamp 21601
transform 1 0 1656 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_14
timestamp 21601
transform 1 0 2392 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_23
timestamp 21601
transform 1 0 3220 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 21601
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_29
timestamp 21601
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_39
timestamp 21601
transform 1 0 4692 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_42
timestamp 21601
transform 1 0 4968 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_50
timestamp 21601
transform 1 0 5704 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_59
timestamp 21601
transform 1 0 6532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_69
timestamp 21601
transform 1 0 7452 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_72
timestamp 21601
transform 1 0 7728 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 21601
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_85
timestamp 21601
transform 1 0 8924 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_89
timestamp 21601
transform 1 0 9292 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_96
timestamp 21601
transform 1 0 9936 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_108
timestamp 21601
transform 1 0 11040 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_116
timestamp 21601
transform 1 0 11776 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_120
timestamp 21601
transform 1 0 12144 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_127
timestamp 21601
transform 1 0 12788 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 21601
transform 1 0 13800 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_141
timestamp 21601
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_148
timestamp 21601
transform 1 0 14720 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_154
timestamp 21601
transform 1 0 15272 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_160
timestamp 21601
transform 1 0 15824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_163
timestamp 21601
transform 1 0 16100 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_171
timestamp 21601
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_174
timestamp 21601
transform 1 0 17112 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_185
timestamp 21601
transform 1 0 18124 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 21601
transform 1 0 18952 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_197
timestamp 21601
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_203
timestamp 21601
transform 1 0 19780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_225
timestamp 21601
transform 1 0 21804 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_233
timestamp 21601
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_236
timestamp 21601
transform 1 0 22816 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_247
timestamp 21601
transform 1 0 23828 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 21601
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_253
timestamp 21601
transform 1 0 24380 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_3
timestamp 21601
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_12
timestamp 21601
transform 1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_28
timestamp 21601
transform 1 0 3680 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_31
timestamp 21601
transform 1 0 3956 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_36
timestamp 21601
transform 1 0 4416 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 21601
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_57
timestamp 21601
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_60
timestamp 21601
transform 1 0 6624 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_70
timestamp 21601
transform 1 0 7544 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_85
timestamp 21601
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_94
timestamp 21601
transform 1 0 9752 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_97
timestamp 21601
transform 1 0 10028 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_108
timestamp 21601
transform 1 0 11040 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 21601
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_113
timestamp 21601
transform 1 0 11500 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_120
timestamp 21601
transform 1 0 12144 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_129
timestamp 21601
transform 1 0 12972 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_140
timestamp 21601
transform 1 0 13984 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_147
timestamp 21601
transform 1 0 14628 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_158
timestamp 21601
transform 1 0 15640 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_164
timestamp 21601
transform 1 0 16192 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 21601
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_169
timestamp 21601
transform 1 0 16652 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_7_192
timestamp 21601
transform 1 0 18768 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_7_214
timestamp 21601
transform 1 0 20792 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_221
timestamp 21601
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_225
timestamp 21601
transform 1 0 21804 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_228
timestamp 21601
transform 1 0 22080 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_234
timestamp 21601
transform 1 0 22632 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_245
timestamp 21601
transform 1 0 23644 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_248
timestamp 21601
transform 1 0 23920 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_254
timestamp 21601
transform 1 0 24472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 21601
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_26
timestamp 21601
transform 1 0 3496 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_29
timestamp 21601
transform 1 0 3772 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_37
timestamp 21601
transform 1 0 4508 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_44
timestamp 21601
transform 1 0 5152 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_55
timestamp 21601
transform 1 0 6164 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_60
timestamp 21601
transform 1 0 6624 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_75
timestamp 21601
transform 1 0 8004 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 21601
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_85
timestamp 21601
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_89
timestamp 21601
transform 1 0 9292 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_101
timestamp 21601
transform 1 0 10396 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_109
timestamp 21601
transform 1 0 11132 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_116
timestamp 21601
transform 1 0 11776 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_119
timestamp 21601
transform 1 0 12052 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_129
timestamp 21601
transform 1 0 12972 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_136
timestamp 21601
transform 1 0 13616 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 21601
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_141
timestamp 21601
transform 1 0 14076 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_146
timestamp 21601
transform 1 0 14536 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_154
timestamp 21601
transform 1 0 15272 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_167
timestamp 21601
transform 1 0 16468 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_8_174
timestamp 21601
transform 1 0 17112 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_177
timestamp 21601
transform 1 0 17388 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_184
timestamp 21601
transform 1 0 18032 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_190
timestamp 21601
transform 1 0 18584 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 21601
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_197
timestamp 21601
transform 1 0 19228 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_202
timestamp 21601
transform 1 0 19688 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_224
timestamp 21601
transform 1 0 21712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_8_229
timestamp 21601
transform 1 0 22172 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 21601
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_253
timestamp 21601
transform 1 0 24380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 21601
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_7
timestamp 21601
transform 1 0 1748 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_17
timestamp 21601
transform 1 0 2668 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34
timestamp 21601
transform 1 0 4232 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_37
timestamp 21601
transform 1 0 4508 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_51
timestamp 21601
transform 1 0 5796 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 21601
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 21601
transform 1 0 6348 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_63
timestamp 21601
transform 1 0 6900 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_68
timestamp 21601
transform 1 0 7360 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_74
timestamp 21601
transform 1 0 7912 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_77
timestamp 21601
transform 1 0 8188 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_86
timestamp 21601
transform 1 0 9016 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_97
timestamp 21601
transform 1 0 10028 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_104
timestamp 21601
transform 1 0 10672 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 21601
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_113
timestamp 21601
transform 1 0 11500 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_136
timestamp 21601
transform 1 0 13616 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_145
timestamp 21601
transform 1 0 14444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_156
timestamp 21601
transform 1 0 15456 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_161
timestamp 21601
transform 1 0 15916 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 21601
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_169
timestamp 21601
transform 1 0 16652 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_179
timestamp 21601
transform 1 0 17572 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_185
timestamp 21601
transform 1 0 18124 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_190
timestamp 21601
transform 1 0 18584 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_201
timestamp 21601
transform 1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_204
timestamp 21601
transform 1 0 19872 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_215
timestamp 21601
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 21601
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_225
timestamp 21601
transform 1 0 21804 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_247
timestamp 21601
transform 1 0 23828 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_254
timestamp 21601
transform 1 0 24472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 21601
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_11
timestamp 21601
transform 1 0 2116 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_19
timestamp 21601
transform 1 0 2852 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 21601
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_29
timestamp 21601
transform 1 0 3772 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_40
timestamp 21601
transform 1 0 4784 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_48
timestamp 21601
transform 1 0 5520 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_56
timestamp 21601
transform 1 0 6256 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_64
timestamp 21601
transform 1 0 6992 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_73
timestamp 21601
transform 1 0 7820 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_76
timestamp 21601
transform 1 0 8096 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 21601
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 21601
transform 1 0 8924 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_97
timestamp 21601
transform 1 0 10028 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_102
timestamp 21601
transform 1 0 10488 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_126
timestamp 21601
transform 1 0 12696 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_138
timestamp 21601
transform 1 0 13800 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_141
timestamp 21601
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_162
timestamp 21601
transform 1 0 16008 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_184
timestamp 21601
transform 1 0 18032 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_191
timestamp 21601
transform 1 0 18676 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 21601
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_197
timestamp 21601
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_10_204
timestamp 21601
transform 1 0 19872 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_226
timestamp 21601
transform 1 0 21896 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_237
timestamp 21601
transform 1 0 22908 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_10_248
timestamp 21601
transform 1 0 23920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 21601
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_253
timestamp 21601
transform 1 0 24380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_3
timestamp 21601
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_24
timestamp 21601
transform 1 0 3312 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_31
timestamp 21601
transform 1 0 3956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_38
timestamp 21601
transform 1 0 4600 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_42
timestamp 21601
transform 1 0 4968 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_47
timestamp 21601
transform 1 0 5428 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 21601
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_57
timestamp 21601
transform 1 0 6348 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_62
timestamp 21601
transform 1 0 6808 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_65
timestamp 21601
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_72
timestamp 21601
transform 1 0 7728 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_79
timestamp 21601
transform 1 0 8372 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_84
timestamp 21601
transform 1 0 8832 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_87
timestamp 21601
transform 1 0 9108 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 21601
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_113
timestamp 21601
transform 1 0 11500 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_11_124
timestamp 21601
transform 1 0 12512 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_132
timestamp 21601
transform 1 0 13248 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_139
timestamp 21601
transform 1 0 13892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_11_142
timestamp 21601
transform 1 0 14168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_148
timestamp 21601
transform 1 0 14720 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_155
timestamp 21601
transform 1 0 15364 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_162
timestamp 21601
transform 1 0 16008 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 21601
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_169
timestamp 21601
transform 1 0 16652 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_172
timestamp 21601
transform 1 0 16928 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_194
timestamp 21601
transform 1 0 18952 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_216
timestamp 21601
transform 1 0 20976 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 21601
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_225
timestamp 21601
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_228
timestamp 21601
transform 1 0 22080 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_250
timestamp 21601
transform 1 0 24104 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_254
timestamp 21601
transform 1 0 24472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 21601
transform 1 0 1380 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_7
timestamp 21601
transform 1 0 1748 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_12
timestamp 21601
transform 1 0 2208 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_23
timestamp 21601
transform 1 0 3220 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 21601
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_29
timestamp 21601
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_53
timestamp 21601
transform 1 0 5980 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_56
timestamp 21601
transform 1 0 6256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_62
timestamp 21601
transform 1 0 6808 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_71
timestamp 21601
transform 1 0 7636 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_74
timestamp 21601
transform 1 0 7912 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 21601
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_85
timestamp 21601
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_94
timestamp 21601
transform 1 0 9752 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_100
timestamp 21601
transform 1 0 10304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_112
timestamp 21601
transform 1 0 11408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_122
timestamp 21601
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_125
timestamp 21601
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_128
timestamp 21601
transform 1 0 12880 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_134
timestamp 21601
transform 1 0 13432 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 21601
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 21601
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_162
timestamp 21601
transform 1 0 16008 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_165
timestamp 21601
transform 1 0 16284 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_171
timestamp 21601
transform 1 0 16836 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_177
timestamp 21601
transform 1 0 17388 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_188
timestamp 21601
transform 1 0 18400 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 21601
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 21601
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_207
timestamp 21601
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_210
timestamp 21601
transform 1 0 20424 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_220
timestamp 21601
transform 1 0 21344 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_224
timestamp 21601
transform 1 0 21712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_235
timestamp 21601
transform 1 0 22724 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_12_246
timestamp 21601
transform 1 0 23736 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 21601
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_253
timestamp 21601
transform 1 0 24380 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_3
timestamp 21601
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_6
timestamp 21601
transform 1 0 1656 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_12
timestamp 21601
transform 1 0 2208 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_23
timestamp 21601
transform 1 0 3220 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_28
timestamp 21601
transform 1 0 3680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_32
timestamp 21601
transform 1 0 4048 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_35
timestamp 21601
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_38
timestamp 21601
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_41
timestamp 21601
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_44
timestamp 21601
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_47
timestamp 21601
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 21601
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 21601
transform 1 0 6348 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_67
timestamp 21601
transform 1 0 7268 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_90
timestamp 21601
transform 1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_93
timestamp 21601
transform 1 0 9660 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_97
timestamp 21601
transform 1 0 10028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_107
timestamp 21601
transform 1 0 10948 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_110
timestamp 21601
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_113
timestamp 21601
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_13_124
timestamp 21601
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_133
timestamp 21601
transform 1 0 13340 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 21601
transform 1 0 14168 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_151
timestamp 21601
transform 1 0 14996 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_158
timestamp 21601
transform 1 0 15640 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_164
timestamp 21601
transform 1 0 16192 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 21601
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_169
timestamp 21601
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_192
timestamp 21601
transform 1 0 18768 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_196
timestamp 21601
transform 1 0 19136 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_207
timestamp 21601
transform 1 0 20148 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_214
timestamp 21601
transform 1 0 20792 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_221
timestamp 21601
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_225
timestamp 21601
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_247
timestamp 21601
transform 1 0 23828 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_254
timestamp 21601
transform 1 0 24472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_3
timestamp 21601
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_25
timestamp 21601
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_29
timestamp 21601
transform 1 0 3772 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 21601
transform 1 0 4048 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_35
timestamp 21601
transform 1 0 4324 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_43
timestamp 21601
transform 1 0 5060 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_53
timestamp 21601
transform 1 0 5980 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_61
timestamp 21601
transform 1 0 6716 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_72
timestamp 21601
transform 1 0 7728 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_75
timestamp 21601
transform 1 0 8004 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_82
timestamp 21601
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_85
timestamp 21601
transform 1 0 8924 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_88
timestamp 21601
transform 1 0 9200 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_96
timestamp 21601
transform 1 0 9936 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_104
timestamp 21601
transform 1 0 10672 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_115
timestamp 21601
transform 1 0 11684 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_127
timestamp 21601
transform 1 0 12788 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 21601
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_141
timestamp 21601
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_163
timestamp 21601
transform 1 0 16100 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_185
timestamp 21601
transform 1 0 18124 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_192
timestamp 21601
transform 1 0 18768 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 21601
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_197
timestamp 21601
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_218
timestamp 21601
transform 1 0 21160 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_14_224
timestamp 21601
transform 1 0 21712 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_14_229
timestamp 21601
transform 1 0 22172 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_14_236
timestamp 21601
transform 1 0 22816 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_244
timestamp 21601
transform 1 0 23552 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_247
timestamp 21601
transform 1 0 23828 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 21601
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_253
timestamp 21601
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_3
timestamp 21601
transform 1 0 1380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_6
timestamp 21601
transform 1 0 1656 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_13
timestamp 21601
transform 1 0 2300 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_24
timestamp 21601
transform 1 0 3312 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_27
timestamp 21601
transform 1 0 3588 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_30
timestamp 21601
transform 1 0 3864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_33
timestamp 21601
transform 1 0 4140 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 21601
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_57
timestamp 21601
transform 1 0 6348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_61
timestamp 21601
transform 1 0 6716 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_69
timestamp 21601
transform 1 0 7452 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_72
timestamp 21601
transform 1 0 7728 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_75
timestamp 21601
transform 1 0 8004 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_78
timestamp 21601
transform 1 0 8280 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_81
timestamp 21601
transform 1 0 8556 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_84
timestamp 21601
transform 1 0 8832 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 21601
transform 1 0 9384 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_96
timestamp 21601
transform 1 0 9936 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_15_99
timestamp 21601
transform 1 0 10212 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 21601
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_113
timestamp 21601
transform 1 0 11500 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 21601
transform 1 0 12788 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_136
timestamp 21601
transform 1 0 13616 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_141
timestamp 21601
transform 1 0 14076 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_151
timestamp 21601
transform 1 0 14996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_160
timestamp 21601
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_165
timestamp 21601
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_15_169
timestamp 21601
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_179
timestamp 21601
transform 1 0 17572 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_190
timestamp 21601
transform 1 0 18584 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_15_197
timestamp 21601
transform 1 0 19228 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_15_200
timestamp 21601
transform 1 0 19504 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_222
timestamp 21601
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_225
timestamp 21601
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_231
timestamp 21601
transform 1 0 22356 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_253
timestamp 21601
transform 1 0 24380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_3
timestamp 21601
transform 1 0 1380 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_26
timestamp 21601
transform 1 0 3496 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_29
timestamp 21601
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 21601
transform 1 0 4048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_37
timestamp 21601
transform 1 0 4508 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_44
timestamp 21601
transform 1 0 5152 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_53
timestamp 21601
transform 1 0 5980 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_56
timestamp 21601
transform 1 0 6256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_59
timestamp 21601
transform 1 0 6532 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 21601
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_85
timestamp 21601
transform 1 0 8924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_106
timestamp 21601
transform 1 0 10856 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_109
timestamp 21601
transform 1 0 11132 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_129
timestamp 21601
transform 1 0 12972 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_136
timestamp 21601
transform 1 0 13616 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 21601
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_141
timestamp 21601
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_144
timestamp 21601
transform 1 0 14352 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_152
timestamp 21601
transform 1 0 15088 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_163
timestamp 21601
transform 1 0 16100 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_168
timestamp 21601
transform 1 0 16560 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_171
timestamp 21601
transform 1 0 16836 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_174
timestamp 21601
transform 1 0 17112 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_16_177
timestamp 21601
transform 1 0 17388 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_183
timestamp 21601
transform 1 0 17940 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_16_190
timestamp 21601
transform 1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_193
timestamp 21601
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_197
timestamp 21601
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_200
timestamp 21601
transform 1 0 19504 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_16_203
timestamp 21601
transform 1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_16_206
timestamp 21601
transform 1 0 20056 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_217
timestamp 21601
transform 1 0 21068 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_221
timestamp 21601
transform 1 0 21436 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_243
timestamp 21601
transform 1 0 23460 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 21601
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_253
timestamp 21601
transform 1 0 24380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_3
timestamp 21601
transform 1 0 1380 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_26
timestamp 21601
transform 1 0 3496 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_29
timestamp 21601
transform 1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 21601
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_57
timestamp 21601
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_64
timestamp 21601
transform 1 0 6992 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_67
timestamp 21601
transform 1 0 7268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_75
timestamp 21601
transform 1 0 8004 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_81
timestamp 21601
transform 1 0 8556 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_84
timestamp 21601
transform 1 0 8832 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_97
timestamp 21601
transform 1 0 10028 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_100
timestamp 21601
transform 1 0 10304 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 21601
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_113
timestamp 21601
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_125
timestamp 21601
transform 1 0 12604 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_130
timestamp 21601
transform 1 0 13064 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_148
timestamp 21601
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_159
timestamp 21601
transform 1 0 15732 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 21601
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_169
timestamp 21601
transform 1 0 16652 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_172
timestamp 21601
transform 1 0 16928 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_193
timestamp 21601
transform 1 0 18860 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_196
timestamp 21601
transform 1 0 19136 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_199
timestamp 21601
transform 1 0 19412 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_202
timestamp 21601
transform 1 0 19688 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_17_205
timestamp 21601
transform 1 0 19964 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_208
timestamp 21601
transform 1 0 20240 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_216
timestamp 21601
transform 1 0 20976 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_17_219
timestamp 21601
transform 1 0 21252 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 21601
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 21601
transform 1 0 21804 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_17_235
timestamp 21601
transform 1 0 22724 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_17_247
timestamp 21601
transform 1 0 23828 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_17_252
timestamp 21601
transform 1 0 24288 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_3
timestamp 21601
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_6
timestamp 21601
transform 1 0 1656 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_13
timestamp 21601
transform 1 0 2300 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_24
timestamp 21601
transform 1 0 3312 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 21601
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_29
timestamp 21601
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_32
timestamp 21601
transform 1 0 4048 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_39
timestamp 21601
transform 1 0 4692 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_61
timestamp 21601
transform 1 0 6716 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_64
timestamp 21601
transform 1 0 6992 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_67
timestamp 21601
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_77
timestamp 21601
transform 1 0 8188 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 21601
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_85
timestamp 21601
transform 1 0 8924 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 21601
transform 1 0 9384 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_100
timestamp 21601
transform 1 0 10304 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_119
timestamp 21601
transform 1 0 12052 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_130
timestamp 21601
transform 1 0 13064 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_137
timestamp 21601
transform 1 0 13708 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_141
timestamp 21601
transform 1 0 14076 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_144
timestamp 21601
transform 1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_18_147
timestamp 21601
transform 1 0 14628 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_150
timestamp 21601
transform 1 0 14904 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_156
timestamp 21601
transform 1 0 15456 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_164
timestamp 21601
transform 1 0 16192 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_167
timestamp 21601
transform 1 0 16468 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_192
timestamp 21601
transform 1 0 18768 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 21601
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_18_197
timestamp 21601
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_18_200
timestamp 21601
transform 1 0 19504 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_208
timestamp 21601
transform 1 0 20240 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_18_218
timestamp 21601
transform 1 0 21160 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_18_221
timestamp 21601
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_231
timestamp 21601
transform 1 0 22356 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_236
timestamp 21601
transform 1 0 22816 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_245
timestamp 21601
transform 1 0 23644 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 21601
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_253
timestamp 21601
transform 1 0 24380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_3
timestamp 21601
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_7
timestamp 21601
transform 1 0 1748 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_11
timestamp 21601
transform 1 0 2116 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_33
timestamp 21601
transform 1 0 4140 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_36
timestamp 21601
transform 1 0 4416 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_39
timestamp 21601
transform 1 0 4692 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_44
timestamp 21601
transform 1 0 5152 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 21601
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_19_57
timestamp 21601
transform 1 0 6348 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_63
timestamp 21601
transform 1 0 6900 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_85
timestamp 21601
transform 1 0 8924 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_88
timestamp 21601
transform 1 0 9200 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_98
timestamp 21601
transform 1 0 10120 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_109
timestamp 21601
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_113
timestamp 21601
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 21601
transform 1 0 12420 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_126
timestamp 21601
transform 1 0 12696 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_129
timestamp 21601
transform 1 0 12972 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_139
timestamp 21601
transform 1 0 13892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_142
timestamp 21601
transform 1 0 14168 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_150
timestamp 21601
transform 1 0 14904 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_158
timestamp 21601
transform 1 0 15640 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_163
timestamp 21601
transform 1 0 16100 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_166
timestamp 21601
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_19_169
timestamp 21601
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_172
timestamp 21601
transform 1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_19_195
timestamp 21601
transform 1 0 19044 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_198
timestamp 21601
transform 1 0 19320 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_203
timestamp 21601
transform 1 0 19780 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_213
timestamp 21601
transform 1 0 20700 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_222
timestamp 21601
transform 1 0 21528 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_225
timestamp 21601
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_233
timestamp 21601
transform 1 0 22540 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_19_236
timestamp 21601
transform 1 0 22816 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_248
timestamp 21601
transform 1 0 23920 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_254
timestamp 21601
transform 1 0 24472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_3
timestamp 21601
transform 1 0 1380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_24
timestamp 21601
transform 1 0 3312 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 21601
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_29
timestamp 21601
transform 1 0 3772 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_39
timestamp 21601
transform 1 0 4692 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_61
timestamp 21601
transform 1 0 6716 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_72
timestamp 21601
transform 1 0 7728 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_80
timestamp 21601
transform 1 0 8464 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 21601
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 21601
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_88
timestamp 21601
transform 1 0 9200 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_98
timestamp 21601
transform 1 0 10120 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_104
timestamp 21601
transform 1 0 10672 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_119
timestamp 21601
transform 1 0 12052 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_128
timestamp 21601
transform 1 0 12880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_138
timestamp 21601
transform 1 0 13800 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_141
timestamp 21601
transform 1 0 14076 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_144
timestamp 21601
transform 1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_147
timestamp 21601
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_156
timestamp 21601
transform 1 0 15456 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_162
timestamp 21601
transform 1 0 16008 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_20_167
timestamp 21601
transform 1 0 16468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_170
timestamp 21601
transform 1 0 16744 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_177
timestamp 21601
transform 1 0 17388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_184
timestamp 21601
transform 1 0 18032 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 21601
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_20_197
timestamp 21601
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_209
timestamp 21601
transform 1 0 20332 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_20_212
timestamp 21601
transform 1 0 20608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_20_222
timestamp 21601
transform 1 0 21528 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_230
timestamp 21601
transform 1 0 22264 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_250
timestamp 21601
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_253
timestamp 21601
transform 1 0 24380 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_3
timestamp 21601
transform 1 0 1380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_7
timestamp 21601
transform 1 0 1748 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_15
timestamp 21601
transform 1 0 2484 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_26
timestamp 21601
transform 1 0 3496 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_33
timestamp 21601
transform 1 0 4140 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_36
timestamp 21601
transform 1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_39
timestamp 21601
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_42
timestamp 21601
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_45
timestamp 21601
transform 1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_48
timestamp 21601
transform 1 0 5520 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 21601
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_57
timestamp 21601
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_60
timestamp 21601
transform 1 0 6624 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_63
timestamp 21601
transform 1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_66
timestamp 21601
transform 1 0 7176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_69
timestamp 21601
transform 1 0 7452 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_75
timestamp 21601
transform 1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_100
timestamp 21601
transform 1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_109
timestamp 21601
transform 1 0 11132 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_113
timestamp 21601
transform 1 0 11500 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_120
timestamp 21601
transform 1 0 12144 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_123
timestamp 21601
transform 1 0 12420 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_132
timestamp 21601
transform 1 0 13248 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_135
timestamp 21601
transform 1 0 13524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_145
timestamp 21601
transform 1 0 14444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_153
timestamp 21601
transform 1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_160
timestamp 21601
transform 1 0 15824 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 21601
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_169
timestamp 21601
transform 1 0 16652 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_190
timestamp 21601
transform 1 0 18584 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_21_211
timestamp 21601
transform 1 0 20516 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_220
timestamp 21601
transform 1 0 21344 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 21601
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_21_225
timestamp 21601
transform 1 0 21804 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_237
timestamp 21601
transform 1 0 22908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_246
timestamp 21601
transform 1 0 23736 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_254
timestamp 21601
transform 1 0 24472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_3
timestamp 21601
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_6
timestamp 21601
transform 1 0 1656 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_13
timestamp 21601
transform 1 0 2300 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_24
timestamp 21601
transform 1 0 3312 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 21601
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_29
timestamp 21601
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_32
timestamp 21601
transform 1 0 4048 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_35
timestamp 21601
transform 1 0 4324 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_38
timestamp 21601
transform 1 0 4600 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_41
timestamp 21601
transform 1 0 4876 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_44
timestamp 21601
transform 1 0 5152 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_56
timestamp 21601
transform 1 0 6256 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_59
timestamp 21601
transform 1 0 6532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_62
timestamp 21601
transform 1 0 6808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_65
timestamp 21601
transform 1 0 7084 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_68
timestamp 21601
transform 1 0 7360 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_71
timestamp 21601
transform 1 0 7636 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_82
timestamp 21601
transform 1 0 8648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_85
timestamp 21601
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_92
timestamp 21601
transform 1 0 9568 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_106
timestamp 21601
transform 1 0 10856 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_111
timestamp 21601
transform 1 0 11316 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_118
timestamp 21601
transform 1 0 11960 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_128
timestamp 21601
transform 1 0 12880 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 21601
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_22_141
timestamp 21601
transform 1 0 14076 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_144
timestamp 21601
transform 1 0 14352 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_147
timestamp 21601
transform 1 0 14628 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_158
timestamp 21601
transform 1 0 15640 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_166
timestamp 21601
transform 1 0 16376 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_173
timestamp 21601
transform 1 0 17020 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_176
timestamp 21601
transform 1 0 17296 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_179
timestamp 21601
transform 1 0 17572 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_22_185
timestamp 21601
transform 1 0 18124 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_194
timestamp 21601
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_22_197
timestamp 21601
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_22_207
timestamp 21601
transform 1 0 20148 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_22_210
timestamp 21601
transform 1 0 20424 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_218
timestamp 21601
transform 1 0 21160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_238
timestamp 21601
transform 1 0 23000 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_247
timestamp 21601
transform 1 0 23828 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 21601
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_22_253
timestamp 21601
transform 1 0 24380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_3
timestamp 21601
transform 1 0 1380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_25
timestamp 21601
transform 1 0 3404 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_32
timestamp 21601
transform 1 0 4048 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 21601
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_57
timestamp 21601
transform 1 0 6348 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_63
timestamp 21601
transform 1 0 6900 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_85
timestamp 21601
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_92
timestamp 21601
transform 1 0 9568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_100
timestamp 21601
transform 1 0 10304 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 21601
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_23_113
timestamp 21601
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_119
timestamp 21601
transform 1 0 12052 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_124
timestamp 21601
transform 1 0 12512 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_127
timestamp 21601
transform 1 0 12788 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_144
timestamp 21601
transform 1 0 14352 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_23_147
timestamp 21601
transform 1 0 14628 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_156
timestamp 21601
transform 1 0 15456 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_163
timestamp 21601
transform 1 0 16100 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_166
timestamp 21601
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_169
timestamp 21601
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_176
timestamp 21601
transform 1 0 17296 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_180
timestamp 21601
transform 1 0 17664 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_200
timestamp 21601
transform 1 0 19504 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_208
timestamp 21601
transform 1 0 20240 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_214
timestamp 21601
transform 1 0 20792 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_218
timestamp 21601
transform 1 0 21160 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 21601
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_225
timestamp 21601
transform 1 0 21804 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_231
timestamp 21601
transform 1 0 22356 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_244
timestamp 21601
transform 1 0 23552 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_253
timestamp 21601
transform 1 0 24380 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_24_3
timestamp 21601
transform 1 0 1380 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_24
timestamp 21601
transform 1 0 3312 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 21601
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_29
timestamp 21601
transform 1 0 3772 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_39
timestamp 21601
transform 1 0 4692 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_62
timestamp 21601
transform 1 0 6808 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_65
timestamp 21601
transform 1 0 7084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_71
timestamp 21601
transform 1 0 7636 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_82
timestamp 21601
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_85
timestamp 21601
transform 1 0 8924 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_92
timestamp 21601
transform 1 0 9568 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_102
timestamp 21601
transform 1 0 10488 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_113
timestamp 21601
transform 1 0 11500 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_122
timestamp 21601
transform 1 0 12328 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_127
timestamp 21601
transform 1 0 12788 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_135
timestamp 21601
transform 1 0 13524 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_138
timestamp 21601
transform 1 0 13800 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_141
timestamp 21601
transform 1 0 14076 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_144
timestamp 21601
transform 1 0 14352 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_156
timestamp 21601
transform 1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_24_159
timestamp 21601
transform 1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_170
timestamp 21601
transform 1 0 16744 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_177
timestamp 21601
transform 1 0 17388 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_180
timestamp 21601
transform 1 0 17664 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_193
timestamp 21601
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_197
timestamp 21601
transform 1 0 19228 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_205
timestamp 21601
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_210
timestamp 21601
transform 1 0 20424 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_24_213
timestamp 21601
transform 1 0 20700 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_218
timestamp 21601
transform 1 0 21160 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_223
timestamp 21601
transform 1 0 21620 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_228
timestamp 21601
transform 1 0 22080 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_24_248
timestamp 21601
transform 1 0 23920 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 21601
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_24_253
timestamp 21601
transform 1 0 24380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_3
timestamp 21601
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_7
timestamp 21601
transform 1 0 1748 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_10
timestamp 21601
transform 1 0 2024 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_16
timestamp 21601
transform 1 0 2576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_19
timestamp 21601
transform 1 0 2852 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_40
timestamp 21601
transform 1 0 4784 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_43
timestamp 21601
transform 1 0 5060 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_46
timestamp 21601
transform 1 0 5336 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_54
timestamp 21601
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_57
timestamp 21601
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_60
timestamp 21601
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_63
timestamp 21601
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_85
timestamp 21601
transform 1 0 8924 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_25_88
timestamp 21601
transform 1 0 9200 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_99
timestamp 21601
transform 1 0 10212 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_110
timestamp 21601
transform 1 0 11224 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_113
timestamp 21601
transform 1 0 11500 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_120
timestamp 21601
transform 1 0 12144 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_123
timestamp 21601
transform 1 0 12420 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_132
timestamp 21601
transform 1 0 13248 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_143
timestamp 21601
transform 1 0 14260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_150
timestamp 21601
transform 1 0 14904 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_160
timestamp 21601
transform 1 0 15824 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 21601
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 21601
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_177
timestamp 21601
transform 1 0 17388 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_180
timestamp 21601
transform 1 0 17664 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_184
timestamp 21601
transform 1 0 18032 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_197
timestamp 21601
transform 1 0 19228 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_202
timestamp 21601
transform 1 0 19688 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_25_205
timestamp 21601
transform 1 0 19964 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_214
timestamp 21601
transform 1 0 20792 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 21601
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_225
timestamp 21601
transform 1 0 21804 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_234
timestamp 21601
transform 1 0 22632 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_243
timestamp 21601
transform 1 0 23460 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_249
timestamp 21601
transform 1 0 24012 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 21601
transform 1 0 24472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_3
timestamp 21601
transform 1 0 1380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_6
timestamp 21601
transform 1 0 1656 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_9
timestamp 21601
transform 1 0 1932 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_21
timestamp 21601
transform 1 0 3036 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_24
timestamp 21601
transform 1 0 3312 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 21601
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_29
timestamp 21601
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_32
timestamp 21601
transform 1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_44
timestamp 21601
transform 1 0 5152 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_51
timestamp 21601
transform 1 0 5796 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_62
timestamp 21601
transform 1 0 6808 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_65
timestamp 21601
transform 1 0 7084 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_68
timestamp 21601
transform 1 0 7360 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_71
timestamp 21601
transform 1 0 7636 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 21601
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 21601
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_88
timestamp 21601
transform 1 0 9200 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_91
timestamp 21601
transform 1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_94
timestamp 21601
transform 1 0 9752 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_97
timestamp 21601
transform 1 0 10028 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_108
timestamp 21601
transform 1 0 11040 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_111
timestamp 21601
transform 1 0 11316 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_121
timestamp 21601
transform 1 0 12236 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_124
timestamp 21601
transform 1 0 12512 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_131
timestamp 21601
transform 1 0 13156 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_134
timestamp 21601
transform 1 0 13432 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_137
timestamp 21601
transform 1 0 13708 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_141
timestamp 21601
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_144
timestamp 21601
transform 1 0 14352 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_152
timestamp 21601
transform 1 0 15088 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_162
timestamp 21601
transform 1 0 16008 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_26_171
timestamp 21601
transform 1 0 16836 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_174
timestamp 21601
transform 1 0 17112 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_194
timestamp 21601
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_197
timestamp 21601
transform 1 0 19228 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_201
timestamp 21601
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_26_212
timestamp 21601
transform 1 0 20608 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_215
timestamp 21601
transform 1 0 20884 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_230
timestamp 21601
transform 1 0 22264 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_26_233
timestamp 21601
transform 1 0 22540 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_246
timestamp 21601
transform 1 0 23736 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 21601
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_253
timestamp 21601
transform 1 0 24380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_3
timestamp 21601
transform 1 0 1380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_7
timestamp 21601
transform 1 0 1748 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_11
timestamp 21601
transform 1 0 2116 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_22
timestamp 21601
transform 1 0 3128 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_25
timestamp 21601
transform 1 0 3404 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_28
timestamp 21601
transform 1 0 3680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_50
timestamp 21601
transform 1 0 5704 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_53
timestamp 21601
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_57
timestamp 21601
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_60
timestamp 21601
transform 1 0 6624 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_63
timestamp 21601
transform 1 0 6900 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_86
timestamp 21601
transform 1 0 9016 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_89
timestamp 21601
transform 1 0 9292 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_92
timestamp 21601
transform 1 0 9568 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_95
timestamp 21601
transform 1 0 9844 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_98
timestamp 21601
transform 1 0 10120 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_106
timestamp 21601
transform 1 0 10856 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 21601
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_113
timestamp 21601
transform 1 0 11500 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_27_132
timestamp 21601
transform 1 0 13248 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_143
timestamp 21601
transform 1 0 14260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_147
timestamp 21601
transform 1 0 14628 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_150
timestamp 21601
transform 1 0 14904 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_153
timestamp 21601
transform 1 0 15180 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_162
timestamp 21601
transform 1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_27_165
timestamp 21601
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 21601
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_176
timestamp 21601
transform 1 0 17296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 21601
transform 1 0 17756 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_190
timestamp 21601
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_199
timestamp 21601
transform 1 0 19412 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_208
timestamp 21601
transform 1 0 20240 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_213
timestamp 21601
transform 1 0 20700 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 21601
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_225
timestamp 21601
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_27_228
timestamp 21601
transform 1 0 22080 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_240
timestamp 21601
transform 1 0 23184 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_249
timestamp 21601
transform 1 0 24012 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_254
timestamp 21601
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_3
timestamp 21601
transform 1 0 1380 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_24
timestamp 21601
transform 1 0 3312 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 21601
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_29
timestamp 21601
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_37
timestamp 21601
transform 1 0 4508 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_48
timestamp 21601
transform 1 0 5520 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_55
timestamp 21601
transform 1 0 6164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_63
timestamp 21601
transform 1 0 6900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_74
timestamp 21601
transform 1 0 7912 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_81
timestamp 21601
transform 1 0 8556 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_85
timestamp 21601
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_88
timestamp 21601
transform 1 0 9200 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_91
timestamp 21601
transform 1 0 9476 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_94
timestamp 21601
transform 1 0 9752 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_98
timestamp 21601
transform 1 0 10120 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_107
timestamp 21601
transform 1 0 10948 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_120
timestamp 21601
transform 1 0 12144 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_126
timestamp 21601
transform 1 0 12696 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_129
timestamp 21601
transform 1 0 12972 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 21601
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 21601
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_145
timestamp 21601
transform 1 0 14444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_150
timestamp 21601
transform 1 0 14904 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_160
timestamp 21601
transform 1 0 15824 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_28_169
timestamp 21601
transform 1 0 16652 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_28_172
timestamp 21601
transform 1 0 16928 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_178
timestamp 21601
transform 1 0 17480 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 21601
transform 1 0 18676 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 21601
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 21601
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_28_202
timestamp 21601
transform 1 0 19688 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_28_205
timestamp 21601
transform 1 0 19964 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_213
timestamp 21601
transform 1 0 20700 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_222
timestamp 21601
transform 1 0 21528 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_230
timestamp 21601
transform 1 0 22264 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 21601
transform 1 0 24104 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_253
timestamp 21601
transform 1 0 24380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 21601
transform 1 0 1380 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_6
timestamp 21601
transform 1 0 1656 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_13
timestamp 21601
transform 1 0 2300 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_24
timestamp 21601
transform 1 0 3312 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_27
timestamp 21601
transform 1 0 3588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_30
timestamp 21601
transform 1 0 3864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_51
timestamp 21601
transform 1 0 5796 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 21601
transform 1 0 6072 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_57
timestamp 21601
transform 1 0 6348 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_78
timestamp 21601
transform 1 0 8280 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_89
timestamp 21601
transform 1 0 9292 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_29_92
timestamp 21601
transform 1 0 9568 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_95
timestamp 21601
transform 1 0 9844 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_102
timestamp 21601
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 21601
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_113
timestamp 21601
transform 1 0 11500 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_125
timestamp 21601
transform 1 0 12604 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_145
timestamp 21601
transform 1 0 14444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_158
timestamp 21601
transform 1 0 15640 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 21601
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_169
timestamp 21601
transform 1 0 16652 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_172
timestamp 21601
transform 1 0 16928 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_192
timestamp 21601
transform 1 0 18768 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_201
timestamp 21601
transform 1 0 19596 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_207
timestamp 21601
transform 1 0 20148 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_212
timestamp 21601
transform 1 0 20608 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_29_215
timestamp 21601
transform 1 0 20884 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 21601
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_225
timestamp 21601
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_29_235
timestamp 21601
transform 1 0 22724 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_250
timestamp 21601
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_254
timestamp 21601
transform 1 0 24472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_3
timestamp 21601
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_30_25
timestamp 21601
transform 1 0 3404 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_29
timestamp 21601
transform 1 0 3772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_32
timestamp 21601
transform 1 0 4048 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_55
timestamp 21601
transform 1 0 6164 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_30_58
timestamp 21601
transform 1 0 6440 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_61
timestamp 21601
transform 1 0 6716 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 21601
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_85
timestamp 21601
transform 1 0 8924 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_30_108
timestamp 21601
transform 1 0 11040 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_128
timestamp 21601
transform 1 0 12880 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_134
timestamp 21601
transform 1 0 13432 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 21601
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 21601
transform 1 0 14076 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_30_144
timestamp 21601
transform 1 0 14352 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 21601
transform 1 0 16100 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_176
timestamp 21601
transform 1 0 17296 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_180
timestamp 21601
transform 1 0 17664 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 21601
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_197
timestamp 21601
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_218
timestamp 21601
transform 1 0 21160 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_224
timestamp 21601
transform 1 0 21712 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_244
timestamp 21601
transform 1 0 23552 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 21601
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_253
timestamp 21601
transform 1 0 24380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_3
timestamp 21601
transform 1 0 1380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_7
timestamp 21601
transform 1 0 1748 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_11
timestamp 21601
transform 1 0 2116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_18
timestamp 21601
transform 1 0 2760 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_23
timestamp 21601
transform 1 0 3220 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_27
timestamp 21601
transform 1 0 3588 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_29
timestamp 21601
transform 1 0 3772 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_34
timestamp 21601
transform 1 0 4232 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_38
timestamp 21601
transform 1 0 4600 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_50
timestamp 21601
transform 1 0 5704 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 21601
transform 1 0 5980 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_57
timestamp 21601
transform 1 0 6348 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 21601
transform 1 0 6808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_66
timestamp 21601
transform 1 0 7176 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp 21601
transform 1 0 7452 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_72
timestamp 21601
transform 1 0 7728 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_75
timestamp 21601
transform 1 0 8004 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_31_81
timestamp 21601
transform 1 0 8556 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_85
timestamp 21601
transform 1 0 8924 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_90
timestamp 21601
transform 1 0 9384 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_94
timestamp 21601
transform 1 0 9752 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_97
timestamp 21601
transform 1 0 10028 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_100
timestamp 21601
transform 1 0 10304 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_103
timestamp 21601
transform 1 0 10580 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_106
timestamp 21601
transform 1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 21601
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_113
timestamp 21601
transform 1 0 11500 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp 21601
transform 1 0 12236 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_126
timestamp 21601
transform 1 0 12696 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_129
timestamp 21601
transform 1 0 12972 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_134
timestamp 21601
transform 1 0 13432 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_139
timestamp 21601
transform 1 0 13892 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_141
timestamp 21601
transform 1 0 14076 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_147
timestamp 21601
transform 1 0 14628 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_156
timestamp 21601
transform 1 0 15456 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_165
timestamp 21601
transform 1 0 16284 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 21601
transform 1 0 16652 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_173
timestamp 21601
transform 1 0 17020 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_178
timestamp 21601
transform 1 0 17480 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_181
timestamp 21601
transform 1 0 17756 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_189
timestamp 21601
transform 1 0 18492 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_195
timestamp 21601
transform 1 0 19044 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_197
timestamp 21601
transform 1 0 19228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_201
timestamp 21601
transform 1 0 19596 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_206
timestamp 21601
transform 1 0 20056 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 21601
transform 1 0 20332 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_216
timestamp 21601
transform 1 0 20976 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 21601
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 21601
transform 1 0 21804 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_233
timestamp 21601
transform 1 0 22540 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_238
timestamp 21601
transform 1 0 23000 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_31_244
timestamp 21601
transform 1 0 23552 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_247
timestamp 21601
transform 1 0 23828 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_251
timestamp 21601
transform 1 0 24196 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_253
timestamp 21601
transform 1 0 24380 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__buf_12  input1
timestamp 21601
transform 1 0 20424 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 21601
transform 1 0 1656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 21601
transform -1 0 3680 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 21601
transform -1 0 4692 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 21601
transform -1 0 4784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 21601
transform -1 0 8372 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 21601
transform -1 0 11868 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 21601
transform 1 0 14168 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 21601
transform -1 0 18124 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 21601
transform -1 0 21712 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 21601
transform 1 0 6440 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 21601
transform -1 0 4232 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 21601
transform -1 0 6808 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 21601
transform -1 0 9384 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 21601
transform 1 0 19320 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 21601
transform 1 0 19780 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 21601
transform -1 0 21160 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 21601
transform -1 0 13892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 21601
transform -1 0 13432 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 21601
transform -1 0 18032 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 21601
transform 1 0 23920 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 21601
transform -1 0 1748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 21601
transform 1 0 24196 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 21601
transform 1 0 23920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 21601
transform 1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 21601
transform -1 0 21620 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input27
timestamp 21601
transform -1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 21601
transform 1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 21601
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input30
timestamp 21601
transform 1 0 1472 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input31
timestamp 21601
transform 1 0 1472 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 21601
transform 1 0 1472 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 21601
transform 1 0 1472 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 21601
transform 1 0 1472 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 21601
transform 1 0 2944 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 21601
transform 1 0 1472 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 21601
transform 1 0 24196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 21601
transform -1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_32
timestamp 21601
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 21601
transform -1 0 24840 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_33
timestamp 21601
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 21601
transform -1 0 24840 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_34
timestamp 21601
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 21601
transform -1 0 24840 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_35
timestamp 21601
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 21601
transform -1 0 24840 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_36
timestamp 21601
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 21601
transform -1 0 24840 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_37
timestamp 21601
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 21601
transform -1 0 24840 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_38
timestamp 21601
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 21601
transform -1 0 24840 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_39
timestamp 21601
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 21601
transform -1 0 24840 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_40
timestamp 21601
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 21601
transform -1 0 24840 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_41
timestamp 21601
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 21601
transform -1 0 24840 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_42
timestamp 21601
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 21601
transform -1 0 24840 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_43
timestamp 21601
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 21601
transform -1 0 24840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_44
timestamp 21601
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 21601
transform -1 0 24840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_45
timestamp 21601
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 21601
transform -1 0 24840 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_46
timestamp 21601
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 21601
transform -1 0 24840 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_47
timestamp 21601
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 21601
transform -1 0 24840 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_48
timestamp 21601
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 21601
transform -1 0 24840 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_49
timestamp 21601
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 21601
transform -1 0 24840 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_50
timestamp 21601
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 21601
transform -1 0 24840 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_51
timestamp 21601
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 21601
transform -1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_52
timestamp 21601
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 21601
transform -1 0 24840 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_53
timestamp 21601
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 21601
transform -1 0 24840 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_54
timestamp 21601
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 21601
transform -1 0 24840 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_55
timestamp 21601
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 21601
transform -1 0 24840 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_56
timestamp 21601
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 21601
transform -1 0 24840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_57
timestamp 21601
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 21601
transform -1 0 24840 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_58
timestamp 21601
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 21601
transform -1 0 24840 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_59
timestamp 21601
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 21601
transform -1 0 24840 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_60
timestamp 21601
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 21601
transform -1 0 24840 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_61
timestamp 21601
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 21601
transform -1 0 24840 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_62
timestamp 21601
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 21601
transform -1 0 24840 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Left_63
timestamp 21601
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_31_Right_31
timestamp 21601
transform -1 0 24840 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer1
timestamp 21601
transform 1 0 10488 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer2
timestamp 21601
transform 1 0 13800 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  rebuffer3
timestamp 21601
transform 1 0 9016 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  rebuffer4
timestamp 21601
transform -1 0 22264 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer5
timestamp 21601
transform 1 0 11868 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer7
timestamp 21601
transform -1 0 14168 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer8
timestamp 21601
transform -1 0 15456 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer9
timestamp 21601
transform -1 0 15640 0 1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer10
timestamp 21601
transform -1 0 10120 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer11
timestamp 21601
transform 1 0 11592 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer12
timestamp 21601
transform 1 0 10672 0 -1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer13
timestamp 21601
transform 1 0 12880 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer14
timestamp 21601
transform -1 0 9292 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  rebuffer15
timestamp 21601
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer16
timestamp 21601
transform -1 0 4232 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer17
timestamp 21601
transform 1 0 3864 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer19
timestamp 21601
transform 1 0 17204 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer20
timestamp 21601
transform -1 0 18952 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer21
timestamp 21601
transform -1 0 16836 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer22
timestamp 21601
transform -1 0 14536 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer23
timestamp 21601
transform -1 0 8740 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer24
timestamp 21601
transform -1 0 9752 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer25
timestamp 21601
transform 1 0 16744 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  rebuffer26
timestamp 21601
transform 1 0 10856 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer27
timestamp 21601
transform 1 0 12972 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  rebuffer28
timestamp 21601
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  rebuffer29
timestamp 21601
transform 1 0 10856 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  rebuffer32
timestamp 21601
transform 1 0 12236 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  rebuffer33
timestamp 21601
transform 1 0 8372 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlygate4sd1_1  rebuffer35
timestamp 21601
transform 1 0 19320 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer36
timestamp 21601
transform 1 0 11776 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  rebuffer37
timestamp 21601
transform -1 0 13892 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  rebuffer38
timestamp 21601
transform -1 0 12604 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  rebuffer39
timestamp 21601
transform 1 0 5152 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s4s_1  rebuffer40
timestamp 21601
transform 1 0 9476 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  rebuffer41
timestamp 21601
transform -1 0 15732 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 21601
transform -1 0 21712 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 21601
transform 1 0 17204 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp 21601
transform 1 0 14812 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 21601
transform 1 0 15640 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0
timestamp 21601
transform 1 0 14444 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1
timestamp 21601
transform 1 0 16284 0 1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 21601
transform -1 0 17020 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 21601
transform -1 0 14628 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 21601
transform -1 0 14904 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 21601
transform 1 0 13064 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 21601
transform -1 0 16468 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 21601
transform 1 0 12788 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 21601
transform -1 0 15640 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 21601
transform -1 0 14444 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 21601
transform -1 0 13432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 21601
transform 1 0 12420 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 21601
transform 1 0 10672 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 21601
transform 1 0 11592 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 21601
transform 1 0 11224 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 21601
transform 1 0 11592 0 -1 17408
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 21601
transform -1 0 11316 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 21601
transform 1 0 12328 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 21601
transform -1 0 10120 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 21601
transform 1 0 11592 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 21601
transform -1 0 10948 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 21601
transform 1 0 11592 0 -1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 21601
transform -1 0 12144 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 21601
transform 1 0 11040 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 21601
transform 1 0 12788 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 21601
transform 1 0 19320 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 21601
transform 1 0 17940 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 21601
transform -1 0 19412 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 21601
transform 1 0 17296 0 1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 21601
transform -1 0 19228 0 -1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 21601
transform -1 0 17756 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 21601
transform -1 0 19688 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 21601
transform -1 0 17480 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 21601
transform 1 0 18952 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 21601
transform -1 0 18492 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 21601
transform 1 0 17112 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 21601
transform 1 0 17664 0 1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 21601
transform 1 0 20332 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 21601
transform -1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 21601
transform 1 0 19412 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 21601
transform 1 0 18308 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 21601
transform -1 0 19964 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 21601
transform 1 0 17848 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 21601
transform 1 0 17848 0 1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 21601
transform -1 0 18124 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 21601
transform -1 0 20792 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 21601
transform 1 0 20148 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 21601
transform 1 0 20700 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 21601
transform 1 0 19504 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 21601
transform 1 0 18860 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 21601
transform 1 0 19320 0 1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 21601
transform -1 0 19780 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 21601
transform -1 0 24472 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 21601
transform 1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 21601
transform 1 0 23184 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 21601
transform 1 0 23000 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 21601
transform 1 0 22448 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 21601
transform 1 0 22908 0 -1 11968
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 21601
transform -1 0 21620 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 21601
transform -1 0 24196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 21601
transform -1 0 22816 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 21601
transform 1 0 20516 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 21601
transform -1 0 23736 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 21601
transform 1 0 21344 0 1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 21601
transform 1 0 21896 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 21601
transform -1 0 21620 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 21601
transform -1 0 22356 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 21601
transform -1 0 22080 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 21601
transform 1 0 22816 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 21601
transform -1 0 24380 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 21601
transform 1 0 22264 0 1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 21601
transform -1 0 23552 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 21601
transform 1 0 23920 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 21601
transform -1 0 24012 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 21601
transform -1 0 20700 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 21601
transform 1 0 22080 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 21601
transform -1 0 24012 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 21601
transform 1 0 22448 0 1 16320
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 21601
transform 1 0 22724 0 1 15232
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 21601
transform -1 0 23552 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 21601
transform 1 0 23736 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 21601
transform -1 0 24104 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 21601
transform -1 0 19044 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 21601
transform -1 0 19044 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1562557784
transform 1 0 22724 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 21601
transform 1 0 21160 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 21601
transform -1 0 21620 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 21601
transform 1 0 21896 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 21601
transform -1 0 21620 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 21601
transform 1 0 21896 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 21601
transform 1 0 22172 0 -1 16320
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 21601
transform -1 0 13892 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0
timestamp 21601
transform 1 0 20516 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 21601
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 21601
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 21601
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 21601
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_68
timestamp 21601
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_69
timestamp 21601
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_70
timestamp 21601
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_71
timestamp 21601
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_72
timestamp 21601
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_73
timestamp 21601
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_74
timestamp 21601
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_75
timestamp 21601
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_76
timestamp 21601
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_77
timestamp 21601
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_78
timestamp 21601
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_79
timestamp 21601
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_80
timestamp 21601
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_81
timestamp 21601
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_82
timestamp 21601
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_83
timestamp 21601
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_84
timestamp 21601
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_85
timestamp 21601
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_86
timestamp 21601
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_87
timestamp 21601
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_88
timestamp 21601
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_89
timestamp 21601
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_90
timestamp 21601
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_91
timestamp 21601
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_92
timestamp 21601
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_93
timestamp 21601
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_94
timestamp 21601
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_95
timestamp 21601
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_96
timestamp 21601
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_97
timestamp 21601
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_98
timestamp 21601
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_99
timestamp 21601
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_100
timestamp 21601
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_101
timestamp 21601
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_102
timestamp 21601
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_103
timestamp 21601
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_104
timestamp 21601
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_105
timestamp 21601
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_106
timestamp 21601
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_107
timestamp 21601
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_108
timestamp 21601
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_109
timestamp 21601
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_110
timestamp 21601
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_111
timestamp 21601
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_112
timestamp 21601
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_113
timestamp 21601
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_114
timestamp 21601
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_115
timestamp 21601
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_116
timestamp 21601
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_117
timestamp 21601
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_118
timestamp 21601
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_119
timestamp 21601
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_120
timestamp 21601
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_121
timestamp 21601
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_122
timestamp 21601
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_123
timestamp 21601
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_124
timestamp 21601
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_125
timestamp 21601
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_126
timestamp 21601
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_127
timestamp 21601
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_128
timestamp 21601
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_129
timestamp 21601
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_130
timestamp 21601
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_131
timestamp 21601
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_132
timestamp 21601
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_133
timestamp 21601
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_134
timestamp 21601
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_135
timestamp 21601
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_136
timestamp 21601
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_137
timestamp 21601
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_138
timestamp 21601
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_139
timestamp 21601
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_140
timestamp 21601
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_141
timestamp 21601
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_142
timestamp 21601
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_143
timestamp 21601
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_144
timestamp 21601
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_145
timestamp 21601
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_146
timestamp 21601
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_147
timestamp 21601
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_148
timestamp 21601
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_149
timestamp 21601
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_150
timestamp 21601
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_151
timestamp 21601
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_152
timestamp 21601
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_153
timestamp 21601
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_154
timestamp 21601
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_155
timestamp 21601
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_156
timestamp 21601
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_157
timestamp 21601
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_158
timestamp 21601
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_159
timestamp 21601
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_160
timestamp 21601
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_161
timestamp 21601
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_162
timestamp 21601
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_163
timestamp 21601
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_164
timestamp 21601
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_165
timestamp 21601
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_166
timestamp 21601
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_167
timestamp 21601
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_168
timestamp 21601
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_169
timestamp 21601
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_170
timestamp 21601
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_171
timestamp 21601
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_172
timestamp 21601
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_173
timestamp 21601
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_174
timestamp 21601
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_175
timestamp 21601
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_176
timestamp 21601
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_177
timestamp 21601
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_178
timestamp 21601
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_179
timestamp 21601
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_180
timestamp 21601
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_181
timestamp 21601
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_182
timestamp 21601
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_183
timestamp 21601
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_184
timestamp 21601
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_185
timestamp 21601
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_186
timestamp 21601
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_187
timestamp 21601
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_188
timestamp 21601
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_189
timestamp 21601
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_190
timestamp 21601
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_191
timestamp 21601
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_192
timestamp 21601
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_193
timestamp 21601
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_194
timestamp 21601
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_195
timestamp 21601
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_196
timestamp 21601
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_197
timestamp 21601
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_198
timestamp 21601
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_199
timestamp 21601
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_200
timestamp 21601
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_201
timestamp 21601
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_202
timestamp 21601
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_203
timestamp 21601
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_204
timestamp 21601
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_205
timestamp 21601
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_206
timestamp 21601
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_207
timestamp 21601
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_208
timestamp 21601
transform 1 0 3680 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_209
timestamp 21601
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_210
timestamp 21601
transform 1 0 8832 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_211
timestamp 21601
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_212
timestamp 21601
transform 1 0 13984 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_213
timestamp 21601
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_214
timestamp 21601
transform 1 0 19136 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_215
timestamp 21601
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_31_216
timestamp 21601
transform 1 0 24288 0 -1 18496
box -38 -48 130 592
<< labels >>
flabel metal2 s 8208 1040 8528 18544 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 16208 1040 16528 18544 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 24208 1040 24528 18544 0 FreeSans 1792 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 1056 8210 24888 8530 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal3 s 1056 16210 24888 16530 0 FreeSans 1920 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal2 s 4208 1040 4528 18544 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 12208 1040 12528 18544 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 20208 1040 20528 18544 0 FreeSans 1792 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 1056 4210 24888 4530 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 1056 12210 24888 12530 0 FreeSans 1920 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal2 s 11610 19200 11666 20000 0 FreeSans 224 90 0 0 clockp[0]
port 2 nsew signal output
flabel metal2 s 14186 19200 14242 20000 0 FreeSans 224 90 0 0 clockp[1]
port 3 nsew signal output
flabel metal2 s 20350 0 20406 800 0 FreeSans 224 90 0 0 dco
port 4 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 div[0]
port 5 nsew signal input
flabel metal2 s 3422 0 3478 800 0 FreeSans 224 90 0 0 div[1]
port 6 nsew signal input
flabel metal2 s 5538 0 5594 800 0 FreeSans 224 90 0 0 div[2]
port 7 nsew signal input
flabel metal2 s 7654 0 7710 800 0 FreeSans 224 90 0 0 div[3]
port 8 nsew signal input
flabel metal2 s 9770 0 9826 800 0 FreeSans 224 90 0 0 div[4]
port 9 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 div[5]
port 10 nsew signal input
flabel metal2 s 14002 0 14058 800 0 FreeSans 224 90 0 0 div[6]
port 11 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 div[7]
port 12 nsew signal input
flabel metal2 s 18234 0 18290 800 0 FreeSans 224 90 0 0 enable
port 13 nsew signal input
flabel metal3 s 0 1096 800 1216 0 FreeSans 480 0 0 0 ext_trim[0]
port 14 nsew signal input
flabel metal2 s 3882 19200 3938 20000 0 FreeSans 224 90 0 0 ext_trim[10]
port 15 nsew signal input
flabel metal2 s 6458 19200 6514 20000 0 FreeSans 224 90 0 0 ext_trim[11]
port 16 nsew signal input
flabel metal2 s 9034 19200 9090 20000 0 FreeSans 224 90 0 0 ext_trim[12]
port 17 nsew signal input
flabel metal2 s 16762 19200 16818 20000 0 FreeSans 224 90 0 0 ext_trim[13]
port 18 nsew signal input
flabel metal2 s 19338 19200 19394 20000 0 FreeSans 224 90 0 0 ext_trim[14]
port 19 nsew signal input
flabel metal2 s 21914 19200 21970 20000 0 FreeSans 224 90 0 0 ext_trim[15]
port 20 nsew signal input
flabel metal2 s 24490 19200 24546 20000 0 FreeSans 224 90 0 0 ext_trim[16]
port 21 nsew signal input
flabel metal3 s 25200 18504 26000 18624 0 FreeSans 480 0 0 0 ext_trim[17]
port 22 nsew signal input
flabel metal3 s 25200 16328 26000 16448 0 FreeSans 480 0 0 0 ext_trim[18]
port 23 nsew signal input
flabel metal3 s 25200 14152 26000 14272 0 FreeSans 480 0 0 0 ext_trim[19]
port 24 nsew signal input
flabel metal3 s 0 3272 800 3392 0 FreeSans 480 0 0 0 ext_trim[1]
port 25 nsew signal input
flabel metal3 s 25200 11976 26000 12096 0 FreeSans 480 0 0 0 ext_trim[20]
port 26 nsew signal input
flabel metal3 s 25200 9800 26000 9920 0 FreeSans 480 0 0 0 ext_trim[21]
port 27 nsew signal input
flabel metal3 s 25200 7624 26000 7744 0 FreeSans 480 0 0 0 ext_trim[22]
port 28 nsew signal input
flabel metal3 s 25200 5448 26000 5568 0 FreeSans 480 0 0 0 ext_trim[23]
port 29 nsew signal input
flabel metal3 s 25200 3272 26000 3392 0 FreeSans 480 0 0 0 ext_trim[24]
port 30 nsew signal input
flabel metal3 s 25200 1096 26000 1216 0 FreeSans 480 0 0 0 ext_trim[25]
port 31 nsew signal input
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 ext_trim[2]
port 32 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 ext_trim[3]
port 33 nsew signal input
flabel metal3 s 0 9800 800 9920 0 FreeSans 480 0 0 0 ext_trim[4]
port 34 nsew signal input
flabel metal3 s 0 11976 800 12096 0 FreeSans 480 0 0 0 ext_trim[5]
port 35 nsew signal input
flabel metal3 s 0 14152 800 14272 0 FreeSans 480 0 0 0 ext_trim[6]
port 36 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 ext_trim[7]
port 37 nsew signal input
flabel metal3 s 0 18504 800 18624 0 FreeSans 480 0 0 0 ext_trim[8]
port 38 nsew signal input
flabel metal2 s 1306 19200 1362 20000 0 FreeSans 224 90 0 0 ext_trim[9]
port 39 nsew signal input
flabel metal2 s 24582 0 24638 800 0 FreeSans 224 90 0 0 osc
port 40 nsew signal input
flabel metal2 s 22466 0 22522 800 0 FreeSans 224 90 0 0 resetb
port 41 nsew signal input
rlabel metal1 12972 18496 12972 18496 0 VGND
rlabel metal1 12972 17952 12972 17952 0 VPWR
rlabel metal2 15226 8738 15226 8738 0 _000_
rlabel metal1 14720 7514 14720 7514 0 _001_
rlabel metal1 9568 9418 9568 9418 0 _002_
rlabel metal2 9522 13294 9522 13294 0 _003_
rlabel metal2 18538 11016 18538 11016 0 _004_
rlabel metal1 17986 10234 17986 10234 0 _005_
rlabel metal1 17710 12342 17710 12342 0 _006_
rlabel metal2 17986 11390 17986 11390 0 _007_
rlabel metal2 4002 14552 4002 14552 0 _008_
rlabel metal1 9108 14246 9108 14246 0 _009_
rlabel metal2 5934 11288 5934 11288 0 _010_
rlabel metal2 18814 8942 18814 8942 0 _011_
rlabel metal2 19734 5032 19734 5032 0 _012_
rlabel metal1 17993 6698 17993 6698 0 _013_
rlabel metal1 2668 18054 2668 18054 0 _014_
rlabel metal2 6854 16966 6854 16966 0 _015_
rlabel metal1 2254 9656 2254 9656 0 _016_
rlabel metal2 23506 9384 23506 9384 0 _017_
rlabel metal2 20102 1122 20102 1122 0 _018_
rlabel metal1 24012 5338 24012 5338 0 _019_
rlabel metal2 2898 13736 2898 13736 0 _020_
rlabel metal1 8885 11798 8885 11798 0 _021_
rlabel metal1 6164 12614 6164 12614 0 _022_
rlabel metal1 18085 8874 18085 8874 0 _023_
rlabel metal2 17986 5406 17986 5406 0 _024_
rlabel metal1 15272 7174 15272 7174 0 _025_
rlabel metal2 5750 17204 5750 17204 0 _026_
rlabel metal2 7958 17816 7958 17816 0 _027_
rlabel metal2 2990 10982 2990 10982 0 _028_
rlabel metal1 22724 9146 22724 9146 0 _029_
rlabel metal2 21666 4556 21666 4556 0 _030_
rlabel metal2 21390 7514 21390 7514 0 _031_
rlabel metal1 4600 7514 4600 7514 0 _032_
rlabel metal2 5106 10472 5106 10472 0 _033_
rlabel metal2 5014 9384 5014 9384 0 _034_
rlabel metal2 8786 8670 8786 8670 0 _035_
rlabel metal1 12834 7480 12834 7480 0 _036_
rlabel metal2 7958 10200 7958 10200 0 _037_
rlabel metal2 2806 16762 2806 16762 0 _038_
rlabel metal2 6026 14552 6026 14552 0 _039_
rlabel metal2 2162 8738 2162 8738 0 _040_
rlabel metal1 24058 8364 24058 8364 0 _041_
rlabel metal1 21942 3128 21942 3128 0 _042_
rlabel metal1 23874 2074 23874 2074 0 _043_
rlabel metal1 5336 15674 5336 15674 0 _044_
rlabel metal1 7636 14586 7636 14586 0 _045_
rlabel metal2 3726 12172 3726 12172 0 _046_
rlabel metal1 20240 8602 20240 8602 0 _047_
rlabel metal1 20424 3910 20424 3910 0 _048_
rlabel metal1 18584 7718 18584 7718 0 _049_
rlabel metal1 22188 2006 22188 2006 0 _050_
rlabel metal1 22678 4998 22678 4998 0 _051_
rlabel metal1 18400 1190 18400 1190 0 _052_
rlabel metal2 2530 14552 2530 14552 0 _053_
rlabel metal1 6486 14008 6486 14008 0 _054_
rlabel metal1 2438 6664 2438 6664 0 _055_
rlabel metal2 24058 6936 24058 6936 0 _056_
rlabel metal2 18262 3672 18262 3672 0 _057_
rlabel metal1 20976 5338 20976 5338 0 _058_
rlabel metal1 4646 16694 4646 16694 0 _059_
rlabel metal1 8556 16422 8556 16422 0 _060_
rlabel metal1 2622 12682 2622 12682 0 _061_
rlabel metal1 21528 9418 21528 9418 0 _062_
rlabel metal1 23966 3638 23966 3638 0 _063_
rlabel metal1 21206 7480 21206 7480 0 _064_
rlabel metal2 1978 1768 1978 1768 0 _065_
rlabel metal1 2392 3706 2392 3706 0 _066_
rlabel metal1 6118 3162 6118 3162 0 _067_
rlabel metal2 7406 3944 7406 3944 0 _068_
rlabel metal1 14490 2074 14490 2074 0 _069_
rlabel metal2 15594 6800 15594 6800 0 _070_
rlabel metal1 17289 4182 17289 4182 0 _071_
rlabel metal1 17342 1530 17342 1530 0 _072_
rlabel metal1 6762 2074 6762 2074 0 _073_
rlabel metal2 14398 8738 14398 8738 0 _074_
rlabel metal1 13984 7922 13984 7922 0 _075_
rlabel metal1 9430 9146 9430 9146 0 _076_
rlabel metal1 9016 12750 9016 12750 0 _077_
rlabel metal1 17434 11662 17434 11662 0 _078_
rlabel metal1 16468 10778 16468 10778 0 _079_
rlabel metal1 16974 12750 16974 12750 0 _080_
rlabel metal1 16192 10234 16192 10234 0 _081_
rlabel metal2 3910 14756 3910 14756 0 _082_
rlabel metal1 7636 13498 7636 13498 0 _083_
rlabel metal1 6670 11186 6670 11186 0 _084_
rlabel metal2 17250 8942 17250 8942 0 _085_
rlabel metal1 19412 5270 19412 5270 0 _086_
rlabel metal2 16790 6562 16790 6562 0 _087_
rlabel metal1 2254 17306 2254 17306 0 _088_
rlabel metal1 7912 16762 7912 16762 0 _089_
rlabel metal2 2530 9894 2530 9894 0 _090_
rlabel metal2 22862 10030 22862 10030 0 _091_
rlabel via1 20095 1530 20095 1530 0 _092_
rlabel metal1 22310 6392 22310 6392 0 _093_
rlabel metal1 2208 13430 2208 13430 0 _094_
rlabel metal2 7406 11560 7406 11560 0 _095_
rlabel metal1 5290 11866 5290 11866 0 _096_
rlabel metal2 16606 9112 16606 9112 0 _097_
rlabel metal2 17342 4964 17342 4964 0 _098_
rlabel metal1 14582 6426 14582 6426 0 _099_
rlabel metal2 4646 17884 4646 17884 0 _100_
rlabel metal1 8648 17306 8648 17306 0 _101_
rlabel metal2 1978 10846 1978 10846 0 _102_
rlabel metal2 21942 10200 21942 10200 0 _103_
rlabel metal1 24012 2958 24012 2958 0 _104_
rlabel metal1 20230 6970 20230 6970 0 _105_
rlabel metal1 6164 7786 6164 7786 0 _106_
rlabel metal2 5382 10404 5382 10404 0 _107_
rlabel metal2 5290 9316 5290 9316 0 _108_
rlabel metal2 7774 8670 7774 8670 0 _109_
rlabel metal2 9522 7582 9522 7582 0 _110_
rlabel metal2 6946 9826 6946 9826 0 _111_
rlabel metal1 2070 16218 2070 16218 0 _112_
rlabel metal1 5428 14314 5428 14314 0 _113_
rlabel metal1 2346 8602 2346 8602 0 _114_
rlabel metal1 22632 8058 22632 8058 0 _115_
rlabel metal1 20378 2958 20378 2958 0 _116_
rlabel metal1 22770 5338 22770 5338 0 _117_
rlabel metal1 4508 15674 4508 15674 0 _118_
rlabel metal2 7866 14756 7866 14756 0 _119_
rlabel metal1 2691 11798 2691 11798 0 _120_
rlabel metal2 19366 8738 19366 8738 0 _121_
rlabel metal1 20240 4250 20240 4250 0 _122_
rlabel metal2 17434 7582 17434 7582 0 _123_
rlabel metal2 1794 14824 1794 14824 0 _124_
rlabel metal2 6210 13600 6210 13600 0 _125_
rlabel metal1 1794 7480 1794 7480 0 _126_
rlabel metal2 22586 7582 22586 7582 0 _127_
rlabel metal1 18492 3162 18492 3162 0 _128_
rlabel metal2 22034 6222 22034 6222 0 _129_
rlabel metal2 4738 16932 4738 16932 0 _130_
rlabel metal2 7958 15844 7958 15844 0 _131_
rlabel metal1 2530 12614 2530 12614 0 _132_
rlabel metal2 20010 9690 20010 9690 0 _133_
rlabel metal2 22586 3876 22586 3876 0 _134_
rlabel metal2 19458 7582 19458 7582 0 _135_
rlabel metal2 2714 2244 2714 2244 0 _136_
rlabel metal1 2024 4182 2024 4182 0 _137_
rlabel metal2 5198 3672 5198 3672 0 _138_
rlabel metal1 6900 4182 6900 4182 0 _139_
rlabel metal1 9522 3570 9522 3570 0 _140_
rlabel metal1 12190 5882 12190 5882 0 _141_
rlabel metal1 16744 3706 16744 3706 0 _142_
rlabel metal2 17066 2244 17066 2244 0 _143_
rlabel metal1 7820 2006 7820 2006 0 _144_
rlabel metal2 22126 1122 22126 1122 0 _145_
rlabel metal1 19642 1326 19642 1326 0 _146_
rlabel metal2 2346 2142 2346 2142 0 _147_
rlabel metal2 1794 6698 1794 6698 0 _148_
rlabel metal1 1978 6324 1978 6324 0 _149_
rlabel metal1 16284 12818 16284 12818 0 _150_
rlabel metal1 11362 7888 11362 7888 0 _151_
rlabel metal1 11086 13158 11086 13158 0 _152_
rlabel metal1 11822 11084 11822 11084 0 _153_
rlabel via1 3634 1173 3634 1173 0 _154_
rlabel metal1 15364 2006 15364 2006 0 _155_
rlabel metal1 18676 2618 18676 2618 0 _156_
rlabel metal1 16330 1904 16330 1904 0 _157_
rlabel metal1 21666 3706 21666 3706 0 _158_
rlabel metal1 15916 2482 15916 2482 0 _159_
rlabel metal1 15640 5134 15640 5134 0 _160_
rlabel metal2 14858 5406 14858 5406 0 _161_
rlabel metal1 15502 2482 15502 2482 0 _162_
rlabel metal1 14996 4046 14996 4046 0 _163_
rlabel metal1 13289 4556 13289 4556 0 _164_
rlabel metal1 14030 4590 14030 4590 0 _165_
rlabel metal2 11730 5066 11730 5066 0 _166_
rlabel metal2 13846 4998 13846 4998 0 _167_
rlabel via1 13588 4590 13588 4590 0 _168_
rlabel metal1 13754 5168 13754 5168 0 _169_
rlabel metal1 12926 4794 12926 4794 0 _170_
rlabel metal2 14950 3774 14950 3774 0 _171_
rlabel metal2 9338 6460 9338 6460 0 _172_
rlabel metal1 10120 6222 10120 6222 0 _173_
rlabel metal2 10258 6596 10258 6596 0 _174_
rlabel metal1 10396 4794 10396 4794 0 _175_
rlabel metal2 11270 4352 11270 4352 0 _176_
rlabel metal2 10442 4828 10442 4828 0 _177_
rlabel metal2 10994 3740 10994 3740 0 _178_
rlabel metal1 11408 3026 11408 3026 0 _179_
rlabel metal1 10902 4114 10902 4114 0 _180_
rlabel metal1 6164 6970 6164 6970 0 _181_
rlabel metal2 6670 6902 6670 6902 0 _182_
rlabel metal2 5934 7072 5934 7072 0 _183_
rlabel metal1 7590 6324 7590 6324 0 _184_
rlabel metal1 8234 6426 8234 6426 0 _185_
rlabel metal2 7866 6562 7866 6562 0 _186_
rlabel metal1 7360 5202 7360 5202 0 _187_
rlabel metal2 7314 4420 7314 4420 0 _188_
rlabel metal2 8694 6188 8694 6188 0 _189_
rlabel metal1 3818 6324 3818 6324 0 _190_
rlabel metal2 2346 6086 2346 6086 0 _191_
rlabel metal2 5198 6528 5198 6528 0 _192_
rlabel metal1 2622 6256 2622 6256 0 _193_
rlabel metal2 5474 6018 5474 6018 0 _194_
rlabel via1 5566 5678 5566 5678 0 _195_
rlabel metal2 5750 6426 5750 6426 0 _196_
rlabel metal1 6762 5610 6762 5610 0 _197_
rlabel metal2 7406 5440 7406 5440 0 _198_
rlabel metal1 3634 5168 3634 5168 0 _199_
rlabel metal1 3036 5678 3036 5678 0 _200_
rlabel metal1 2530 5202 2530 5202 0 _201_
rlabel metal2 2254 3978 2254 3978 0 _202_
rlabel metal2 3542 4794 3542 4794 0 _203_
rlabel metal1 3174 3502 3174 3502 0 _204_
rlabel metal1 3496 4250 3496 4250 0 _205_
rlabel metal1 5888 5134 5888 5134 0 _206_
rlabel metal1 7498 5100 7498 5100 0 _207_
rlabel metal1 7544 5610 7544 5610 0 _208_
rlabel metal2 10718 4896 10718 4896 0 _209_
rlabel metal1 15318 4522 15318 4522 0 _210_
rlabel metal1 13294 4114 13294 4114 0 _211_
rlabel metal1 13708 3910 13708 3910 0 _212_
rlabel metal1 15088 3026 15088 3026 0 _213_
rlabel metal1 15272 2890 15272 2890 0 _214_
rlabel via1 15962 2363 15962 2363 0 _215_
rlabel metal1 16422 5202 16422 5202 0 _216_
rlabel metal1 17756 1462 17756 1462 0 _217_
rlabel metal2 15226 3196 15226 3196 0 _218_
rlabel metal1 13570 3060 13570 3060 0 _219_
rlabel metal2 13294 2380 13294 2380 0 _220_
rlabel metal1 4830 1394 4830 1394 0 _221_
rlabel metal1 8188 2482 8188 2482 0 _222_
rlabel metal1 4554 3060 4554 3060 0 _223_
rlabel metal2 16146 4692 16146 4692 0 _224_
rlabel metal2 16698 3740 16698 3740 0 _225_
rlabel metal1 16376 2482 16376 2482 0 _226_
rlabel metal1 17572 1530 17572 1530 0 _227_
rlabel metal2 16054 3298 16054 3298 0 _228_
rlabel metal1 12466 5644 12466 5644 0 _229_
rlabel metal2 12650 5508 12650 5508 0 _230_
rlabel metal1 10212 4114 10212 4114 0 _231_
rlabel metal1 10074 4080 10074 4080 0 _232_
rlabel metal1 7084 4658 7084 4658 0 _233_
rlabel metal2 7038 4794 7038 4794 0 _234_
rlabel metal1 5060 4794 5060 4794 0 _235_
rlabel metal2 5290 4556 5290 4556 0 _236_
rlabel metal2 5382 4284 5382 4284 0 _237_
rlabel via2 2990 4675 2990 4675 0 _238_
rlabel metal2 2668 3638 2668 3638 0 _239_
rlabel metal1 4278 4114 4278 4114 0 _240_
rlabel metal1 2438 2516 2438 2516 0 _241_
rlabel viali 7490 7446 7490 7446 0 _242_
rlabel metal1 8418 7888 8418 7888 0 _243_
rlabel metal2 7406 8194 7406 8194 0 _244_
rlabel metal1 9246 7820 9246 7820 0 _245_
rlabel metal2 7222 8704 7222 8704 0 _246_
rlabel via1 7153 8874 7153 8874 0 _247_
rlabel metal1 6072 8942 6072 8942 0 _248_
rlabel via1 5819 8942 5819 8942 0 _249_
rlabel metal1 7038 10642 7038 10642 0 _250_
rlabel metal2 5842 10268 5842 10268 0 _251_
rlabel metal1 7452 6426 7452 6426 0 _252_
rlabel metal1 10442 1360 10442 1360 0 _253_
rlabel metal1 7774 2380 7774 2380 0 _254_
rlabel via2 8878 2499 8878 2499 0 _255_
rlabel metal2 12926 3740 12926 3740 0 _256_
rlabel metal1 12788 4590 12788 4590 0 _257_
rlabel metal2 12650 3638 12650 3638 0 _258_
rlabel metal1 11040 1734 11040 1734 0 _259_
rlabel metal1 12466 2006 12466 2006 0 _260_
rlabel metal1 11914 1904 11914 1904 0 _261_
rlabel metal1 13202 2448 13202 2448 0 _262_
rlabel metal1 11316 2890 11316 2890 0 _263_
rlabel metal1 13110 3162 13110 3162 0 _264_
rlabel metal1 14398 5576 14398 5576 0 _265_
rlabel via2 11086 1309 11086 1309 0 _266_
rlabel metal1 10672 2414 10672 2414 0 _267_
rlabel metal1 11500 6766 11500 6766 0 _268_
rlabel metal1 7268 2414 7268 2414 0 _269_
rlabel metal2 6854 1904 6854 1904 0 _270_
rlabel metal1 5842 2482 5842 2482 0 _271_
rlabel metal1 6716 1530 6716 1530 0 _272_
rlabel metal1 5796 2414 5796 2414 0 _273_
rlabel metal2 6762 2244 6762 2244 0 _274_
rlabel metal1 3588 1938 3588 1938 0 _275_
rlabel metal2 3082 1938 3082 1938 0 _276_
rlabel metal2 4002 2244 4002 2244 0 _277_
rlabel metal1 4554 2074 4554 2074 0 _278_
rlabel metal1 3450 2584 3450 2584 0 _279_
rlabel metal1 10994 6188 10994 6188 0 _280_
rlabel metal1 11776 7854 11776 7854 0 _281_
rlabel metal1 12006 8942 12006 8942 0 _282_
rlabel metal1 15042 10642 15042 10642 0 _283_
rlabel metal1 14306 9350 14306 9350 0 _284_
rlabel metal1 14398 9588 14398 9588 0 _285_
rlabel metal1 13386 11696 13386 11696 0 _286_
rlabel metal1 13662 11764 13662 11764 0 _287_
rlabel metal1 10626 11186 10626 11186 0 _288_
rlabel metal1 11316 8466 11316 8466 0 _289_
rlabel metal1 10577 8942 10577 8942 0 _290_
rlabel metal1 14858 6154 14858 6154 0 _291_
rlabel metal1 13202 9384 13202 9384 0 _292_
rlabel metal2 12926 9656 12926 9656 0 _293_
rlabel metal1 10350 7922 10350 7922 0 _294_
rlabel metal2 10534 8262 10534 8262 0 _295_
rlabel metal2 10810 9792 10810 9792 0 _296_
rlabel metal2 9982 12002 9982 12002 0 _297_
rlabel metal1 13294 11152 13294 11152 0 _298_
rlabel metal1 14674 11730 14674 11730 0 _299_
rlabel metal1 15686 9690 15686 9690 0 _300_
rlabel metal1 15134 9554 15134 9554 0 _301_
rlabel metal1 15226 10166 15226 10166 0 _302_
rlabel metal1 13202 12818 13202 12818 0 _303_
rlabel metal1 15318 14314 15318 14314 0 _304_
rlabel metal1 11684 9554 11684 9554 0 _305_
rlabel metal2 12650 9792 12650 9792 0 _306_
rlabel metal1 22172 14994 22172 14994 0 _307_
rlabel metal1 13386 10166 13386 10166 0 _308_
rlabel metal2 13754 11356 13754 11356 0 _309_
rlabel metal2 13386 10268 13386 10268 0 _310_
rlabel via1 6762 1819 6762 1819 0 _311_
rlabel metal2 9062 2176 9062 2176 0 _312_
rlabel metal1 16054 12614 16054 12614 0 _313_
rlabel metal2 12650 10438 12650 10438 0 _314_
rlabel metal1 14674 12614 14674 12614 0 _315_
rlabel metal2 15226 12206 15226 12206 0 _316_
rlabel metal1 15410 11764 15410 11764 0 _317_
rlabel metal1 15916 12682 15916 12682 0 _318_
rlabel metal1 16054 12750 16054 12750 0 _319_
rlabel metal1 16422 10676 16422 10676 0 _320_
rlabel metal1 16100 10574 16100 10574 0 _321_
rlabel metal1 14950 9418 14950 9418 0 _322_
rlabel metal1 12190 12206 12190 12206 0 _323_
rlabel metal1 13478 11322 13478 11322 0 _324_
rlabel metal2 10350 11900 10350 11900 0 _325_
rlabel metal2 10810 11492 10810 11492 0 _326_
rlabel metal2 9522 12002 9522 12002 0 _327_
rlabel metal1 9890 8976 9890 8976 0 _328_
rlabel metal1 10143 9146 10143 9146 0 _329_
rlabel metal2 9430 9996 9430 9996 0 _330_
rlabel metal1 14996 7378 14996 7378 0 _331_
rlabel metal1 14904 8058 14904 8058 0 _332_
rlabel metal1 13018 8364 13018 8364 0 _333_
rlabel metal2 12098 13056 12098 13056 0 _334_
rlabel metal1 14582 14348 14582 14348 0 _335_
rlabel metal1 16192 14042 16192 14042 0 _336_
rlabel metal1 12742 14586 12742 14586 0 _337_
rlabel metal2 16974 13702 16974 13702 0 _338_
rlabel metal2 16790 14144 16790 14144 0 _339_
rlabel metal1 14030 15096 14030 15096 0 _340_
rlabel metal2 11822 14790 11822 14790 0 _341_
rlabel metal1 10488 14314 10488 14314 0 _342_
rlabel metal2 13294 14229 13294 14229 0 _343_
rlabel metal1 10994 13906 10994 13906 0 _344_
rlabel metal2 17342 14756 17342 14756 0 _345_
rlabel metal1 15088 15334 15088 15334 0 _346_
rlabel metal1 15410 14416 15410 14416 0 _347_
rlabel metal1 16192 16558 16192 16558 0 _348_
rlabel metal2 10258 16320 10258 16320 0 _349_
rlabel metal2 10166 15436 10166 15436 0 _350_
rlabel metal2 16054 16490 16054 16490 0 _351_
rlabel metal1 19642 16116 19642 16116 0 _352_
rlabel metal1 20528 11798 20528 11798 0 _353_
rlabel metal1 15916 15130 15916 15130 0 _354_
rlabel metal2 15318 16337 15318 16337 0 _355_
rlabel metal1 21482 15538 21482 15538 0 _356_
rlabel metal1 21712 14994 21712 14994 0 _357_
rlabel metal1 20746 16218 20746 16218 0 _358_
rlabel metal1 20608 15674 20608 15674 0 _359_
rlabel metal2 21482 15674 21482 15674 0 _360_
rlabel metal1 21390 11118 21390 11118 0 _361_
rlabel metal2 21022 12036 21022 12036 0 _362_
rlabel metal1 11316 17714 11316 17714 0 clockp[0]
rlabel metal2 20654 18088 20654 18088 0 clockp[1]
rlabel metal1 23966 1394 23966 1394 0 clockp_buffer_in\[0\]
rlabel metal1 19182 17578 19182 17578 0 clockp_buffer_in\[1\]
rlabel metal2 20654 1581 20654 1581 0 dco
rlabel metal1 1702 2380 1702 2380 0 div[0]
rlabel metal1 3680 8466 3680 8466 0 div[1]
rlabel metal1 4784 3502 4784 3502 0 div[2]
rlabel metal1 4692 1326 4692 1326 0 div[3]
rlabel metal2 9798 1761 9798 1761 0 div[4]
rlabel metal1 11776 1326 11776 1326 0 div[5]
rlabel metal1 14122 1326 14122 1326 0 div[6]
rlabel metal2 16146 1761 16146 1761 0 div[7]
rlabel metal1 2898 3604 2898 3604 0 dll_control.accum\[0\]
rlabel metal1 4922 1938 4922 1938 0 dll_control.accum\[1\]
rlabel metal1 5842 1258 5842 1258 0 dll_control.accum\[2\]
rlabel metal2 7866 1428 7866 1428 0 dll_control.accum\[3\]
rlabel metal1 12604 3978 12604 3978 0 dll_control.accum\[4\]
rlabel metal2 12650 1853 12650 1853 0 dll_control.accum\[5\]
rlabel metal2 15778 1870 15778 1870 0 dll_control.accum\[6\]
rlabel metal1 11362 3502 11362 3502 0 dll_control.accum\[7\]
rlabel metal1 9706 1938 9706 1938 0 dll_control.accum\[8\]
rlabel metal2 2070 5372 2070 5372 0 dll_control.count0\[0\]
rlabel metal1 1702 6358 1702 6358 0 dll_control.count0\[1\]
rlabel metal1 5980 9486 5980 9486 0 dll_control.count0\[2\]
rlabel metal1 15318 8568 15318 8568 0 dll_control.count0\[3\]
rlabel metal1 9522 7854 9522 7854 0 dll_control.count0\[4\]
rlabel metal1 8142 10098 8142 10098 0 dll_control.count0\[5\]
rlabel metal2 3358 14144 3358 14144 0 dll_control.count1\[0\]
rlabel metal1 8234 13226 8234 13226 0 dll_control.count1\[1\]
rlabel metal1 6670 12104 6670 12104 0 dll_control.count1\[2\]
rlabel metal1 17710 9622 17710 9622 0 dll_control.count1\[3\]
rlabel metal1 18906 5338 18906 5338 0 dll_control.count1\[4\]
rlabel metal1 16606 6630 16606 6630 0 dll_control.count1\[5\]
rlabel metal1 4784 15130 4784 15130 0 dll_control.count2\[0\]
rlabel metal1 8510 14042 8510 14042 0 dll_control.count2\[1\]
rlabel metal1 4370 12342 4370 12342 0 dll_control.count2\[2\]
rlabel metal2 18722 9078 18722 9078 0 dll_control.count2\[3\]
rlabel metal2 20746 5882 20746 5882 0 dll_control.count2\[4\]
rlabel metal1 18032 6970 18032 6970 0 dll_control.count2\[5\]
rlabel metal1 5520 15946 5520 15946 0 dll_control.count3\[0\]
rlabel metal2 8878 15232 8878 15232 0 dll_control.count3\[1\]
rlabel metal1 3726 12206 3726 12206 0 dll_control.count3\[2\]
rlabel metal1 20424 8806 20424 8806 0 dll_control.count3\[3\]
rlabel metal2 21758 4012 21758 4012 0 dll_control.count3\[4\]
rlabel metal1 19366 7514 19366 7514 0 dll_control.count3\[5\]
rlabel metal1 5566 17034 5566 17034 0 dll_control.count4\[0\]
rlabel metal2 8970 16660 8970 16660 0 dll_control.count4\[1\]
rlabel metal1 3174 12886 3174 12886 0 dll_control.count4\[2\]
rlabel metal1 21528 9486 21528 9486 0 dll_control.count4\[3\]
rlabel metal2 23322 3978 23322 3978 0 dll_control.count4\[4\]
rlabel metal1 20378 7786 20378 7786 0 dll_control.count4\[5\]
rlabel metal2 5290 17782 5290 17782 0 dll_control.count5\[0\]
rlabel metal2 7406 17068 7406 17068 0 dll_control.count5\[1\]
rlabel metal1 3174 10778 3174 10778 0 dll_control.count5\[2\]
rlabel metal1 22908 10710 22908 10710 0 dll_control.count5\[3\]
rlabel metal1 21160 2482 21160 2482 0 dll_control.count5\[4\]
rlabel metal1 21390 6970 21390 6970 0 dll_control.count5\[5\]
rlabel metal1 3128 17306 3128 17306 0 dll_control.count6\[0\]
rlabel metal1 7130 16558 7130 16558 0 dll_control.count6\[1\]
rlabel metal2 2898 9792 2898 9792 0 dll_control.count6\[2\]
rlabel metal1 23874 9486 23874 9486 0 dll_control.count6\[3\]
rlabel metal1 21344 1530 21344 1530 0 dll_control.count6\[4\]
rlabel metal1 23552 6086 23552 6086 0 dll_control.count6\[5\]
rlabel metal2 2714 16320 2714 16320 0 dll_control.count7\[0\]
rlabel metal2 6762 13804 6762 13804 0 dll_control.count7\[1\]
rlabel metal1 3082 8602 3082 8602 0 dll_control.count7\[2\]
rlabel metal2 23322 8092 23322 8092 0 dll_control.count7\[3\]
rlabel metal1 20654 3162 20654 3162 0 dll_control.count7\[4\]
rlabel metal1 23138 5338 23138 5338 0 dll_control.count7\[5\]
rlabel metal1 2668 15334 2668 15334 0 dll_control.count8\[0\]
rlabel metal1 4186 13702 4186 13702 0 dll_control.count8\[1\]
rlabel metal2 3266 7616 3266 7616 0 dll_control.count8\[2\]
rlabel metal1 22632 7786 22632 7786 0 dll_control.count8\[3\]
rlabel metal1 17250 3400 17250 3400 0 dll_control.count8\[4\]
rlabel metal1 20010 5882 20010 5882 0 dll_control.count8\[5\]
rlabel metal2 22034 1632 22034 1632 0 dll_control.oscbuf\[0\]
rlabel metal1 20194 1870 20194 1870 0 dll_control.oscbuf\[1\]
rlabel metal1 18814 2074 18814 2074 0 dll_control.oscbuf\[2\]
rlabel metal1 19826 13906 19826 13906 0 dll_control.tint\[0\]
rlabel metal1 23966 12716 23966 12716 0 dll_control.tint\[1\]
rlabel metal1 20378 15028 20378 15028 0 dll_control.tint\[2\]
rlabel metal1 19780 12954 19780 12954 0 dll_control.tint\[3\]
rlabel metal1 16238 15028 16238 15028 0 dll_control.tint\[4\]
rlabel via2 13202 7837 13202 7837 0 dll_control.tval\[0\]
rlabel metal1 13294 7820 13294 7820 0 dll_control.tval\[1\]
rlabel metal1 13340 10234 13340 10234 0 dll_control.tval\[2\]
rlabel metal2 18262 840 18262 840 0 enable
rlabel metal1 6440 1326 6440 1326 0 ext_trim[0]
rlabel metal1 3956 18258 3956 18258 0 ext_trim[10]
rlabel metal1 6532 18258 6532 18258 0 ext_trim[11]
rlabel metal1 9108 18258 9108 18258 0 ext_trim[12]
rlabel metal1 17158 17782 17158 17782 0 ext_trim[13]
rlabel metal1 20010 18292 20010 18292 0 ext_trim[14]
rlabel metal1 21528 14042 21528 14042 0 ext_trim[15]
rlabel metal2 24426 19193 24426 19193 0 ext_trim[16]
rlabel via2 23506 18581 23506 18581 0 ext_trim[17]
rlabel metal1 22954 14824 22954 14824 0 ext_trim[18]
rlabel metal1 24242 17306 24242 17306 0 ext_trim[19]
rlabel metal2 1518 2329 1518 2329 0 ext_trim[1]
rlabel metal1 24288 14994 24288 14994 0 ext_trim[20]
rlabel metal2 24150 9401 24150 9401 0 ext_trim[21]
rlabel metal2 21666 9078 21666 9078 0 ext_trim[22]
rlabel metal3 24388 5508 24388 5508 0 ext_trim[23]
rlabel metal2 18998 6392 18998 6392 0 ext_trim[24]
rlabel metal3 23560 1156 23560 1156 0 ext_trim[25]
rlabel metal1 1472 4794 1472 4794 0 ext_trim[2]
rlabel metal1 1472 7854 1472 7854 0 ext_trim[3]
rlabel metal1 1426 11730 1426 11730 0 ext_trim[4]
rlabel metal1 1426 12818 1426 12818 0 ext_trim[5]
rlabel metal1 1472 14994 1472 14994 0 ext_trim[6]
rlabel via2 1518 16099 1518 16099 0 ext_trim[7]
rlabel metal2 2990 18411 2990 18411 0 ext_trim[8]
rlabel metal1 1426 18258 1426 18258 0 ext_trim[9]
rlabel metal1 23966 16218 23966 16218 0 ireset
rlabel metal2 14490 15572 14490 15572 0 itrim\[0\]
rlabel metal1 22862 14892 22862 14892 0 itrim\[10\]
rlabel metal1 22310 17102 22310 17102 0 itrim\[11\]
rlabel metal1 21022 18258 21022 18258 0 itrim\[12\]
rlabel metal1 16238 17646 16238 17646 0 itrim\[13\]
rlabel metal2 15594 16966 15594 16966 0 itrim\[14\]
rlabel metal2 20930 16864 20930 16864 0 itrim\[15\]
rlabel metal1 17572 16694 17572 16694 0 itrim\[16\]
rlabel metal2 19366 15776 19366 15776 0 itrim\[17\]
rlabel metal2 17710 16660 17710 16660 0 itrim\[18\]
rlabel metal1 19918 14484 19918 14484 0 itrim\[19\]
rlabel metal2 13110 15878 13110 15878 0 itrim\[1\]
rlabel metal2 19366 11968 19366 11968 0 itrim\[20\]
rlabel metal1 22678 11186 22678 11186 0 itrim\[21\]
rlabel metal1 23690 12852 23690 12852 0 itrim\[22\]
rlabel metal1 24196 13838 24196 13838 0 itrim\[23\]
rlabel metal1 23000 15470 23000 15470 0 itrim\[24\]
rlabel metal2 22218 15606 22218 15606 0 itrim\[25\]
rlabel metal2 10718 15164 10718 15164 0 itrim\[2\]
rlabel metal2 11638 15810 11638 15810 0 itrim\[3\]
rlabel metal2 17342 15742 17342 15742 0 itrim\[4\]
rlabel metal1 16836 17170 16836 17170 0 itrim\[5\]
rlabel metal1 17894 13940 17894 13940 0 itrim\[6\]
rlabel metal1 18906 12784 18906 12784 0 itrim\[7\]
rlabel metal1 23230 13430 23230 13430 0 itrim\[8\]
rlabel metal1 20562 13226 20562 13226 0 itrim\[9\]
rlabel metal1 21988 2414 21988 2414 0 net1
rlabel metal1 16054 816 16054 816 0 net10
rlabel metal2 14122 8670 14122 8670 0 net101
rlabel metal2 13478 9214 13478 9214 0 net102
rlabel metal2 14674 8602 14674 8602 0 net103
rlabel metal1 5474 6290 5474 6290 0 net105
rlabel metal1 10856 4046 10856 4046 0 net106
rlabel metal1 19182 3706 19182 3706 0 net107
rlabel metal1 10657 1938 10657 1938 0 net108
rlabel metal2 13570 3842 13570 3842 0 net109
rlabel metal1 12880 13362 12880 13362 0 net11
rlabel metal1 11868 10710 11868 10710 0 net110
rlabel metal2 15134 11628 15134 11628 0 net111
rlabel metal1 9246 14994 9246 14994 0 net12
rlabel metal1 13202 18088 13202 18088 0 net13
rlabel metal1 9660 17170 9660 17170 0 net14
rlabel metal2 19458 17238 19458 17238 0 net15
rlabel via1 15663 16490 15663 16490 0 net16
rlabel metal2 21114 15572 21114 15572 0 net17
rlabel metal1 20148 16558 20148 16558 0 net18
rlabel metal2 13386 18530 13386 18530 0 net19
rlabel metal1 4048 1734 4048 1734 0 net2
rlabel metal2 22494 15045 22494 15045 0 net20
rlabel metal1 23874 18054 23874 18054 0 net21
rlabel metal2 1702 1088 1702 1088 0 net22
rlabel viali 20654 11733 20654 11733 0 net23
rlabel metal1 23828 9146 23828 9146 0 net24
rlabel metal1 22540 11730 22540 11730 0 net25
rlabel metal2 21574 3944 21574 3944 0 net26
rlabel metal1 21160 15062 21160 15062 0 net27
rlabel via1 22404 14994 22404 14994 0 net28
rlabel metal1 2116 3638 2116 3638 0 net29
rlabel metal1 4140 1802 4140 1802 0 net3
rlabel metal2 7774 8041 7774 8041 0 net30
rlabel metal1 17204 14994 17204 14994 0 net31
rlabel metal2 9798 13668 9798 13668 0 net32
rlabel metal1 2231 14858 2231 14858 0 net33
rlabel metal2 13846 15300 13846 15300 0 net34
rlabel metal1 10833 15470 10833 15470 0 net35
rlabel metal2 9154 16150 9154 16150 0 net36
rlabel metal1 23690 2006 23690 2006 0 net37
rlabel metal2 15962 1632 15962 1632 0 net38
rlabel metal2 12926 10370 12926 10370 0 net39
rlabel metal2 4692 1292 4692 1292 0 net4
rlabel metal1 5382 16626 5382 16626 0 net40
rlabel metal1 5980 15538 5980 15538 0 net41
rlabel metal1 8280 12886 8280 12886 0 net42
rlabel metal1 23414 2482 23414 2482 0 net43
rlabel metal1 23184 9690 23184 9690 0 net44
rlabel metal2 19734 14246 19734 14246 0 net45
rlabel metal1 20562 14994 20562 14994 0 net46
rlabel metal1 24242 12920 24242 12920 0 net47
rlabel metal2 1886 17782 1886 17782 0 net48
rlabel metal1 9522 13192 9522 13192 0 net49
rlabel metal2 5658 1530 5658 1530 0 net5
rlabel metal1 9522 14280 9522 14280 0 net50
rlabel metal1 24564 2006 24564 2006 0 net51
rlabel metal1 21666 7446 21666 7446 0 net52
rlabel metal1 19780 6222 19780 6222 0 net53
rlabel metal1 2270 17238 2270 17238 0 net54
rlabel metal1 7736 16422 7736 16422 0 net55
rlabel via1 2154 1258 2154 1258 0 net56
rlabel metal1 24185 2006 24185 2006 0 net57
rlabel metal1 19642 7888 19642 7888 0 net58
rlabel metal1 24564 16082 24564 16082 0 net59
rlabel metal1 12834 1326 12834 1326 0 net6
rlabel metal1 2300 16966 2300 16966 0 net60
rlabel metal1 8326 16728 8326 16728 0 net61
rlabel metal1 2208 1530 2208 1530 0 net62
rlabel metal1 24104 1734 24104 1734 0 net63
rlabel metal1 17112 1530 17112 1530 0 net64
rlabel metal1 23782 15878 23782 15878 0 net65
rlabel metal2 10626 16354 10626 16354 0 net66
rlabel metal1 22034 11016 22034 11016 0 net67
rlabel metal1 21298 12308 21298 12308 0 net68
rlabel metal1 2024 1326 2024 1326 0 net69
rlabel metal1 12052 1326 12052 1326 0 net7
rlabel metal1 17756 16082 17756 16082 0 net70
rlabel metal2 11270 9248 11270 9248 0 net71
rlabel metal2 13570 7820 13570 7820 0 net73
rlabel metal1 15318 13294 15318 13294 0 net74
rlabel metal2 14674 12988 14674 12988 0 net75
rlabel metal1 4554 2482 4554 2482 0 net76
rlabel metal1 13202 5712 13202 5712 0 net77
rlabel metal1 12926 6732 12926 6732 0 net78
rlabel metal2 12650 7344 12650 7344 0 net79
rlabel metal1 14674 1938 14674 1938 0 net8
rlabel metal1 8786 2924 8786 2924 0 net80
rlabel via1 4117 1326 4117 1326 0 net81
rlabel metal1 3910 5678 3910 5678 0 net82
rlabel via1 3817 7378 3817 7378 0 net83
rlabel metal1 17756 2618 17756 2618 0 net85
rlabel metal1 16790 4692 16790 4692 0 net86
rlabel metal1 16146 3536 16146 3536 0 net87
rlabel metal2 11960 7854 11960 7854 0 net88
rlabel metal1 9430 5134 9430 5134 0 net89
rlabel metal1 13570 1904 13570 1904 0 net9
rlabel metal2 7406 4828 7406 4828 0 net90
rlabel metal1 17894 2414 17894 2414 0 net91
rlabel metal1 14689 5678 14689 5678 0 net92
rlabel metal1 12006 1972 12006 1972 0 net93
rlabel metal2 13386 5882 13386 5882 0 net95
rlabel metal2 13662 10608 13662 10608 0 net98
rlabel metal1 7958 3026 7958 3026 0 net99
rlabel metal1 21206 3400 21206 3400 0 osc
rlabel metal1 18814 7480 18814 7480 0 resetb
rlabel metal2 23966 17340 23966 17340 0 ringosc.c\[0\]
rlabel metal2 18814 17850 18814 17850 0 ringosc.c\[1\]
rlabel metal1 16238 18156 16238 18156 0 ringosc.dstage\[0\].id.d0
rlabel metal1 16560 18326 16560 18326 0 ringosc.dstage\[0\].id.d1
rlabel metal1 16100 18258 16100 18258 0 ringosc.dstage\[0\].id.d2
rlabel metal1 22402 18088 22402 18088 0 ringosc.dstage\[0\].id.in
rlabel metal2 15318 17952 15318 17952 0 ringosc.dstage\[0\].id.out
rlabel metal1 17250 17680 17250 17680 0 ringosc.dstage\[0\].id.ts
rlabel metal2 23782 14110 23782 14110 0 ringosc.dstage\[10\].id.d0
rlabel metal1 23920 13974 23920 13974 0 ringosc.dstage\[10\].id.d1
rlabel metal2 23414 15300 23414 15300 0 ringosc.dstage\[10\].id.d2
rlabel metal2 22218 13668 22218 13668 0 ringosc.dstage\[10\].id.in
rlabel metal1 23598 14994 23598 14994 0 ringosc.dstage\[10\].id.out
rlabel metal2 22586 14178 22586 14178 0 ringosc.dstage\[10\].id.ts
rlabel metal1 23414 15980 23414 15980 0 ringosc.dstage\[11\].id.d0
rlabel metal2 23506 15810 23506 15810 0 ringosc.dstage\[11\].id.d1
rlabel metal1 23046 17238 23046 17238 0 ringosc.dstage\[11\].id.d2
rlabel metal2 23322 17170 23322 17170 0 ringosc.dstage\[11\].id.out
rlabel metal1 23414 16524 23414 16524 0 ringosc.dstage\[11\].id.ts
rlabel metal1 14858 16456 14858 16456 0 ringosc.dstage\[1\].id.d0
rlabel metal1 15456 17238 15456 17238 0 ringosc.dstage\[1\].id.d1
rlabel metal1 13938 16490 13938 16490 0 ringosc.dstage\[1\].id.d2
rlabel metal2 13570 17136 13570 17136 0 ringosc.dstage\[1\].id.out
rlabel metal2 14306 17646 14306 17646 0 ringosc.dstage\[1\].id.ts
rlabel metal1 12190 18156 12190 18156 0 ringosc.dstage\[2\].id.d0
rlabel metal2 12098 17680 12098 17680 0 ringosc.dstage\[2\].id.d1
rlabel metal1 11224 17238 11224 17238 0 ringosc.dstage\[2\].id.d2
rlabel metal1 12650 16558 12650 16558 0 ringosc.dstage\[2\].id.out
rlabel metal2 12742 17952 12742 17952 0 ringosc.dstage\[2\].id.ts
rlabel metal1 10350 16456 10350 16456 0 ringosc.dstage\[3\].id.d0
rlabel metal2 11086 16456 11086 16456 0 ringosc.dstage\[3\].id.d1
rlabel metal1 12098 15538 12098 15538 0 ringosc.dstage\[3\].id.d2
rlabel metal2 12926 15708 12926 15708 0 ringosc.dstage\[3\].id.out
rlabel metal2 12650 16286 12650 16286 0 ringosc.dstage\[3\].id.ts
rlabel metal1 19090 15674 19090 15674 0 ringosc.dstage\[4\].id.d0
rlabel metal1 18906 16184 18906 16184 0 ringosc.dstage\[4\].id.d1
rlabel metal1 18078 16150 18078 16150 0 ringosc.dstage\[4\].id.d2
rlabel metal1 18998 16082 18998 16082 0 ringosc.dstage\[4\].id.out
rlabel metal1 18216 15470 18216 15470 0 ringosc.dstage\[4\].id.ts
rlabel metal1 17664 16422 17664 16422 0 ringosc.dstage\[5\].id.d0
rlabel via1 18354 17306 18354 17306 0 ringosc.dstage\[5\].id.d1
rlabel metal1 20010 17102 20010 17102 0 ringosc.dstage\[5\].id.d2
rlabel metal2 18722 17748 18722 17748 0 ringosc.dstage\[5\].id.out
rlabel metal1 18224 16558 18224 16558 0 ringosc.dstage\[5\].id.ts
rlabel metal1 19412 14450 19412 14450 0 ringosc.dstage\[6\].id.d0
rlabel metal2 18538 13770 18538 13770 0 ringosc.dstage\[6\].id.d1
rlabel via2 18906 13243 18906 13243 0 ringosc.dstage\[6\].id.d2
rlabel metal1 20056 13974 20056 13974 0 ringosc.dstage\[6\].id.out
rlabel metal2 19642 16014 19642 16014 0 ringosc.dstage\[6\].id.ts
rlabel metal2 20102 13804 20102 13804 0 ringosc.dstage\[7\].id.d0
rlabel metal1 19872 11866 19872 11866 0 ringosc.dstage\[7\].id.d1
rlabel metal1 20470 11526 20470 11526 0 ringosc.dstage\[7\].id.d2
rlabel metal1 21298 12682 21298 12682 0 ringosc.dstage\[7\].id.out
rlabel metal1 20516 12818 20516 12818 0 ringosc.dstage\[7\].id.ts
rlabel metal1 23828 10778 23828 10778 0 ringosc.dstage\[8\].id.d0
rlabel metal1 23460 11050 23460 11050 0 ringosc.dstage\[8\].id.d1
rlabel metal1 23644 13294 23644 13294 0 ringosc.dstage\[8\].id.d2
rlabel metal1 23736 12342 23736 12342 0 ringosc.dstage\[8\].id.out
rlabel metal2 23874 12002 23874 12002 0 ringosc.dstage\[8\].id.ts
rlabel metal1 22954 11322 22954 11322 0 ringosc.dstage\[9\].id.d0
rlabel metal1 22356 12818 22356 12818 0 ringosc.dstage\[9\].id.d1
rlabel metal1 21298 13362 21298 13362 0 ringosc.dstage\[9\].id.d2
rlabel metal2 22862 13056 22862 13056 0 ringosc.dstage\[9\].id.ts
rlabel metal1 21896 17646 21896 17646 0 ringosc.iss.ctrl0
rlabel metal1 21482 14586 21482 14586 0 ringosc.iss.d0
rlabel metal1 22586 16150 22586 16150 0 ringosc.iss.d1
rlabel metal2 22494 18020 22494 18020 0 ringosc.iss.d2
rlabel metal2 20930 18292 20930 18292 0 ringosc.iss.one
<< properties >>
string FIXED_BBOX 0 0 26000 20000
<< end >>
