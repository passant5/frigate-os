VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO dll
  CLASS BLOCK ;
  FOREIGN dll ;
  ORIGIN 0.000 0.000 ;
  SIZE 130.000 BY 100.000 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 41.040 5.200 42.640 92.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 81.040 5.200 82.640 92.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 121.040 5.200 122.640 92.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 41.050 124.440 42.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 81.050 124.440 82.650 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 21.040 5.200 22.640 92.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 61.040 5.200 62.640 92.720 ;
    END
    PORT
      LAYER met2 ;
        RECT 101.040 5.200 102.640 92.720 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 21.050 124.440 22.650 ;
    END
    PORT
      LAYER met3 ;
        RECT 5.280 61.050 124.440 62.650 ;
    END
  END VPWR
  PIN clockp[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 58.050 96.000 58.330 100.000 ;
    END
  END clockp[0]
  PIN clockp[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.180800 ;
    PORT
      LAYER met2 ;
        RECT 70.930 96.000 71.210 100.000 ;
    END
  END clockp[1]
  PIN dco
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.424700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 101.750 0.000 102.030 4.000 ;
    END
  END dco
  PIN div[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END div[0]
  PIN div[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 17.110 0.000 17.390 4.000 ;
    END
  END div[1]
  PIN div[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 27.690 0.000 27.970 4.000 ;
    END
  END div[2]
  PIN div[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.270 0.000 38.550 4.000 ;
    END
  END div[3]
  PIN div[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.850 0.000 49.130 4.000 ;
    END
  END div[4]
  PIN div[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END div[5]
  PIN div[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.560700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END div[6]
  PIN div[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END div[7]
  PIN enable
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 91.170 0.000 91.450 4.000 ;
    END
  END enable
  PIN ext_trim[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 5.480 4.000 6.080 ;
    END
  END ext_trim[0]
  PIN ext_trim[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.410 96.000 19.690 100.000 ;
    END
  END ext_trim[10]
  PIN ext_trim[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 96.000 32.570 100.000 ;
    END
  END ext_trim[11]
  PIN ext_trim[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 96.000 45.450 100.000 ;
    END
  END ext_trim[12]
  PIN ext_trim[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 83.810 96.000 84.090 100.000 ;
    END
  END ext_trim[13]
  PIN ext_trim[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 96.690 96.000 96.970 100.000 ;
    END
  END ext_trim[14]
  PIN ext_trim[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 109.570 96.000 109.850 100.000 ;
    END
  END ext_trim[15]
  PIN ext_trim[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 122.450 96.000 122.730 100.000 ;
    END
  END ext_trim[16]
  PIN ext_trim[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 92.520 130.000 93.120 ;
    END
  END ext_trim[17]
  PIN ext_trim[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 81.640 130.000 82.240 ;
    END
  END ext_trim[18]
  PIN ext_trim[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 70.760 130.000 71.360 ;
    END
  END ext_trim[19]
  PIN ext_trim[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 16.360 4.000 16.960 ;
    END
  END ext_trim[1]
  PIN ext_trim[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 59.880 130.000 60.480 ;
    END
  END ext_trim[20]
  PIN ext_trim[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 49.000 130.000 49.600 ;
    END
  END ext_trim[21]
  PIN ext_trim[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 38.120 130.000 38.720 ;
    END
  END ext_trim[22]
  PIN ext_trim[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 27.240 130.000 27.840 ;
    END
  END ext_trim[23]
  PIN ext_trim[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 16.360 130.000 16.960 ;
    END
  END ext_trim[24]
  PIN ext_trim[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 126.000 5.480 130.000 6.080 ;
    END
  END ext_trim[25]
  PIN ext_trim[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END ext_trim[2]
  PIN ext_trim[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.120 4.000 38.720 ;
    END
  END ext_trim[3]
  PIN ext_trim[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END ext_trim[4]
  PIN ext_trim[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END ext_trim[5]
  PIN ext_trim[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END ext_trim[6]
  PIN ext_trim[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END ext_trim[7]
  PIN ext_trim[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END ext_trim[8]
  PIN ext_trim[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 6.530 96.000 6.810 100.000 ;
    END
  END ext_trim[9]
  PIN osc
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 122.910 0.000 123.190 4.000 ;
    END
  END osc
  PIN resetb
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END resetb
  OBS
      LAYER nwell ;
        RECT 5.330 5.355 124.390 92.565 ;
      LAYER li1 ;
        RECT 5.520 5.355 124.200 92.565 ;
      LAYER met1 ;
        RECT 5.520 3.440 125.510 96.520 ;
      LAYER met2 ;
        RECT 7.090 95.720 19.130 96.550 ;
        RECT 19.970 95.720 32.010 96.550 ;
        RECT 32.850 95.720 44.890 96.550 ;
        RECT 45.730 95.720 57.770 96.550 ;
        RECT 58.610 95.720 70.650 96.550 ;
        RECT 71.490 95.720 83.530 96.550 ;
        RECT 84.370 95.720 96.410 96.550 ;
        RECT 97.250 95.720 109.290 96.550 ;
        RECT 110.130 95.720 122.170 96.550 ;
        RECT 123.010 95.720 125.490 96.550 ;
        RECT 6.530 93.000 125.490 95.720 ;
        RECT 6.530 4.920 20.760 93.000 ;
        RECT 22.920 4.920 40.760 93.000 ;
        RECT 42.920 4.920 60.760 93.000 ;
        RECT 62.920 4.920 80.760 93.000 ;
        RECT 82.920 4.920 100.760 93.000 ;
        RECT 102.920 4.920 120.760 93.000 ;
        RECT 122.920 4.920 125.490 93.000 ;
        RECT 6.530 4.280 125.490 4.920 ;
        RECT 7.090 3.410 16.830 4.280 ;
        RECT 17.670 3.410 27.410 4.280 ;
        RECT 28.250 3.410 37.990 4.280 ;
        RECT 38.830 3.410 48.570 4.280 ;
        RECT 49.410 3.410 59.150 4.280 ;
        RECT 59.990 3.410 69.730 4.280 ;
        RECT 70.570 3.410 80.310 4.280 ;
        RECT 81.150 3.410 90.890 4.280 ;
        RECT 91.730 3.410 101.470 4.280 ;
        RECT 102.310 3.410 112.050 4.280 ;
        RECT 112.890 3.410 122.630 4.280 ;
        RECT 123.470 3.410 125.490 4.280 ;
      LAYER met3 ;
        RECT 4.400 92.120 125.600 92.985 ;
        RECT 3.990 83.050 126.000 92.120 ;
        RECT 3.990 82.640 4.880 83.050 ;
        RECT 4.400 81.240 4.880 82.640 ;
        RECT 3.990 80.650 4.880 81.240 ;
        RECT 124.840 82.640 126.000 83.050 ;
        RECT 124.840 81.240 125.600 82.640 ;
        RECT 124.840 80.650 126.000 81.240 ;
        RECT 3.990 71.760 126.000 80.650 ;
        RECT 4.400 70.360 125.600 71.760 ;
        RECT 3.990 63.050 126.000 70.360 ;
        RECT 3.990 60.880 4.880 63.050 ;
        RECT 4.400 60.650 4.880 60.880 ;
        RECT 124.840 60.880 126.000 63.050 ;
        RECT 124.840 60.650 125.600 60.880 ;
        RECT 4.400 59.480 125.600 60.650 ;
        RECT 3.990 50.000 126.000 59.480 ;
        RECT 4.400 48.600 125.600 50.000 ;
        RECT 3.990 43.050 126.000 48.600 ;
        RECT 3.990 40.650 4.880 43.050 ;
        RECT 124.840 40.650 126.000 43.050 ;
        RECT 3.990 39.120 126.000 40.650 ;
        RECT 4.400 37.720 125.600 39.120 ;
        RECT 3.990 28.240 126.000 37.720 ;
        RECT 4.400 26.840 125.600 28.240 ;
        RECT 3.990 23.050 126.000 26.840 ;
        RECT 3.990 20.650 4.880 23.050 ;
        RECT 124.840 20.650 126.000 23.050 ;
        RECT 3.990 17.360 126.000 20.650 ;
        RECT 4.400 15.960 125.600 17.360 ;
        RECT 3.990 6.480 126.000 15.960 ;
        RECT 4.400 5.615 125.600 6.480 ;
  END
END dll
END LIBRARY

