module analog_ctrl_regs_APB (IRQ,
    PCLK,
    PENABLE,
    PREADY,
    PRESETn,
    PSEL,
    PWRITE,
    adc0_to_analog1,
    adc0_to_dac0,
    adc0_to_left_vref,
    adc0_to_tempsense,
    adc0_to_vbgtc,
    adc0_to_voutref,
    adc1_to_analog0,
    adc1_to_dac1,
    adc1_to_right_vref,
    adc1_to_vbgsc,
    adc1_to_vinref,
    bandgap_ena,
    bandgap_sel,
    brownout_ena,
    brownout_filt,
    brownout_isrc_sel,
    brownout_oneshot,
    brownout_rc_dis,
    brownout_rc_ena,
    brownout_timeout,
    brownout_unfilt,
    brownout_vunder,
    comp_ena,
    comp_n_to_analog0,
    comp_n_to_dac1,
    comp_n_to_right_vref,
    comp_n_to_sio1,
    comp_n_to_vbgsc,
    comp_n_to_vinref,
    comp_out,
    comp_p_to_analog1,
    comp_p_to_dac0,
    comp_p_to_left_vref,
    comp_p_to_sio0,
    comp_p_to_tempsense,
    comp_p_to_vbgtc,
    comp_p_to_voutref,
    dac0_to_analog1,
    dac0_to_user,
    dac1_to_analog0,
    dac1_to_user,
    ibias_ena,
    ibias_ref_select,
    idac_ena,
    ldo_ena,
    ldo_ref_sel,
    left_hgbw_opamp_ena,
    left_hgbw_opamp_n_to_amuxbusB,
    left_hgbw_opamp_n_to_analog1,
    left_hgbw_opamp_n_to_dac1,
    left_hgbw_opamp_n_to_rheostat_out,
    left_hgbw_opamp_n_to_rheostat_tap,
    left_hgbw_opamp_n_to_right_vref,
    left_hgbw_opamp_n_to_sio1,
    left_hgbw_opamp_n_to_vbgtc,
    left_hgbw_opamp_n_to_vinref,
    left_hgbw_opamp_p_to_amuxbusA,
    left_hgbw_opamp_p_to_analog0,
    left_hgbw_opamp_p_to_dac0,
    left_hgbw_opamp_p_to_left_vref,
    left_hgbw_opamp_p_to_rheostat_out,
    left_hgbw_opamp_p_to_sio0,
    left_hgbw_opamp_p_to_tempsense,
    left_hgbw_opamp_p_to_voutref,
    left_instramp_ena,
    left_instramp_n_to_amuxbusB,
    left_instramp_n_to_analog1,
    left_instramp_n_to_right_vref,
    left_instramp_n_to_sio1,
    left_instramp_n_to_vinref,
    left_instramp_p_to_amuxbusA,
    left_instramp_p_to_analog0,
    left_instramp_p_to_left_vref,
    left_instramp_p_to_sio0,
    left_instramp_p_to_tempsense,
    left_instramp_p_to_voutref,
    left_lp_opamp_ena,
    left_lp_opamp_n_to_amuxbusB,
    left_lp_opamp_n_to_analog1,
    left_lp_opamp_n_to_dac1,
    left_lp_opamp_n_to_rheostat_out,
    left_lp_opamp_n_to_rheostat_tap,
    left_lp_opamp_n_to_right_vref,
    left_lp_opamp_n_to_sio1,
    left_lp_opamp_n_to_vbgsc,
    left_lp_opamp_n_to_vinref,
    left_lp_opamp_p_to_amuxbusA,
    left_lp_opamp_p_to_analog0,
    left_lp_opamp_p_to_dac0,
    left_lp_opamp_p_to_left_vref,
    left_lp_opamp_p_to_rheostat_out,
    left_lp_opamp_p_to_sio0,
    left_lp_opamp_p_to_voutref,
    left_vref_to_user,
    overvoltage_ena,
    overvoltage_out,
    rdac0_ena,
    rdac1_ena,
    right_hgbw_opamp_ena,
    right_hgbw_opamp_n_to_amuxbusB,
    right_hgbw_opamp_n_to_analog1,
    right_hgbw_opamp_n_to_dac1,
    right_hgbw_opamp_n_to_rheostat_out,
    right_hgbw_opamp_n_to_rheostat_tap,
    right_hgbw_opamp_n_to_right_vref,
    right_hgbw_opamp_n_to_sio1,
    right_hgbw_opamp_n_to_vbgsc,
    right_hgbw_opamp_n_to_vinref,
    right_hgbw_opamp_p_to_amuxbusA,
    right_hgbw_opamp_p_to_analog0,
    right_hgbw_opamp_p_to_dac0,
    right_hgbw_opamp_p_to_left_vref,
    right_hgbw_opamp_p_to_rheostat_out,
    right_hgbw_opamp_p_to_sio0,
    right_hgbw_opamp_p_to_voutref,
    right_instramp_ena,
    right_instramp_n_to_amuxbusB,
    right_instramp_n_to_analog1,
    right_instramp_n_to_right_vref,
    right_instramp_n_to_sio1,
    right_instramp_n_to_vinref,
    right_instramp_p_to_amuxbusA,
    right_instramp_p_to_analog0,
    right_instramp_p_to_left_vref,
    right_instramp_p_to_sio0,
    right_instramp_p_to_tempsense,
    right_instramp_p_to_voutref,
    right_lp_opamp_ena,
    right_lp_opamp_n_to_amuxbusB,
    right_lp_opamp_n_to_analog1,
    right_lp_opamp_n_to_dac1,
    right_lp_opamp_n_to_rheostat_out,
    right_lp_opamp_n_to_rheostat_tap,
    right_lp_opamp_n_to_right_vref,
    right_lp_opamp_n_to_sio1,
    right_lp_opamp_n_to_vbgtc,
    right_lp_opamp_n_to_vinref,
    right_lp_opamp_p_to_amuxbusA,
    right_lp_opamp_p_to_analog0,
    right_lp_opamp_p_to_dac0,
    right_lp_opamp_p_to_left_vref,
    right_lp_opamp_p_to_rheostat_out,
    right_lp_opamp_p_to_sio0,
    right_lp_opamp_p_to_tempsense,
    right_lp_opamp_p_to_voutref,
    right_vref_to_user,
    tempsense_ena,
    tempsense_sel,
    tempsense_to_user,
    ulpcomp_clk,
    ulpcomp_ena,
    ulpcomp_n_to_analog0,
    ulpcomp_n_to_dac1,
    ulpcomp_n_to_right_vref,
    ulpcomp_n_to_sio1,
    ulpcomp_n_to_vbgsc,
    ulpcomp_n_to_vinref,
    ulpcomp_out,
    ulpcomp_p_to_analog1,
    ulpcomp_p_to_dac0,
    ulpcomp_p_to_left_vref,
    ulpcomp_p_to_sio0,
    ulpcomp_p_to_tempsense,
    ulpcomp_p_to_vbgtc,
    ulpcomp_p_to_voutref,
    vbgsc_to_user,
    vbgtc_to_user,
    vccd1_pwr_good,
    vccd2_pwr_good,
    vdda1_pwr_good,
    vdda2_pwr_good,
    vinref_to_user,
    voutref_to_user,
    vccd0,
    vssd0,
    PADDR,
    PRDATA,
    PWDATA,
    adc0_to_gpio1_3,
    adc0_to_gpio6_4,
    adc1_to_gpio1_2,
    adc1_to_gpio6_5,
    adc_refh_to_gpio6_6,
    adc_refl_to_gpio6_7,
    analog0_connect,
    analog1_connect,
    audiodac_out_to_analog1,
    audiodac_outb_to_analog0,
    bandgap_trim,
    brownout_otrip,
    brownout_vtrip,
    comp_hyst,
    comp_n_to_gpio1_4,
    comp_n_to_gpio6_3,
    comp_p_to_gpio1_5,
    comp_p_to_gpio6_2,
    comp_trim,
    dac_refh_to_gpio1_1,
    dac_refl_to_gpio1_0,
    ibias_snk_ena,
    ibias_src_ena,
    ibias_test_to_gpio1_2,
    idac_to_gpio1_2,
    idac_to_gpio1_3,
    idac_value,
    left_hgbw_opamp_n_to_gpio2_0,
    left_hgbw_opamp_n_to_gpio5_3,
    left_hgbw_opamp_p_to_gpio2_1,
    left_hgbw_opamp_p_to_gpio5_2,
    left_hgbw_opamp_to_adc0,
    left_hgbw_opamp_to_amuxbusB,
    left_hgbw_opamp_to_analog1,
    left_hgbw_opamp_to_comp_p,
    left_hgbw_opamp_to_gpio3_1,
    left_hgbw_opamp_to_gpio3_5,
    left_hgbw_opamp_to_gpio4_1,
    left_hgbw_opamp_to_gpio4_5,
    left_hgbw_opamp_to_ulpcomp_p,
    left_instramp_G1,
    left_instramp_G2,
    left_instramp_n_to_gpio5_7,
    left_instramp_p_to_gpio5_6,
    left_instramp_to_adc0,
    left_instramp_to_amuxbusB,
    left_instramp_to_analog1,
    left_instramp_to_comp_p,
    left_instramp_to_gpio4_4,
    left_instramp_to_ulpcomp_p,
    left_lp_opamp_n_to_gpio5_5,
    left_lp_opamp_p_to_gpio5_4,
    left_lp_opamp_to_adc1,
    left_lp_opamp_to_amuxbusA,
    left_lp_opamp_to_analog0,
    left_lp_opamp_to_comp_n,
    left_lp_opamp_to_gpio3_4,
    left_lp_opamp_to_gpio4_0,
    left_lp_opamp_to_ulpcomp_n,
    left_rheostat1_b,
    left_rheostat2_b,
    overvoltage_trim,
    rdac0_value,
    rdac1_value,
    right_hgbw_opamp_n_to_gpio2_2,
    right_hgbw_opamp_n_to_gpio5_1,
    right_hgbw_opamp_p_to_gpio2_3,
    right_hgbw_opamp_p_to_gpio5_0,
    right_hgbw_opamp_to_adc1,
    right_hgbw_opamp_to_amuxbusA,
    right_hgbw_opamp_to_analog0,
    right_hgbw_opamp_to_comp_n,
    right_hgbw_opamp_to_gpio3_2,
    right_hgbw_opamp_to_gpio3_6,
    right_hgbw_opamp_to_gpio4_2,
    right_hgbw_opamp_to_gpio4_6,
    right_hgbw_opamp_to_ulpcomp_n,
    right_instramp_G1,
    right_instramp_G2,
    right_instramp_n_to_gpio2_6,
    right_instramp_p_to_gpio2_7,
    right_instramp_to_adc1,
    right_instramp_to_amuxbusA,
    right_instramp_to_analog0,
    right_instramp_to_comp_n,
    right_instramp_to_gpio3_0,
    right_instramp_to_ulpcomp_n,
    right_lp_opamp_n_to_gpio2_4,
    right_lp_opamp_p_to_gpio2_5,
    right_lp_opamp_to_adc0,
    right_lp_opamp_to_amuxbusB,
    right_lp_opamp_to_analog1,
    right_lp_opamp_to_comp_p,
    right_lp_opamp_to_gpio3_3,
    right_lp_opamp_to_gpio3_7,
    right_lp_opamp_to_gpio4_3,
    right_lp_opamp_to_gpio4_7,
    right_lp_opamp_to_ulpcomp_p,
    right_rheostat1_b,
    right_rheostat2_b,
    sio0_connect,
    sio1_connect,
    ulpcomp_n_to_gpio1_6,
    ulpcomp_n_to_gpio6_1,
    ulpcomp_p_to_gpio1_7,
    ulpcomp_p_to_gpio6_0,
    user_to_adc0,
    user_to_adc1,
    user_to_comp_n,
    user_to_comp_p,
    user_to_ulpcomp_n,
    user_to_ulpcomp_p,
    vbg_test_to_gpio1_1);
 output IRQ;
 input PCLK;
 input PENABLE;
 output PREADY;
 input PRESETn;
 input PSEL;
 input PWRITE;
 output adc0_to_analog1;
 output adc0_to_dac0;
 output adc0_to_left_vref;
 output adc0_to_tempsense;
 output adc0_to_vbgtc;
 output adc0_to_voutref;
 output adc1_to_analog0;
 output adc1_to_dac1;
 output adc1_to_right_vref;
 output adc1_to_vbgsc;
 output adc1_to_vinref;
 output bandgap_ena;
 output bandgap_sel;
 output brownout_ena;
 input brownout_filt;
 output brownout_isrc_sel;
 output brownout_oneshot;
 output brownout_rc_dis;
 output brownout_rc_ena;
 input brownout_timeout;
 input brownout_unfilt;
 input brownout_vunder;
 output comp_ena;
 output comp_n_to_analog0;
 output comp_n_to_dac1;
 output comp_n_to_right_vref;
 output comp_n_to_sio1;
 output comp_n_to_vbgsc;
 output comp_n_to_vinref;
 input comp_out;
 output comp_p_to_analog1;
 output comp_p_to_dac0;
 output comp_p_to_left_vref;
 output comp_p_to_sio0;
 output comp_p_to_tempsense;
 output comp_p_to_vbgtc;
 output comp_p_to_voutref;
 output dac0_to_analog1;
 output dac0_to_user;
 output dac1_to_analog0;
 output dac1_to_user;
 output ibias_ena;
 output ibias_ref_select;
 output idac_ena;
 output ldo_ena;
 output ldo_ref_sel;
 output left_hgbw_opamp_ena;
 output left_hgbw_opamp_n_to_amuxbusB;
 output left_hgbw_opamp_n_to_analog1;
 output left_hgbw_opamp_n_to_dac1;
 output left_hgbw_opamp_n_to_rheostat_out;
 output left_hgbw_opamp_n_to_rheostat_tap;
 output left_hgbw_opamp_n_to_right_vref;
 output left_hgbw_opamp_n_to_sio1;
 output left_hgbw_opamp_n_to_vbgtc;
 output left_hgbw_opamp_n_to_vinref;
 output left_hgbw_opamp_p_to_amuxbusA;
 output left_hgbw_opamp_p_to_analog0;
 output left_hgbw_opamp_p_to_dac0;
 output left_hgbw_opamp_p_to_left_vref;
 output left_hgbw_opamp_p_to_rheostat_out;
 output left_hgbw_opamp_p_to_sio0;
 output left_hgbw_opamp_p_to_tempsense;
 output left_hgbw_opamp_p_to_voutref;
 output left_instramp_ena;
 output left_instramp_n_to_amuxbusB;
 output left_instramp_n_to_analog1;
 output left_instramp_n_to_right_vref;
 output left_instramp_n_to_sio1;
 output left_instramp_n_to_vinref;
 output left_instramp_p_to_amuxbusA;
 output left_instramp_p_to_analog0;
 output left_instramp_p_to_left_vref;
 output left_instramp_p_to_sio0;
 output left_instramp_p_to_tempsense;
 output left_instramp_p_to_voutref;
 output left_lp_opamp_ena;
 output left_lp_opamp_n_to_amuxbusB;
 output left_lp_opamp_n_to_analog1;
 output left_lp_opamp_n_to_dac1;
 output left_lp_opamp_n_to_rheostat_out;
 output left_lp_opamp_n_to_rheostat_tap;
 output left_lp_opamp_n_to_right_vref;
 output left_lp_opamp_n_to_sio1;
 output left_lp_opamp_n_to_vbgsc;
 output left_lp_opamp_n_to_vinref;
 output left_lp_opamp_p_to_amuxbusA;
 output left_lp_opamp_p_to_analog0;
 output left_lp_opamp_p_to_dac0;
 output left_lp_opamp_p_to_left_vref;
 output left_lp_opamp_p_to_rheostat_out;
 output left_lp_opamp_p_to_sio0;
 output left_lp_opamp_p_to_voutref;
 output left_vref_to_user;
 output overvoltage_ena;
 input overvoltage_out;
 output rdac0_ena;
 output rdac1_ena;
 output right_hgbw_opamp_ena;
 output right_hgbw_opamp_n_to_amuxbusB;
 output right_hgbw_opamp_n_to_analog1;
 output right_hgbw_opamp_n_to_dac1;
 output right_hgbw_opamp_n_to_rheostat_out;
 output right_hgbw_opamp_n_to_rheostat_tap;
 output right_hgbw_opamp_n_to_right_vref;
 output right_hgbw_opamp_n_to_sio1;
 output right_hgbw_opamp_n_to_vbgsc;
 output right_hgbw_opamp_n_to_vinref;
 output right_hgbw_opamp_p_to_amuxbusA;
 output right_hgbw_opamp_p_to_analog0;
 output right_hgbw_opamp_p_to_dac0;
 output right_hgbw_opamp_p_to_left_vref;
 output right_hgbw_opamp_p_to_rheostat_out;
 output right_hgbw_opamp_p_to_sio0;
 output right_hgbw_opamp_p_to_voutref;
 output right_instramp_ena;
 output right_instramp_n_to_amuxbusB;
 output right_instramp_n_to_analog1;
 output right_instramp_n_to_right_vref;
 output right_instramp_n_to_sio1;
 output right_instramp_n_to_vinref;
 output right_instramp_p_to_amuxbusA;
 output right_instramp_p_to_analog0;
 output right_instramp_p_to_left_vref;
 output right_instramp_p_to_sio0;
 output right_instramp_p_to_tempsense;
 output right_instramp_p_to_voutref;
 output right_lp_opamp_ena;
 output right_lp_opamp_n_to_amuxbusB;
 output right_lp_opamp_n_to_analog1;
 output right_lp_opamp_n_to_dac1;
 output right_lp_opamp_n_to_rheostat_out;
 output right_lp_opamp_n_to_rheostat_tap;
 output right_lp_opamp_n_to_right_vref;
 output right_lp_opamp_n_to_sio1;
 output right_lp_opamp_n_to_vbgtc;
 output right_lp_opamp_n_to_vinref;
 output right_lp_opamp_p_to_amuxbusA;
 output right_lp_opamp_p_to_analog0;
 output right_lp_opamp_p_to_dac0;
 output right_lp_opamp_p_to_left_vref;
 output right_lp_opamp_p_to_rheostat_out;
 output right_lp_opamp_p_to_sio0;
 output right_lp_opamp_p_to_tempsense;
 output right_lp_opamp_p_to_voutref;
 output right_vref_to_user;
 output tempsense_ena;
 output tempsense_sel;
 output tempsense_to_user;
 output ulpcomp_clk;
 output ulpcomp_ena;
 output ulpcomp_n_to_analog0;
 output ulpcomp_n_to_dac1;
 output ulpcomp_n_to_right_vref;
 output ulpcomp_n_to_sio1;
 output ulpcomp_n_to_vbgsc;
 output ulpcomp_n_to_vinref;
 input ulpcomp_out;
 output ulpcomp_p_to_analog1;
 output ulpcomp_p_to_dac0;
 output ulpcomp_p_to_left_vref;
 output ulpcomp_p_to_sio0;
 output ulpcomp_p_to_tempsense;
 output ulpcomp_p_to_vbgtc;
 output ulpcomp_p_to_voutref;
 output vbgsc_to_user;
 output vbgtc_to_user;
 input vccd1_pwr_good;
 input vccd2_pwr_good;
 input vdda1_pwr_good;
 input vdda2_pwr_good;
 output vinref_to_user;
 output voutref_to_user;
 inout vccd0;
 inout vssd0;
 input [31:0] PADDR;
 output [31:0] PRDATA;
 input [31:0] PWDATA;
 output [1:0] adc0_to_gpio1_3;
 output [1:0] adc0_to_gpio6_4;
 output [1:0] adc1_to_gpio1_2;
 output [1:0] adc1_to_gpio6_5;
 output [1:0] adc_refh_to_gpio6_6;
 output [1:0] adc_refl_to_gpio6_7;
 output [1:0] analog0_connect;
 output [1:0] analog1_connect;
 output [1:0] audiodac_out_to_analog1;
 output [1:0] audiodac_outb_to_analog0;
 output [15:0] bandgap_trim;
 output [2:0] brownout_otrip;
 output [2:0] brownout_vtrip;
 output [1:0] comp_hyst;
 output [1:0] comp_n_to_gpio1_4;
 output [1:0] comp_n_to_gpio6_3;
 output [1:0] comp_p_to_gpio1_5;
 output [1:0] comp_p_to_gpio6_2;
 output [5:0] comp_trim;
 output [1:0] dac_refh_to_gpio1_1;
 output [1:0] dac_refl_to_gpio1_0;
 output [3:0] ibias_snk_ena;
 output [23:0] ibias_src_ena;
 output [1:0] ibias_test_to_gpio1_2;
 output [1:0] idac_to_gpio1_2;
 output [1:0] idac_to_gpio1_3;
 output [11:0] idac_value;
 output [1:0] left_hgbw_opamp_n_to_gpio2_0;
 output [1:0] left_hgbw_opamp_n_to_gpio5_3;
 output [1:0] left_hgbw_opamp_p_to_gpio2_1;
 output [1:0] left_hgbw_opamp_p_to_gpio5_2;
 output [1:0] left_hgbw_opamp_to_adc0;
 output [1:0] left_hgbw_opamp_to_amuxbusB;
 output [1:0] left_hgbw_opamp_to_analog1;
 output [1:0] left_hgbw_opamp_to_comp_p;
 output [1:0] left_hgbw_opamp_to_gpio3_1;
 output [1:0] left_hgbw_opamp_to_gpio3_5;
 output [1:0] left_hgbw_opamp_to_gpio4_1;
 output [1:0] left_hgbw_opamp_to_gpio4_5;
 output [1:0] left_hgbw_opamp_to_ulpcomp_p;
 output [4:0] left_instramp_G1;
 output [4:0] left_instramp_G2;
 output [1:0] left_instramp_n_to_gpio5_7;
 output [1:0] left_instramp_p_to_gpio5_6;
 output [1:0] left_instramp_to_adc0;
 output [1:0] left_instramp_to_amuxbusB;
 output [1:0] left_instramp_to_analog1;
 output [1:0] left_instramp_to_comp_p;
 output [1:0] left_instramp_to_gpio4_4;
 output [1:0] left_instramp_to_ulpcomp_p;
 output [1:0] left_lp_opamp_n_to_gpio5_5;
 output [1:0] left_lp_opamp_p_to_gpio5_4;
 output [1:0] left_lp_opamp_to_adc1;
 output [1:0] left_lp_opamp_to_amuxbusA;
 output [1:0] left_lp_opamp_to_analog0;
 output [1:0] left_lp_opamp_to_comp_n;
 output [1:0] left_lp_opamp_to_gpio3_4;
 output [1:0] left_lp_opamp_to_gpio4_0;
 output [1:0] left_lp_opamp_to_ulpcomp_n;
 output [7:0] left_rheostat1_b;
 output [7:0] left_rheostat2_b;
 output [3:0] overvoltage_trim;
 output [11:0] rdac0_value;
 output [11:0] rdac1_value;
 output [1:0] right_hgbw_opamp_n_to_gpio2_2;
 output [1:0] right_hgbw_opamp_n_to_gpio5_1;
 output [1:0] right_hgbw_opamp_p_to_gpio2_3;
 output [1:0] right_hgbw_opamp_p_to_gpio5_0;
 output [1:0] right_hgbw_opamp_to_adc1;
 output [1:0] right_hgbw_opamp_to_amuxbusA;
 output [1:0] right_hgbw_opamp_to_analog0;
 output [1:0] right_hgbw_opamp_to_comp_n;
 output [1:0] right_hgbw_opamp_to_gpio3_2;
 output [1:0] right_hgbw_opamp_to_gpio3_6;
 output [1:0] right_hgbw_opamp_to_gpio4_2;
 output [1:0] right_hgbw_opamp_to_gpio4_6;
 output [1:0] right_hgbw_opamp_to_ulpcomp_n;
 output [4:0] right_instramp_G1;
 output [4:0] right_instramp_G2;
 output [1:0] right_instramp_n_to_gpio2_6;
 output [1:0] right_instramp_p_to_gpio2_7;
 output [1:0] right_instramp_to_adc1;
 output [1:0] right_instramp_to_amuxbusA;
 output [1:0] right_instramp_to_analog0;
 output [1:0] right_instramp_to_comp_n;
 output [1:0] right_instramp_to_gpio3_0;
 output [1:0] right_instramp_to_ulpcomp_n;
 output [1:0] right_lp_opamp_n_to_gpio2_4;
 output [1:0] right_lp_opamp_p_to_gpio2_5;
 output [1:0] right_lp_opamp_to_adc0;
 output [1:0] right_lp_opamp_to_amuxbusB;
 output [1:0] right_lp_opamp_to_analog1;
 output [1:0] right_lp_opamp_to_comp_p;
 output [1:0] right_lp_opamp_to_gpio3_3;
 output [1:0] right_lp_opamp_to_gpio3_7;
 output [1:0] right_lp_opamp_to_gpio4_3;
 output [1:0] right_lp_opamp_to_gpio4_7;
 output [1:0] right_lp_opamp_to_ulpcomp_p;
 output [7:0] right_rheostat1_b;
 output [7:0] right_rheostat2_b;
 output [1:0] sio0_connect;
 output [1:0] sio1_connect;
 output [1:0] ulpcomp_n_to_gpio1_6;
 output [1:0] ulpcomp_n_to_gpio6_1;
 output [1:0] ulpcomp_p_to_gpio1_7;
 output [1:0] ulpcomp_p_to_gpio6_0;
 output [1:0] user_to_adc0;
 output [1:0] user_to_adc1;
 output [1:0] user_to_comp_n;
 output [1:0] user_to_comp_p;
 output [1:0] user_to_ulpcomp_n;
 output [1:0] user_to_ulpcomp_p;
 output [1:0] vbg_test_to_gpio1_1;

 wire n1000;
 wire n1001;
 wire n1002;
 wire n1003;
 wire n1004;
 wire n1005;
 wire n1006;
 wire n1007;
 wire n1008;
 wire n1009;
 wire n1010;
 wire n1011;
 wire n1012;
 wire n1013;
 wire n1015;
 wire n1016;
 wire n1017;
 wire n1018;
 wire n1019;
 wire n1020;
 wire n1021;
 wire n1022;
 wire n1023;
 wire n1024;
 wire n1025;
 wire n1026;
 wire n1027;
 wire n1028;
 wire n1029;
 wire n1030;
 wire n1031;
 wire n1032;
 wire n1033;
 wire n1034;
 wire n1035;
 wire n1036;
 wire n1037;
 wire n1038;
 wire n1039;
 wire n1040;
 wire n1041;
 wire n1042;
 wire n1043;
 wire n1044;
 wire n1045;
 wire n1046;
 wire n1048;
 wire n1049;
 wire n1051;
 wire n1052;
 wire n1053;
 wire n1054;
 wire n1055;
 wire n1056;
 wire n1057;
 wire n1058;
 wire n1059;
 wire n1060;
 wire n1061;
 wire n1062;
 wire n1063;
 wire n1064;
 wire n1065;
 wire n1066;
 wire n1067;
 wire n1068;
 wire n1069;
 wire n1070;
 wire n1071;
 wire n1072;
 wire n1073;
 wire n1074;
 wire n1075;
 wire n1076;
 wire n1077;
 wire n1078;
 wire n1079;
 wire n1080;
 wire n1081;
 wire n1082;
 wire n1083;
 wire n1084;
 wire n1085;
 wire n1086;
 wire n1087;
 wire n1088;
 wire n1089;
 wire n1090;
 wire n1091;
 wire n1092;
 wire n1093;
 wire n1094;
 wire n1095;
 wire n1096;
 wire n1097;
 wire n1098;
 wire n1099;
 wire n1100;
 wire n1101;
 wire n1102;
 wire n1103;
 wire n1104;
 wire n1105;
 wire n1106;
 wire n1107;
 wire n1108;
 wire n1109;
 wire n1110;
 wire n1111;
 wire n1112;
 wire n1113;
 wire n1114;
 wire n1115;
 wire n1116;
 wire n1117;
 wire n1118;
 wire n1119;
 wire n1120;
 wire n1121;
 wire n1122;
 wire n1123;
 wire n1124;
 wire n1125;
 wire n1126;
 wire n1127;
 wire n1129;
 wire n1130;
 wire n1131;
 wire n1132;
 wire n1133;
 wire n1134;
 wire n1135;
 wire n1136;
 wire n1137;
 wire n1138;
 wire n1139;
 wire n1140;
 wire n1141;
 wire n1142;
 wire n1146;
 wire n1147;
 wire n1148;
 wire n1149;
 wire n1150;
 wire n1151;
 wire n1152;
 wire n1153;
 wire n1154;
 wire n1155;
 wire n1156;
 wire n1157;
 wire n1158;
 wire n1159;
 wire n1160;
 wire n1161;
 wire n1162;
 wire n1163;
 wire n1164;
 wire n1165;
 wire n1166;
 wire n1167;
 wire n1168;
 wire n1169;
 wire n1170;
 wire n1171;
 wire n1172;
 wire n1173;
 wire n1174;
 wire n1175;
 wire n1176;
 wire n1177;
 wire n1178;
 wire n1179;
 wire n1180;
 wire n1181;
 wire n1182;
 wire n1183;
 wire n1184;
 wire n1185;
 wire n1186;
 wire n1187;
 wire n1188;
 wire n1189;
 wire n1190;
 wire n1191;
 wire n1192;
 wire n1193;
 wire n1194;
 wire n1195;
 wire n1197;
 wire n1198;
 wire n1199;
 wire n1200;
 wire n1201;
 wire n1202;
 wire n1203;
 wire n1204;
 wire n1205;
 wire n1206;
 wire n1207;
 wire n1208;
 wire n1209;
 wire n1210;
 wire n1211;
 wire n1212;
 wire n1213;
 wire n1214;
 wire n1215;
 wire n1216;
 wire n1217;
 wire n1218;
 wire n1219;
 wire n1220;
 wire n1221;
 wire n1222;
 wire n1223;
 wire n1224;
 wire n1225;
 wire n1228;
 wire n1229;
 wire n1230;
 wire n1231;
 wire n1232;
 wire n1233;
 wire n1234;
 wire n1235;
 wire n1236;
 wire n1237;
 wire n1238;
 wire n1239;
 wire n1240;
 wire n1241;
 wire n1242;
 wire n1243;
 wire n1244;
 wire n1245;
 wire n1246;
 wire n1247;
 wire n1248;
 wire n1249;
 wire n1250;
 wire n1251;
 wire n1252;
 wire n1253;
 wire n1254;
 wire n1255;
 wire n1256;
 wire n1260;
 wire n1261;
 wire n1262;
 wire n1263;
 wire n1264;
 wire n1265;
 wire n1266;
 wire n1267;
 wire n1268;
 wire n1269;
 wire n1270;
 wire n1271;
 wire n1272;
 wire n1273;
 wire n1274;
 wire n1275;
 wire n1276;
 wire n1277;
 wire n1278;
 wire n1280;
 wire n1281;
 wire n1282;
 wire n1283;
 wire n1284;
 wire n1285;
 wire n1287;
 wire n1288;
 wire n1290;
 wire n1291;
 wire n1292;
 wire n1294;
 wire n1295;
 wire n1296;
 wire n1297;
 wire n1298;
 wire n1299;
 wire n1300;
 wire n1301;
 wire n1302;
 wire n1303;
 wire n1304;
 wire n1305;
 wire n1306;
 wire n1307;
 wire n1308;
 wire n1309;
 wire n1310;
 wire n1311;
 wire n1312;
 wire n1313;
 wire n1314;
 wire n1315;
 wire n1316;
 wire n1317;
 wire n1318;
 wire n1319;
 wire n1320;
 wire n1321;
 wire n1322;
 wire n1323;
 wire n1324;
 wire n1325;
 wire n1326;
 wire n1327;
 wire n1328;
 wire n1329;
 wire n1330;
 wire n1331;
 wire n1332;
 wire n1333;
 wire n1336;
 wire n1337;
 wire n1338;
 wire n1339;
 wire n1340;
 wire n1341;
 wire n1342;
 wire n1343;
 wire n1344;
 wire n1345;
 wire n1346;
 wire n1347;
 wire n1348;
 wire n1349;
 wire n1350;
 wire n1351;
 wire n1352;
 wire n1353;
 wire n1354;
 wire n1355;
 wire n1356;
 wire n1357;
 wire n1358;
 wire n1359;
 wire n1360;
 wire n1361;
 wire n1362;
 wire n1363;
 wire n1366;
 wire n1367;
 wire n1368;
 wire n1369;
 wire n1370;
 wire n1371;
 wire n1372;
 wire n1373;
 wire n1374;
 wire n1375;
 wire n1376;
 wire n1377;
 wire n1378;
 wire n1379;
 wire n1380;
 wire n1381;
 wire n1382;
 wire n1383;
 wire n1384;
 wire n1385;
 wire n1386;
 wire n1387;
 wire n1388;
 wire n1389;
 wire n1390;
 wire n1391;
 wire n1392;
 wire n1393;
 wire n1394;
 wire n1395;
 wire n1396;
 wire n1397;
 wire n1398;
 wire n1399;
 wire n1400;
 wire n1401;
 wire n1402;
 wire n1403;
 wire n1404;
 wire n1405;
 wire n1406;
 wire n1407;
 wire n1408;
 wire n1409;
 wire n1410;
 wire n1411;
 wire n1412;
 wire n1413;
 wire n1414;
 wire n1415;
 wire n1416;
 wire n1417;
 wire n1418;
 wire n1419;
 wire n1420;
 wire n1421;
 wire n1422;
 wire n1423;
 wire n1424;
 wire n1425;
 wire n1426;
 wire n1427;
 wire n1428;
 wire n1429;
 wire n1430;
 wire n1431;
 wire n1432;
 wire n1433;
 wire n1434;
 wire n1435;
 wire n1436;
 wire n1437;
 wire n1438;
 wire n1439;
 wire n1440;
 wire n1441;
 wire n1442;
 wire n1443;
 wire n1444;
 wire n1445;
 wire n1446;
 wire n1447;
 wire n1448;
 wire n1449;
 wire n1450;
 wire n1451;
 wire n1452;
 wire n1453;
 wire n1454;
 wire n1455;
 wire n1456;
 wire n1457;
 wire n1458;
 wire n1459;
 wire n1460;
 wire n1461;
 wire n1462;
 wire n1463;
 wire n1464;
 wire n1465;
 wire n1466;
 wire n1467;
 wire n1469;
 wire n1470;
 wire n1475;
 wire n1476;
 wire n1477;
 wire n1478;
 wire n1479;
 wire n1480;
 wire n1481;
 wire n1482;
 wire n1483;
 wire n1484;
 wire n1485;
 wire n1486;
 wire n1487;
 wire n1488;
 wire n498;
 wire n499;
 wire n500;
 wire n501;
 wire n502;
 wire n503;
 wire n504;
 wire n505;
 wire n506;
 wire n507;
 wire n508;
 wire n509;
 wire n510;
 wire n511;
 wire n512;
 wire n513;
 wire n514;
 wire n515;
 wire n516;
 wire n517;
 wire n518;
 wire n519;
 wire n520;
 wire n521;
 wire n522;
 wire n523;
 wire n524;
 wire n525;
 wire n526;
 wire n527;
 wire n528;
 wire n529;
 wire n530;
 wire n531;
 wire n532;
 wire n533;
 wire n534;
 wire n535;
 wire n536;
 wire n537;
 wire n538;
 wire n539;
 wire n540;
 wire n541;
 wire n542;
 wire n543;
 wire n544;
 wire n545;
 wire n546;
 wire n547;
 wire n548;
 wire n549;
 wire n550;
 wire n551;
 wire n552;
 wire n553;
 wire n554;
 wire n555;
 wire n556;
 wire n557;
 wire n558;
 wire n559;
 wire n560;
 wire n561;
 wire n562;
 wire n563;
 wire n564;
 wire n565;
 wire n566;
 wire n567;
 wire n568;
 wire n569;
 wire n570;
 wire n571;
 wire n572;
 wire n573;
 wire n574;
 wire n575;
 wire n576;
 wire n577;
 wire n578;
 wire n579;
 wire n580;
 wire n581;
 wire n582;
 wire n583;
 wire n584;
 wire n585;
 wire n586;
 wire n587;
 wire n588;
 wire n589;
 wire n590;
 wire n591;
 wire n592;
 wire n593;
 wire n594;
 wire n595;
 wire n596;
 wire n597;
 wire n598;
 wire n599;
 wire n600;
 wire n601;
 wire n602;
 wire n603;
 wire n604;
 wire n605;
 wire n606;
 wire n607;
 wire n608;
 wire n609;
 wire n610;
 wire n611;
 wire n612;
 wire n613;
 wire n614;
 wire n615;
 wire n616;
 wire n617;
 wire n618;
 wire n619;
 wire n620;
 wire n621;
 wire n622;
 wire n623;
 wire n624;
 wire n625;
 wire n626;
 wire n627;
 wire n628;
 wire n629;
 wire n630;
 wire n631;
 wire n632;
 wire n633;
 wire n634;
 wire n635;
 wire n636;
 wire n637;
 wire n638;
 wire n639;
 wire n640;
 wire n641;
 wire n642;
 wire n643;
 wire n644;
 wire n645;
 wire n646;
 wire n647;
 wire n648;
 wire n649;
 wire n650;
 wire n651;
 wire n652;
 wire n653;
 wire n654;
 wire n655;
 wire n656;
 wire n657;
 wire n658;
 wire n659;
 wire n660;
 wire n661;
 wire n662;
 wire n663;
 wire n664;
 wire n665;
 wire n666;
 wire n667;
 wire n668;
 wire n669;
 wire n670;
 wire n671;
 wire n672;
 wire n673;
 wire n674;
 wire n675;
 wire n676;
 wire n677;
 wire n678;
 wire n679;
 wire n680;
 wire n681;
 wire n682;
 wire n683;
 wire n684;
 wire n685;
 wire n686;
 wire n687;
 wire n688;
 wire n689;
 wire n690;
 wire n691;
 wire n692;
 wire n693;
 wire n694;
 wire n695;
 wire n696;
 wire n697;
 wire n698;
 wire n699;
 wire n700;
 wire n701;
 wire n702;
 wire n703;
 wire n704;
 wire n705;
 wire n706;
 wire n707;
 wire n708;
 wire n709;
 wire n710;
 wire n711;
 wire n712;
 wire n713;
 wire n714;
 wire n715;
 wire n716;
 wire n717;
 wire n718;
 wire n719;
 wire n720;
 wire n721;
 wire n722;
 wire n723;
 wire n724;
 wire n725;
 wire n726;
 wire n727;
 wire n728;
 wire n729;
 wire n730;
 wire n731;
 wire n732;
 wire n733;
 wire n734;
 wire n735;
 wire n736;
 wire n737;
 wire n738;
 wire n739;
 wire n740;
 wire n741;
 wire n742;
 wire n743;
 wire n744;
 wire n745;
 wire n746;
 wire n747;
 wire n748;
 wire n749;
 wire n750;
 wire n751;
 wire n752;
 wire n753;
 wire n754;
 wire n755;
 wire n756;
 wire n757;
 wire n758;
 wire n759;
 wire n760;
 wire n761;
 wire n762;
 wire n763;
 wire n764;
 wire n765;
 wire n766;
 wire n767;
 wire n768;
 wire n769;
 wire n770;
 wire n771;
 wire n772;
 wire n773;
 wire n774;
 wire n775;
 wire n776;
 wire n777;
 wire n778;
 wire n779;
 wire n780;
 wire n781;
 wire n782;
 wire n783;
 wire n784;
 wire n785;
 wire n786;
 wire n787;
 wire n788;
 wire n789;
 wire n790;
 wire n791;
 wire n792;
 wire n793;
 wire n794;
 wire n795;
 wire n796;
 wire n797;
 wire n798;
 wire n799;
 wire n800;
 wire n801;
 wire n802;
 wire n803;
 wire n804;
 wire n805;
 wire n806;
 wire n807;
 wire n808;
 wire n809;
 wire n810;
 wire n811;
 wire n812;
 wire n813;
 wire n814;
 wire n815;
 wire n816;
 wire n817;
 wire n818;
 wire n819;
 wire n820;
 wire n821;
 wire n822;
 wire n823;
 wire n824;
 wire n825;
 wire n826;
 wire n827;
 wire n828;
 wire n829;
 wire n830;
 wire n831;
 wire n832;
 wire n833;
 wire n834;
 wire n835;
 wire n836;
 wire n837;
 wire n838;
 wire n839;
 wire n840;
 wire n841;
 wire n842;
 wire n843;
 wire n844;
 wire n845;
 wire n846;
 wire n847;
 wire n848;
 wire n849;
 wire n850;
 wire n851;
 wire n852;
 wire n853;
 wire n854;
 wire n855;
 wire n856;
 wire n857;
 wire n858;
 wire n859;
 wire n860;
 wire n861;
 wire n862;
 wire n863;
 wire n864;
 wire n865;
 wire n866;
 wire n867;
 wire n868;
 wire n869;
 wire n870;
 wire n871;
 wire n872;
 wire n873;
 wire n874;
 wire n875;
 wire n876;
 wire n877;
 wire n878;
 wire n879;
 wire n880;
 wire n881;
 wire n882;
 wire n883;
 wire n884;
 wire n885;
 wire n886;
 wire n887;
 wire n888;
 wire n889;
 wire n890;
 wire n891;
 wire n892;
 wire n893;
 wire n894;
 wire n895;
 wire n896;
 wire n897;
 wire n898;
 wire n899;
 wire n900;
 wire n901;
 wire n902;
 wire n903;
 wire n904;
 wire n905;
 wire n906;
 wire n907;
 wire n908;
 wire n909;
 wire n910;
 wire n911;
 wire n912;
 wire n913;
 wire n914;
 wire n915;
 wire n916;
 wire n917;
 wire n918;
 wire n919;
 wire n920;
 wire n921;
 wire n922;
 wire n923;
 wire n924;
 wire n925;
 wire n926;
 wire n927;
 wire n928;
 wire n929;
 wire n930;
 wire n931;
 wire n932;
 wire n933;
 wire n934;
 wire n935;
 wire n936;
 wire n937;
 wire n938;
 wire n939;
 wire n940;
 wire n941;
 wire n942;
 wire n943;
 wire n944;
 wire n945;
 wire n946;
 wire n947;
 wire n948;
 wire n949;
 wire n950;
 wire n951;
 wire n952;
 wire n953;
 wire n954;
 wire n955;
 wire n956;
 wire n957;
 wire n958;
 wire n959;
 wire n960;
 wire n961;
 wire n962;
 wire n963;
 wire n964;
 wire n965;
 wire n966;
 wire n967;
 wire n968;
 wire n969;
 wire n970;
 wire n971;
 wire n972;
 wire n973;
 wire n974;
 wire n975;
 wire n976;
 wire n977;
 wire n978;
 wire n979;
 wire n980;
 wire n981;
 wire n982;
 wire n983;
 wire n984;
 wire n985;
 wire n986;
 wire n987;
 wire n988;
 wire n989;
 wire n990;
 wire n991;
 wire n992;
 wire n993;
 wire n994;
 wire n995;
 wire n996;
 wire n997;
 wire clknet_leaf_0_PCLK;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire clknet_leaf_1_PCLK;
 wire clknet_leaf_2_PCLK;
 wire clknet_leaf_3_PCLK;
 wire clknet_leaf_4_PCLK;
 wire clknet_leaf_5_PCLK;
 wire clknet_leaf_6_PCLK;
 wire clknet_leaf_7_PCLK;
 wire clknet_leaf_8_PCLK;
 wire clknet_leaf_9_PCLK;
 wire clknet_leaf_10_PCLK;
 wire clknet_leaf_11_PCLK;
 wire clknet_leaf_12_PCLK;
 wire clknet_leaf_13_PCLK;
 wire clknet_leaf_14_PCLK;
 wire clknet_leaf_15_PCLK;
 wire clknet_leaf_16_PCLK;
 wire clknet_leaf_17_PCLK;
 wire clknet_leaf_18_PCLK;
 wire clknet_leaf_19_PCLK;
 wire clknet_0_PCLK;
 wire clknet_1_0__leaf_PCLK;
 wire clknet_1_1__leaf_PCLK;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;

 sky130_fd_sc_hd__or4_1 U1032 (.A(n1326),
    .B(n1325),
    .C(n1324),
    .D(n1323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1351));
 sky130_fd_sc_hd__or4_1 U1033 (.A(n1355),
    .B(n1354),
    .C(n1353),
    .D(n1352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1381));
 sky130_fd_sc_hd__or4_1 U1034 (.A(n1219),
    .B(n1218),
    .C(n1217),
    .D(n1216),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1244));
 sky130_fd_sc_hd__or4_1 U1035 (.A(n1253),
    .B(n1252),
    .C(n1251),
    .D(n1250),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1269));
 sky130_fd_sc_hd__or4_1 U1036 (.A(n1278),
    .B(n1277),
    .C(n1276),
    .D(n1275),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1321));
 sky130_fd_sc_hd__or4_1 U1037 (.A(n1274),
    .B(n1273),
    .C(n1272),
    .D(n1271),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1322));
 sky130_fd_sc_hd__or4_1 U1038 (.A(n1330),
    .B(n1329),
    .C(n1328),
    .D(n1327),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1350));
 sky130_fd_sc_hd__or4_1 U1039 (.A(n1359),
    .B(n1358),
    .C(n1357),
    .D(n1356),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1380));
 sky130_fd_sc_hd__or4_1 U1040 (.A(n1164),
    .B(n1163),
    .C(n1162),
    .D(n1161),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1183));
 sky130_fd_sc_hd__or4_1 U1041 (.A(n1345),
    .B(n1344),
    .C(n1343),
    .D(n1342),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1346));
 sky130_fd_sc_hd__or4_4 U1042 (.A(n1341),
    .B(n1340),
    .C(n1339),
    .D(n1338),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1347));
 sky130_fd_sc_hd__or4_4 U1043 (.A(n1195),
    .B(n1192),
    .C(n1193),
    .D(n1194),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1205));
 sky130_fd_sc_hd__or4_1 U1044 (.A(n1126),
    .B(n1125),
    .C(n1124),
    .D(n1123),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1137));
 sky130_fd_sc_hd__or4_4 U1045 (.A(n1134),
    .B(n1133),
    .C(n1132),
    .D(n1131),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1135));
 sky130_fd_sc_hd__or4_1 U1046 (.A(n1172),
    .B(n1171),
    .C(n1170),
    .D(n1169),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1180));
 sky130_fd_sc_hd__or2_1 U1047 (.A(n1261),
    .B(n1260),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1265));
 sky130_fd_sc_hd__mux2_1 U1048 (.A0(net638),
    .A1(net123),
    .S(n1470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n678));
 sky130_fd_sc_hd__nand2_2 U1049 (.A(net620),
    .B(n1407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1470));
 sky130_fd_sc_hd__and2_4 U1050 (.A(net12),
    .B(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1038));
 sky130_fd_sc_hd__or2_1 U1051 (.A(n1475),
    .B(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net79));
 sky130_fd_sc_hd__or2_4 U1052 (.A(n1314),
    .B(n1315),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1316));
 sky130_fd_sc_hd__or4_1 U1053 (.A(n1235),
    .B(n1234),
    .C(n1233),
    .D(n1232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1241));
 sky130_fd_sc_hd__or4_4 U1054 (.A(n1371),
    .B(n1370),
    .C(n1369),
    .D(n1368),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1377));
 sky130_fd_sc_hd__nand4bb_4 U1055 (.A_N(n1037),
    .B_N(n1036),
    .C(n1035),
    .D(n1034),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1044));
 sky130_fd_sc_hd__or3_4 U1056 (.A(n1112),
    .B(n1111),
    .C(n1110),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net93));
 sky130_fd_sc_hd__or3_1 U1057 (.A(n1137),
    .B(n1136),
    .C(n1135),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1138));
 sky130_fd_sc_hd__nand4bb_2 U1058 (.A_N(n1097),
    .B_N(n1096),
    .C(n1095),
    .D(n1094),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1098));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_0_PCLK));
 sky130_fd_sc_hd__inv_2 U1060 (.A(net704),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(PREADY));
 sky130_fd_sc_hd__nor2_1 U1061 (.A(n1101),
    .B(n1281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1000));
 sky130_fd_sc_hd__nor2_2 U1062 (.A(n1117),
    .B(n1281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1001));
 sky130_fd_sc_hd__nor2_8 U1063 (.A(n1015),
    .B(net14),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1033));
 sky130_fd_sc_hd__or4_1 U1064 (.A(n1239),
    .B(n1238),
    .C(n1237),
    .D(n1236),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1240));
 sky130_fd_sc_hd__or4_1 U1065 (.A(n1375),
    .B(n1374),
    .C(n1373),
    .D(n1372),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1376));
 sky130_fd_sc_hd__or4_4 U1066 (.A(n1201),
    .B(n1200),
    .C(n1199),
    .D(n1198),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1202));
 sky130_fd_sc_hd__or4_1 U1067 (.A(n1212),
    .B(n1211),
    .C(n1210),
    .D(n1209),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1245));
 sky130_fd_sc_hd__or4_1 U1068 (.A(n1249),
    .B(n1248),
    .C(n1247),
    .D(n1246),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1270));
 sky130_fd_sc_hd__clkbuf_4 U1069 (.A(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1466));
 sky130_fd_sc_hd__or3_4 U1070 (.A(n1160),
    .B(n1159),
    .C(n1158),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net92));
 sky130_fd_sc_hd__inv_6 U1071 (.A(n1297),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(net85));
 sky130_fd_sc_hd__nor2_1 U1072 (.A(net2),
    .B(net3),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1003));
 sky130_fd_sc_hd__nor2_1 U1073 (.A(net4),
    .B(net5),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1002));
 sky130_fd_sc_hd__nand2_2 U1074 (.A(n1002),
    .B(n1003),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1008));
 sky130_fd_sc_hd__nor2_1 U1075 (.A(net6),
    .B(net7),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1006));
 sky130_fd_sc_hd__nor2_2 U1076 (.A(net1),
    .B(net8),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1005));
 sky130_fd_sc_hd__nor2_2 U1077 (.A(net16),
    .B(net15),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1004));
 sky130_fd_sc_hd__nand3_4 U1078 (.A(n1006),
    .B(n1005),
    .C(n1004),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1007));
 sky130_fd_sc_hd__nor2_8 U1079 (.A(n1007),
    .B(n1008),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1010));
 sky130_fd_sc_hd__nor2_8 U1080 (.A(net12),
    .B(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1013));
 sky130_fd_sc_hd__clkinv_4 U1081 (.A(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1023));
 sky130_fd_sc_hd__nand2_8 U1082 (.A(n1013),
    .B(n1023),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1215));
 sky130_fd_sc_hd__and2_1 U1083 (.A(net13),
    .B(net14),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1295));
 sky130_fd_sc_hd__nand2_1 U1084 (.A(n1215),
    .B(n1295),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1009));
 sky130_fd_sc_hd__nand2_4 U1085 (.A(n1010),
    .B(n1009),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1221));
 sky130_fd_sc_hd__inv_2 U1086 (.A(n1221),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1297));
 sky130_fd_sc_hd__clkbuf_1 U1087 (.A(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net86));
 sky130_fd_sc_hd__inv_2 U1088 (.A(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1021));
 sky130_fd_sc_hd__nand3_4 U1089 (.A(n1023),
    .B(n1021),
    .C(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1122));
 sky130_fd_sc_hd__inv_6 U1090 (.A(n1010),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1015));
 sky130_fd_sc_hd__inv_2 U1091 (.A(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1032));
 sky130_fd_sc_hd__nor2_2 U1092 (.A(net13),
    .B(n1032),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1011));
 sky130_fd_sc_hd__nand2_8 U1093 (.A(n1033),
    .B(n1011),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1214));
 sky130_fd_sc_hd__nor2_8 U1094 (.A(n1122),
    .B(n1214),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1012));
 sky130_fd_sc_hd__nand2_8 U1095 (.A(net715),
    .B(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1117));
 sky130_fd_sc_hd__a22o_1 U1096 (.A1(net398),
    .A2(net615),
    .B1(net194),
    .B2(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1475));
 sky130_fd_sc_hd__or4_4 U1097 (.A(n1476),
    .B(n1049),
    .C(net619),
    .D(n1048),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1051));
 sky130_fd_sc_hd__nor2_4 U1098 (.A(n1016),
    .B(n1015),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1017));
 sky130_fd_sc_hd__nand2_8 U1099 (.A(n1017),
    .B(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1220));
 sky130_fd_sc_hd__nor2_8 U1100 (.A(n1117),
    .B(n1220),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1469));
 sky130_fd_sc_hd__a22o_1 U1101 (.A1(net612),
    .A2(net513),
    .B1(n1469),
    .B2(net200),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1031));
 sky130_fd_sc_hd__nand2_8 U1102 (.A(n1017),
    .B(n1032),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1281));
 sky130_fd_sc_hd__nor2_4 U1103 (.A(n1122),
    .B(n1281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1399));
 sky130_fd_sc_hd__inv_2 U1104 (.A(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1024));
 sky130_fd_sc_hd__nand2_8 U1105 (.A(n1038),
    .B(n1024),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1290));
 sky130_fd_sc_hd__nor2_2 U1106 (.A(net9),
    .B(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1018));
 sky130_fd_sc_hd__nand2_8 U1107 (.A(n1033),
    .B(n1018),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1213));
 sky130_fd_sc_hd__nor2_8 U1108 (.A(n1290),
    .B(n1213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1019));
 sky130_fd_sc_hd__a22o_1 U1109 (.A1(net611),
    .A2(net539),
    .B1(n1019),
    .B2(net248),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1020));
 sky130_fd_sc_hd__a211o_1 U1110 (.A1(net129),
    .A2(net613),
    .B1(net619),
    .C1(n1020),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1030));
 sky130_fd_sc_hd__nand3_4 U1111 (.A(n1021),
    .B(net10),
    .C(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1287));
 sky130_fd_sc_hd__nor2_8 U1112 (.A(n1213),
    .B(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1452));
 sky130_fd_sc_hd__nand3_4 U1113 (.A(n1033),
    .B(net13),
    .C(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1231));
 sky130_fd_sc_hd__nor2_8 U1114 (.A(net618),
    .B(n1290),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1408));
 sky130_fd_sc_hd__a22o_1 U1115 (.A1(net717),
    .A2(net354),
    .B1(n1408),
    .B2(net578),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1028));
 sky130_fd_sc_hd__nor2_8 U1116 (.A(n1215),
    .B(n1281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1403));
 sky130_fd_sc_hd__nand3_4 U1117 (.A(n1023),
    .B(net10),
    .C(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1280));
 sky130_fd_sc_hd__nor2_8 U1118 (.A(n1280),
    .B(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1445));
 sky130_fd_sc_hd__a22o_1 U1119 (.A1(net609),
    .A2(net370),
    .B1(n1445),
    .B2(net413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1027));
 sky130_fd_sc_hd__nor2_8 U1120 (.A(n1117),
    .B(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1455));
 sky130_fd_sc_hd__nor2_8 U1121 (.A(n1287),
    .B(n1281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1393));
 sky130_fd_sc_hd__a22o_1 U1122 (.A1(net608),
    .A2(net435),
    .B1(n1393),
    .B2(net224),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1026));
 sky130_fd_sc_hd__nor2_8 U1123 (.A(n1117),
    .B(n1214),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1022));
 sky130_fd_sc_hd__nand3_4 U1124 (.A(n1023),
    .B(n1024),
    .C(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1101));
 sky130_fd_sc_hd__a22o_4 U1125 (.A1(net607),
    .A2(net271),
    .B1(net615),
    .B2(net385),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1025));
 sky130_fd_sc_hd__or4_1 U1126 (.A(n1028),
    .B(n1027),
    .C(n1026),
    .D(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1029));
 sky130_fd_sc_hd__or3_4 U1127 (.A(n1031),
    .B(n1030),
    .C(n1029),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net65));
 sky130_fd_sc_hd__nand3_4 U1128 (.A(n1033),
    .B(net13),
    .C(n1032),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1230));
 sky130_fd_sc_hd__nor2_8 U1129 (.A(n1215),
    .B(n1230),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1434));
 sky130_fd_sc_hd__a22o_2 U1130 (.A1(n1445),
    .A2(net412),
    .B1(n1434),
    .B2(net486),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1037));
 sky130_fd_sc_hd__a22o_1 U1131 (.A1(net608),
    .A2(net438),
    .B1(n1408),
    .B2(net577),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1036));
 sky130_fd_sc_hd__a22oi_4 U1132 (.A1(net613),
    .A2(net128),
    .B1(net717),
    .B2(net349),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1035));
 sky130_fd_sc_hd__a22oi_2 U1133 (.A1(n1019),
    .A2(net247),
    .B1(net609),
    .B2(net369),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1034));
 sky130_fd_sc_hd__nor2_8 U1134 (.A(n1280),
    .B(n1214),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1443));
 sky130_fd_sc_hd__a22o_1 U1135 (.A1(net607),
    .A2(net274),
    .B1(n1443),
    .B2(net261),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1043));
 sky130_fd_sc_hd__nand2_8 U1136 (.A(n1038),
    .B(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1127));
 sky130_fd_sc_hd__nor2_8 U1137 (.A(n1127),
    .B(net712),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1436));
 sky130_fd_sc_hd__a22o_1 U1138 (.A1(n1436),
    .A2(net316),
    .B1(net612),
    .B2(net516),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1042));
 sky130_fd_sc_hd__a21o_1 U1139 (.A1(net611),
    .A2(net538),
    .B1(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1040));
 sky130_fd_sc_hd__a22o_1 U1140 (.A1(n1393),
    .A2(net231),
    .B1(net616),
    .B2(net384),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1039));
 sky130_fd_sc_hd__a211o_1 U1141 (.A1(net606),
    .A2(net199),
    .B1(n1040),
    .C1(n1039),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1041));
 sky130_fd_sc_hd__or4_4 U1142 (.A(n1044),
    .B(n1043),
    .C(n1042),
    .D(n1041),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net64));
 sky130_fd_sc_hd__a22o_2 U1143 (.A1(net614),
    .A2(net378),
    .B1(net718),
    .B2(net593),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1046));
 sky130_fd_sc_hd__a22o_1 U1144 (.A1(net615),
    .A2(net404),
    .B1(n1469),
    .B2(net208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1045));
 sky130_fd_sc_hd__or2_1 U1145 (.A(n1046),
    .B(n1045),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net74));
 sky130_fd_sc_hd__a22o_4 U1146 (.A1(net608),
    .A2(net436),
    .B1(n1012),
    .B2(net514),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1053));
 sky130_fd_sc_hd__a22o_1 U1147 (.A1(net607),
    .A2(net272),
    .B1(net615),
    .B2(net395),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1052));
 sky130_fd_sc_hd__a22o_1 U1148 (.A1(net540),
    .A2(net611),
    .B1(net201),
    .B2(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1476));
 sky130_fd_sc_hd__nand2b_1 U1149 (.A_N(n1290),
    .B(net57),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1283));
 sky130_fd_sc_hd__a22o_1 U1150 (.A1(net613),
    .A2(net130),
    .B1(net717),
    .B2(net355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1049));
 sky130_fd_sc_hd__a22o_1 U1151 (.A1(net609),
    .A2(net371),
    .B1(net718),
    .B2(net579),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1048));
 sky130_fd_sc_hd__nand2b_1 U1152 (.A_N(net59),
    .B(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1294));
 sky130_fd_sc_hd__or3_2 U1153 (.A(n1053),
    .B(n1052),
    .C(n1051),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net66));
 sky130_fd_sc_hd__a22o_1 U1154 (.A1(net608),
    .A2(net441),
    .B1(n1403),
    .B2(net374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1058));
 sky130_fd_sc_hd__a22o_4 U1155 (.A1(net607),
    .A2(net277),
    .B1(n1012),
    .B2(net519),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1057));
 sky130_fd_sc_hd__a22o_1 U1156 (.A1(net616),
    .A2(net400),
    .B1(n1469),
    .B2(net204),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1056));
 sky130_fd_sc_hd__a22o_1 U1157 (.A1(net613),
    .A2(net133),
    .B1(n1408),
    .B2(net552),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1054));
 sky130_fd_sc_hd__a211o_1 U1158 (.A1(net543),
    .A2(n1399),
    .B1(net619),
    .C1(n1054),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1055));
 sky130_fd_sc_hd__or4_4 U1159 (.A(n1058),
    .B(n1057),
    .C(n1056),
    .D(n1055),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net69));
 sky130_fd_sc_hd__a22o_1 U1160 (.A1(net608),
    .A2(net444),
    .B1(n1403),
    .B2(net373),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1063));
 sky130_fd_sc_hd__a22o_4 U1161 (.A1(net607),
    .A2(net280),
    .B1(n1012),
    .B2(net522),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1062));
 sky130_fd_sc_hd__a22o_1 U1162 (.A1(net616),
    .A2(net399),
    .B1(n1469),
    .B2(net203),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1061));
 sky130_fd_sc_hd__a22o_1 U1163 (.A1(net613),
    .A2(net132),
    .B1(n1408),
    .B2(net187),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1059));
 sky130_fd_sc_hd__a211o_1 U1164 (.A1(net542),
    .A2(n1399),
    .B1(net619),
    .C1(n1059),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1060));
 sky130_fd_sc_hd__or4_4 U1165 (.A(n1063),
    .B(n1062),
    .C(n1061),
    .D(n1060),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net68));
 sky130_fd_sc_hd__and2_1 U1166 (.A(n1469),
    .B(net193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net83));
 sky130_fd_sc_hd__a22o_1 U1167 (.A1(net609),
    .A2(net375),
    .B1(net718),
    .B2(net545),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1068));
 sky130_fd_sc_hd__a22o_4 U1168 (.A1(net608),
    .A2(net442),
    .B1(net607),
    .B2(net278),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1067));
 sky130_fd_sc_hd__a22o_1 U1169 (.A1(net612),
    .A2(net520),
    .B1(n1469),
    .B2(net205),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1065));
 sky130_fd_sc_hd__a22o_1 U1170 (.A1(net613),
    .A2(net126),
    .B1(net611),
    .B2(net544),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1064));
 sky130_fd_sc_hd__a211o_1 U1171 (.A1(net616),
    .A2(net401),
    .B1(n1065),
    .C1(n1064),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1066));
 sky130_fd_sc_hd__or3_4 U1172 (.A(n1068),
    .B(n1067),
    .C(n1066),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net70));
 sky130_fd_sc_hd__a22o_1 U1173 (.A1(net609),
    .A2(net372),
    .B1(net718),
    .B2(net185),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1073));
 sky130_fd_sc_hd__a22o_4 U1174 (.A1(net608),
    .A2(net443),
    .B1(net607),
    .B2(net279),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1072));
 sky130_fd_sc_hd__a22o_1 U1175 (.A1(net612),
    .A2(net521),
    .B1(n1469),
    .B2(net202),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1070));
 sky130_fd_sc_hd__a22o_1 U1176 (.A1(net613),
    .A2(net131),
    .B1(net611),
    .B2(net541),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1069));
 sky130_fd_sc_hd__a211o_1 U1177 (.A1(net616),
    .A2(net396),
    .B1(n1070),
    .C1(n1069),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1071));
 sky130_fd_sc_hd__or3_4 U1178 (.A(n1073),
    .B(n1072),
    .C(n1071),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net67));
 sky130_fd_sc_hd__a22o_1 U1179 (.A1(net607),
    .A2(net273),
    .B1(n1393),
    .B2(net230),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1092));
 sky130_fd_sc_hd__nor2_8 U1180 (.A(net707),
    .B(n1220),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1074));
 sky130_fd_sc_hd__a22o_2 U1181 (.A1(n1074),
    .A2(net149),
    .B1(net615),
    .B2(net394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1091));
 sky130_fd_sc_hd__a22oi_1 U1182 (.A1(net612),
    .A2(net515),
    .B1(net606),
    .B2(net221),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1077));
 sky130_fd_sc_hd__nor2_8 U1183 (.A(n1117),
    .B(net705),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1424));
 sky130_fd_sc_hd__a22oi_4 U1184 (.A1(net611),
    .A2(net537),
    .B1(n1424),
    .B2(net568),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1076));
 sky130_fd_sc_hd__a21oi_1 U1185 (.A1(net613),
    .A2(net142),
    .B1(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1075));
 sky130_fd_sc_hd__nand3_1 U1186 (.A(n1077),
    .B(n1076),
    .C(n1075),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1090));
 sky130_fd_sc_hd__a22o_1 U1187 (.A1(n1436),
    .A2(net315),
    .B1(n1434),
    .B2(net485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1088));
 sky130_fd_sc_hd__nor2_8 U1188 (.A(n1127),
    .B(n1213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1438));
 sky130_fd_sc_hd__a22o_1 U1189 (.A1(n1438),
    .A2(net336),
    .B1(n1443),
    .B2(net260),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1087));
 sky130_fd_sc_hd__nor2_8 U1190 (.A(n1122),
    .B(n1220),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1397));
 sky130_fd_sc_hd__a22o_1 U1191 (.A1(n1397),
    .A2(net553),
    .B1(n1445),
    .B2(net421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1082));
 sky130_fd_sc_hd__nor2_8 U1192 (.A(net707),
    .B(n1213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1078));
 sky130_fd_sc_hd__a22o_1 U1193 (.A1(n1019),
    .A2(net256),
    .B1(n1078),
    .B2(net494),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1081));
 sky130_fd_sc_hd__a22o_1 U1194 (.A1(net609),
    .A2(net368),
    .B1(net610),
    .B2(net576),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1080));
 sky130_fd_sc_hd__nor2_8 U1195 (.A(net707),
    .B(net712),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1447));
 sky130_fd_sc_hd__a22o_1 U1196 (.A1(n1447),
    .A2(net426),
    .B1(net717),
    .B2(net348),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1079));
 sky130_fd_sc_hd__nor4_1 U1197 (.A(n1082),
    .B(n1081),
    .C(n1080),
    .D(n1079),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1086));
 sky130_fd_sc_hd__nor2_8 U1198 (.A(net722),
    .B(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1420));
 sky130_fd_sc_hd__a22o_2 U1199 (.A1(net608),
    .A2(net437),
    .B1(n1420),
    .B2(net170),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1084));
 sky130_fd_sc_hd__nor2_8 U1200 (.A(n1215),
    .B(n1220),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1401));
 sky130_fd_sc_hd__nor2_8 U1201 (.A(net618),
    .B(n1127),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1405));
 sky130_fd_sc_hd__a22o_1 U1202 (.A1(n1401),
    .A2(net460),
    .B1(n1405),
    .B2(net296),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1083));
 sky130_fd_sc_hd__nor2_1 U1203 (.A(n1084),
    .B(n1083),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1085));
 sky130_fd_sc_hd__or4bb_4 U1204 (.A(n1088),
    .B(n1087),
    .C_N(n1086),
    .D_N(n1085),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1089));
 sky130_fd_sc_hd__or4_4 U1205 (.A(n1092),
    .B(n1091),
    .C(n1090),
    .D(n1089),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net63));
 sky130_fd_sc_hd__a22o_1 U1206 (.A1(net612),
    .A2(net524),
    .B1(n1469),
    .B2(net220),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1100));
 sky130_fd_sc_hd__nor2_8 U1207 (.A(net708),
    .B(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1418));
 sky130_fd_sc_hd__a22o_1 U1208 (.A1(net614),
    .A2(net141),
    .B1(n1424),
    .B2(net567),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1093));
 sky130_fd_sc_hd__a211o_1 U1209 (.A1(net160),
    .A2(n1418),
    .B1(net619),
    .C1(n1093),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1099));
 sky130_fd_sc_hd__a22o_1 U1210 (.A1(net609),
    .A2(net367),
    .B1(net610),
    .B2(net587),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1097));
 sky130_fd_sc_hd__nor2_8 U1211 (.A(net617),
    .B(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1422));
 sky130_fd_sc_hd__a22o_1 U1212 (.A1(net717),
    .A2(net351),
    .B1(net716),
    .B2(net558),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1096));
 sky130_fd_sc_hd__a22oi_1 U1213 (.A1(net611),
    .A2(net536),
    .B1(net253),
    .B2(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1095));
 sky130_fd_sc_hd__a22oi_4 U1214 (.A1(n1078),
    .A2(net493),
    .B1(n1447),
    .B2(net425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1094));
 sky130_fd_sc_hd__or3_1 U1215 (.A(n1100),
    .B(n1099),
    .C(n1098),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1112));
 sky130_fd_sc_hd__nor2_8 U1216 (.A(net618),
    .B(net707),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1416));
 sky130_fd_sc_hd__a22o_1 U1217 (.A1(n1397),
    .A2(net554),
    .B1(net706),
    .B2(net97),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1105));
 sky130_fd_sc_hd__a22o_2 U1218 (.A1(n1445),
    .A2(net418),
    .B1(net721),
    .B2(net169),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1104));
 sky130_fd_sc_hd__a22o_1 U1219 (.A1(net608),
    .A2(net446),
    .B1(n1401),
    .B2(net459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1103));
 sky130_fd_sc_hd__nor2_8 U1220 (.A(n1287),
    .B(net713),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1450));
 sky130_fd_sc_hd__a22o_1 U1221 (.A1(n1450),
    .A2(net505),
    .B1(net720),
    .B2(net295),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1102));
 sky130_fd_sc_hd__or4_1 U1222 (.A(n1105),
    .B(n1104),
    .C(n1103),
    .D(n1102),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1111));
 sky130_fd_sc_hd__a22o_2 U1223 (.A1(n1443),
    .A2(net268),
    .B1(n1434),
    .B2(net480),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1109));
 sky130_fd_sc_hd__a22o_1 U1224 (.A1(n1438),
    .A2(net333),
    .B1(n1022),
    .B2(net282),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1108));
 sky130_fd_sc_hd__a22o_1 U1225 (.A1(n1436),
    .A2(net318),
    .B1(n1393),
    .B2(net240),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1107));
 sky130_fd_sc_hd__a22o_4 U1226 (.A1(n1074),
    .A2(net150),
    .B1(net615),
    .B2(net393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1106));
 sky130_fd_sc_hd__or4_1 U1227 (.A(n1109),
    .B(n1108),
    .C(n1107),
    .D(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1110));
 sky130_fd_sc_hd__a22o_1 U1228 (.A1(net716),
    .A2(net561),
    .B1(n1397),
    .B2(net181),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1116));
 sky130_fd_sc_hd__nor2_8 U1229 (.A(net711),
    .B(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1430));
 sky130_fd_sc_hd__a22o_1 U1230 (.A1(net609),
    .A2(net362),
    .B1(n1430),
    .B2(net310),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1115));
 sky130_fd_sc_hd__a22o_1 U1231 (.A1(n1445),
    .A2(net409),
    .B1(net706),
    .B2(net100),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1114));
 sky130_fd_sc_hd__nor2_8 U1232 (.A(net711),
    .B(net618),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1428));
 sky130_fd_sc_hd__a22o_1 U1233 (.A1(net721),
    .A2(net175),
    .B1(n1428),
    .B2(net468),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1113));
 sky130_fd_sc_hd__or4_4 U1234 (.A(n1116),
    .B(n1115),
    .C(n1114),
    .D(n1113),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1140));
 sky130_fd_sc_hd__nor2_8 U1235 (.A(n1280),
    .B(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1414));
 sky130_fd_sc_hd__a22o_1 U1236 (.A1(net608),
    .A2(net433),
    .B1(n1414),
    .B2(net112),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1121));
 sky130_fd_sc_hd__nor2_8 U1237 (.A(n1117),
    .B(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1426));
 sky130_fd_sc_hd__a22o_4 U1238 (.A1(n1450),
    .A2(net508),
    .B1(n1426),
    .B2(net473),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1120));
 sky130_fd_sc_hd__a22o_1 U1239 (.A1(n1401),
    .A2(net454),
    .B1(n1443),
    .B2(net257),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1119));
 sky130_fd_sc_hd__a22o_1 U1240 (.A1(net720),
    .A2(net290),
    .B1(n1434),
    .B2(net477),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1118));
 sky130_fd_sc_hd__or4_1 U1241 (.A(n1121),
    .B(n1120),
    .C(n1119),
    .D(n1118),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1139));
 sky130_fd_sc_hd__a22o_1 U1242 (.A1(n1438),
    .A2(net326),
    .B1(n1436),
    .B2(net313),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1126));
 sky130_fd_sc_hd__nor2_8 U1243 (.A(net710),
    .B(n1213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1458));
 sky130_fd_sc_hd__nor2_8 U1244 (.A(n1215),
    .B(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1432));
 sky130_fd_sc_hd__a22o_1 U1245 (.A1(n1458),
    .A2(net115),
    .B1(n1432),
    .B2(net303),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1125));
 sky130_fd_sc_hd__a22o_1 U1246 (.A1(n1074),
    .A2(net146),
    .B1(net607),
    .B2(net269),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1124));
 sky130_fd_sc_hd__a22o_1 U1247 (.A1(n1393),
    .A2(net235),
    .B1(net612),
    .B2(net511),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1123));
 sky130_fd_sc_hd__nor2_8 U1248 (.A(n1290),
    .B(net712),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1440));
 sky130_fd_sc_hd__a22o_1 U1249 (.A1(net606),
    .A2(net215),
    .B1(n1440),
    .B2(net337),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1130));
 sky130_fd_sc_hd__inv_2 U1250 (.A(n1127),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1288));
 sky130_fd_sc_hd__or2_1 U1251 (.A(net617),
    .B(n1127),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1302));
 sky130_fd_sc_hd__nand2b_1 U1252 (.A_N(net13),
    .B(net14),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1016));
 sky130_fd_sc_hd__inv_2 U1253 (.A(n1302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1407));
 sky130_fd_sc_hd__a22o_1 U1254 (.A1(n1407),
    .A2(net123),
    .B1(n1418),
    .B2(net163),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1129));
 sky130_fd_sc_hd__a211o_1 U1255 (.A1(net615),
    .A2(net388),
    .B1(n1130),
    .C1(n1129),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1136));
 sky130_fd_sc_hd__a22o_1 U1256 (.A1(net614),
    .A2(net136),
    .B1(n1424),
    .B2(net573),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1134));
 sky130_fd_sc_hd__a22o_1 U1257 (.A1(net611),
    .A2(net531),
    .B1(n1019),
    .B2(net244),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1133));
 sky130_fd_sc_hd__a22o_1 U1258 (.A1(n1447),
    .A2(net422),
    .B1(n1452),
    .B2(net346),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1132));
 sky130_fd_sc_hd__a22o_1 U1259 (.A1(n1078),
    .A2(net496),
    .B1(net610),
    .B2(net582),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1131));
 sky130_fd_sc_hd__or3_4 U1260 (.A(n1140),
    .B(n1139),
    .C(n1138),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net88));
 sky130_fd_sc_hd__a22o_1 U1261 (.A1(n1418),
    .A2(net159),
    .B1(n1424),
    .B2(net570),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1141));
 sky130_fd_sc_hd__a21o_1 U1262 (.A1(net616),
    .A2(net392),
    .B1(n1141),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1149));
 sky130_fd_sc_hd__a22o_1 U1263 (.A1(net614),
    .A2(net140),
    .B1(n1019),
    .B2(net255),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1148));
 sky130_fd_sc_hd__a22o_1 U1264 (.A1(net611),
    .A2(net535),
    .B1(n1078),
    .B2(net500),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1147));
 sky130_fd_sc_hd__inv_2 U1265 (.A(n1302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1477));
 sky130_fd_sc_hd__a22o_1 U1266 (.A1(net124),
    .A2(n1477),
    .B1(net571),
    .B2(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1197));
 sky130_fd_sc_hd__inv_2 U1267 (.A(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1478));
 sky130_fd_sc_hd__a22o_2 U1268 (.A1(n1397),
    .A2(net156),
    .B1(n1420),
    .B2(net172),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1142));
 sky130_fd_sc_hd__a22o_1 U1269 (.A1(n1478),
    .A2(net550),
    .B1(n1285),
    .B2(net55),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1292));
 sky130_fd_sc_hd__or4_1 U1270 (.A(n1149),
    .B(n1148),
    .C(n1147),
    .D(n1146),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1160));
 sky130_fd_sc_hd__a22o_2 U1271 (.A1(n1445),
    .A2(net420),
    .B1(n1414),
    .B2(net107),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1153));
 sky130_fd_sc_hd__a22o_1 U1272 (.A1(n1455),
    .A2(net445),
    .B1(n1401),
    .B2(net458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1152));
 sky130_fd_sc_hd__a22o_1 U1273 (.A1(n1450),
    .A2(net504),
    .B1(n1405),
    .B2(net294),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1151));
 sky130_fd_sc_hd__a22o_2 U1274 (.A1(n1443),
    .A2(net264),
    .B1(n1434),
    .B2(net479),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1150));
 sky130_fd_sc_hd__or4_1 U1275 (.A(n1153),
    .B(n1152),
    .C(n1151),
    .D(n1150),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1159));
 sky130_fd_sc_hd__a22o_1 U1276 (.A1(n1438),
    .A2(net335),
    .B1(net607),
    .B2(net281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1157));
 sky130_fd_sc_hd__a22o_1 U1277 (.A1(n1436),
    .A2(net317),
    .B1(n1393),
    .B2(net239),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1156));
 sky130_fd_sc_hd__a22o_1 U1278 (.A1(n1074),
    .A2(net145),
    .B1(n1440),
    .B2(net345),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1155));
 sky130_fd_sc_hd__a22o_1 U1279 (.A1(net612),
    .A2(net523),
    .B1(net606),
    .B2(net219),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1154));
 sky130_fd_sc_hd__or4_2 U1280 (.A(n1157),
    .B(n1156),
    .C(n1155),
    .D(n1154),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1158));
 sky130_fd_sc_hd__a22o_1 U1281 (.A1(n1019),
    .A2(net254),
    .B1(net717),
    .B2(net357),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1164));
 sky130_fd_sc_hd__a22o_1 U1282 (.A1(n1078),
    .A2(net497),
    .B1(net610),
    .B2(net585),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1163));
 sky130_fd_sc_hd__a22o_1 U1283 (.A1(net716),
    .A2(net560),
    .B1(n1397),
    .B2(net155),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1162));
 sky130_fd_sc_hd__a22o_1 U1284 (.A1(net609),
    .A2(net365),
    .B1(n1430),
    .B2(net312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1161));
 sky130_fd_sc_hd__a22o_1 U1285 (.A1(n1445),
    .A2(net419),
    .B1(net706),
    .B2(net99),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1168));
 sky130_fd_sc_hd__a22o_4 U1286 (.A1(net608),
    .A2(net448),
    .B1(net721),
    .B2(net171),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1167));
 sky130_fd_sc_hd__a22o_2 U1287 (.A1(n1450),
    .A2(net510),
    .B1(n1414),
    .B2(net106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1166));
 sky130_fd_sc_hd__a22o_1 U1288 (.A1(n1401),
    .A2(net457),
    .B1(n1426),
    .B2(net472),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1165));
 sky130_fd_sc_hd__or4_1 U1289 (.A(n1168),
    .B(n1167),
    .C(n1166),
    .D(n1165),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1182));
 sky130_fd_sc_hd__a22o_1 U1290 (.A1(n1405),
    .A2(net293),
    .B1(n1443),
    .B2(net267),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1172));
 sky130_fd_sc_hd__a22o_1 U1291 (.A1(n1438),
    .A2(net334),
    .B1(n1436),
    .B2(net322),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1171));
 sky130_fd_sc_hd__a22o_1 U1292 (.A1(n1022),
    .A2(net284),
    .B1(n1434),
    .B2(net482),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1170));
 sky130_fd_sc_hd__a22o_1 U1293 (.A1(n1458),
    .A2(net191),
    .B1(n1393),
    .B2(net238),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1169));
 sky130_fd_sc_hd__a22o_1 U1294 (.A1(n1074),
    .A2(net144),
    .B1(n1440),
    .B2(net342),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1179));
 sky130_fd_sc_hd__a22o_4 U1295 (.A1(net612),
    .A2(net526),
    .B1(net616),
    .B2(net391),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1178));
 sky130_fd_sc_hd__a21o_1 U1296 (.A1(net613),
    .A2(net139),
    .B1(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1173));
 sky130_fd_sc_hd__a21o_1 U1297 (.A1(net606),
    .A2(net218),
    .B1(n1173),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1176));
 sky130_fd_sc_hd__a22o_1 U1298 (.A1(net611),
    .A2(net534),
    .B1(n1418),
    .B2(net162),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1175));
 sky130_fd_sc_hd__a22o_1 U1299 (.A1(n1447),
    .A2(net429),
    .B1(n1424),
    .B2(net569),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1174));
 sky130_fd_sc_hd__or3_1 U1300 (.A(n1176),
    .B(n1175),
    .C(n1174),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1177));
 sky130_fd_sc_hd__or4_1 U1301 (.A(n1180),
    .B(n1179),
    .C(n1178),
    .D(n1177),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1181));
 sky130_fd_sc_hd__or3_4 U1302 (.A(n1183),
    .B(n1181),
    .C(n1182),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net91));
 sky130_fd_sc_hd__a22o_1 U1303 (.A1(net609),
    .A2(net363),
    .B1(net706),
    .B2(net103),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1187));
 sky130_fd_sc_hd__a22o_1 U1304 (.A1(n1397),
    .A2(net182),
    .B1(n1445),
    .B2(net416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1186));
 sky130_fd_sc_hd__a22o_1 U1305 (.A1(n1430),
    .A2(net311),
    .B1(net721),
    .B2(net173),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1185));
 sky130_fd_sc_hd__a22o_1 U1306 (.A1(n1455),
    .A2(net434),
    .B1(n1428),
    .B2(net464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1184));
 sky130_fd_sc_hd__or4_4 U1307 (.A(n1187),
    .B(n1186),
    .C(n1185),
    .D(n1184),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1208));
 sky130_fd_sc_hd__a22o_1 U1308 (.A1(n1450),
    .A2(net509),
    .B1(n1414),
    .B2(net108),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1191));
 sky130_fd_sc_hd__a22o_1 U1309 (.A1(n1401),
    .A2(net455),
    .B1(n1426),
    .B2(net476),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1190));
 sky130_fd_sc_hd__a22o_2 U1310 (.A1(n1405),
    .A2(net291),
    .B1(n1443),
    .B2(net265),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1189));
 sky130_fd_sc_hd__a22o_1 U1311 (.A1(n1438),
    .A2(net331),
    .B1(n1432),
    .B2(net302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1188));
 sky130_fd_sc_hd__or4_1 U1312 (.A(n1191),
    .B(n1190),
    .C(n1189),
    .D(n1188),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1207));
 sky130_fd_sc_hd__a22o_1 U1313 (.A1(n1458),
    .A2(net116),
    .B1(n1434),
    .B2(net478),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1195));
 sky130_fd_sc_hd__a22o_1 U1314 (.A1(n1436),
    .A2(net314),
    .B1(net607),
    .B2(net270),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1194));
 sky130_fd_sc_hd__a22o_2 U1315 (.A1(n1074),
    .A2(net147),
    .B1(n1393),
    .B2(net236),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1193));
 sky130_fd_sc_hd__a22o_1 U1316 (.A1(net612),
    .A2(net512),
    .B1(n1440),
    .B2(net343),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1192));
 sky130_fd_sc_hd__a22o_1 U1317 (.A1(net616),
    .A2(net389),
    .B1(net606),
    .B2(net216),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1204));
 sky130_fd_sc_hd__inv_2 U1318 (.A(n1290),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1479));
 sky130_fd_sc_hd__a211o_1 U1319 (.A1(net166),
    .A2(n1418),
    .B1(net85),
    .C1(n1197),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1203));
 sky130_fd_sc_hd__a22o_4 U1320 (.A1(net613),
    .A2(net137),
    .B1(n1019),
    .B2(net251),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1201));
 sky130_fd_sc_hd__a22o_1 U1321 (.A1(net611),
    .A2(net532),
    .B1(n1447),
    .B2(net430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1200));
 sky130_fd_sc_hd__a22o_1 U1322 (.A1(n1078),
    .A2(net498),
    .B1(n1452),
    .B2(net347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1199));
 sky130_fd_sc_hd__a22o_1 U1323 (.A1(n1422),
    .A2(net564),
    .B1(net610),
    .B2(net583),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1198));
 sky130_fd_sc_hd__or4_4 U1324 (.A(n1205),
    .B(n1204),
    .C(n1203),
    .D(n1202),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1206));
 sky130_fd_sc_hd__or3_4 U1325 (.A(n1208),
    .B(n1206),
    .C(n1207),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net89));
 sky130_fd_sc_hd__a22o_1 U1326 (.A1(net608),
    .A2(net450),
    .B1(n1426),
    .B2(net469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1212));
 sky130_fd_sc_hd__a22o_4 U1327 (.A1(n1450),
    .A2(net502),
    .B1(n1401),
    .B2(net451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1211));
 sky130_fd_sc_hd__a22o_1 U1328 (.A1(n1405),
    .A2(net287),
    .B1(n1443),
    .B2(net263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1210));
 sky130_fd_sc_hd__a22o_2 U1329 (.A1(n1438),
    .A2(net330),
    .B1(n1432),
    .B2(net301),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1209));
 sky130_fd_sc_hd__a22o_1 U1330 (.A1(n1436),
    .A2(net324),
    .B1(n1434),
    .B2(net488),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1219));
 sky130_fd_sc_hd__nor2_8 U1331 (.A(n1215),
    .B(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1463));
 sky130_fd_sc_hd__a22o_1 U1332 (.A1(n1463),
    .A2(net223),
    .B1(n1458),
    .B2(net114),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1218));
 sky130_fd_sc_hd__nor2_4 U1333 (.A(n1215),
    .B(n1214),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1460));
 sky130_fd_sc_hd__a22o_1 U1334 (.A1(n1460),
    .A2(net228),
    .B1(net607),
    .B2(net286),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1217));
 sky130_fd_sc_hd__a22o_1 U1335 (.A1(n1074),
    .A2(net151),
    .B1(net612),
    .B2(net528),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1216));
 sky130_fd_sc_hd__a22o_1 U1336 (.A1(n1393),
    .A2(net232),
    .B1(n1440),
    .B2(net341),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1229));
 sky130_fd_sc_hd__a22o_1 U1337 (.A1(net616),
    .A2(net383),
    .B1(net606),
    .B2(net198),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1228));
 sky130_fd_sc_hd__nor2_2 U1338 (.A(n1280),
    .B(n1281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1361));
 sky130_fd_sc_hd__inv_2 U1339 (.A(n1220),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1391));
 sky130_fd_sc_hd__inv_2 U1340 (.A(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1390));
 sky130_fd_sc_hd__a31o_1 U1341 (.A1(n1391),
    .A2(n1390),
    .A3(net551),
    .B1(n1221),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1222));
 sky130_fd_sc_hd__a21o_1 U1342 (.A1(n1418),
    .A2(net157),
    .B1(n1222),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1223));
 sky130_fd_sc_hd__a22o_1 U1343 (.A1(n1479),
    .A2(net56),
    .B1(net58),
    .B2(n1288),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1291));
 sky130_fd_sc_hd__a22o_1 U1344 (.A1(net614),
    .A2(net127),
    .B1(n1407),
    .B2(net186),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1225));
 sky130_fd_sc_hd__a22o_4 U1345 (.A1(net611),
    .A2(net489),
    .B1(n1424),
    .B2(net565),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1224));
 sky130_fd_sc_hd__or3_4 U1346 (.A(n1378),
    .B(n1377),
    .C(n1376),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1379));
 sky130_fd_sc_hd__or3_4 U1347 (.A(n1348),
    .B(n1347),
    .C(n1346),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1349));
 sky130_fd_sc_hd__a22o_1 U1348 (.A1(n1019),
    .A2(net250),
    .B1(n1078),
    .B2(net491),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1235));
 sky130_fd_sc_hd__a22o_1 U1349 (.A1(n1447),
    .A2(net428),
    .B1(n1452),
    .B2(net359),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1234));
 sky130_fd_sc_hd__nor2_4 U1350 (.A(n1290),
    .B(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1410));
 sky130_fd_sc_hd__a22o_1 U1351 (.A1(n1422),
    .A2(net555),
    .B1(n1410),
    .B2(net118),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1233));
 sky130_fd_sc_hd__nor2_8 U1352 (.A(n1280),
    .B(net618),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1412));
 sky130_fd_sc_hd__a22o_2 U1353 (.A1(net610),
    .A2(net590),
    .B1(n1412),
    .B2(net547),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1232));
 sky130_fd_sc_hd__a22o_1 U1354 (.A1(net609),
    .A2(net325),
    .B1(n1416),
    .B2(net94),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1239));
 sky130_fd_sc_hd__a22o_1 U1355 (.A1(n1397),
    .A2(net178),
    .B1(n1430),
    .B2(net308),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1238));
 sky130_fd_sc_hd__a22o_2 U1356 (.A1(n1445),
    .A2(net415),
    .B1(n1420),
    .B2(net167),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1237));
 sky130_fd_sc_hd__a22o_1 U1357 (.A1(n1414),
    .A2(net104),
    .B1(n1428),
    .B2(net462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1236));
 sky130_fd_sc_hd__or3_4 U1358 (.A(n1242),
    .B(n1241),
    .C(n1240),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1243));
 sky130_fd_sc_hd__or3_4 U1359 (.A(n1245),
    .B(n1244),
    .C(n1243),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net73));
 sky130_fd_sc_hd__a22o_1 U1360 (.A1(net609),
    .A2(net364),
    .B1(net718),
    .B2(net584),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1249));
 sky130_fd_sc_hd__a22o_1 U1361 (.A1(n1397),
    .A2(net183),
    .B1(n1416),
    .B2(net98),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1248));
 sky130_fd_sc_hd__a22o_2 U1362 (.A1(n1445),
    .A2(net417),
    .B1(n1430),
    .B2(net309),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1247));
 sky130_fd_sc_hd__a22o_1 U1363 (.A1(net608),
    .A2(net447),
    .B1(net721),
    .B2(net177),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1246));
 sky130_fd_sc_hd__a22o_2 U1364 (.A1(n1450),
    .A2(net506),
    .B1(n1428),
    .B2(net465),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1253));
 sky130_fd_sc_hd__a22o_1 U1365 (.A1(n1401),
    .A2(net456),
    .B1(n1414),
    .B2(net109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1252));
 sky130_fd_sc_hd__a22o_1 U1366 (.A1(n1426),
    .A2(net471),
    .B1(n1405),
    .B2(net292),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1251));
 sky130_fd_sc_hd__a22o_1 U1367 (.A1(n1438),
    .A2(net332),
    .B1(n1443),
    .B2(net266),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1250));
 sky130_fd_sc_hd__a22o_1 U1368 (.A1(n1074),
    .A2(net148),
    .B1(n1440),
    .B2(net344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1267));
 sky130_fd_sc_hd__a22o_1 U1369 (.A1(n1022),
    .A2(net283),
    .B1(n1393),
    .B2(net237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1266));
 sky130_fd_sc_hd__a21o_1 U1370 (.A1(net613),
    .A2(net138),
    .B1(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1255));
 sky130_fd_sc_hd__a22o_4 U1371 (.A1(net612),
    .A2(net525),
    .B1(net615),
    .B2(net390),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1254));
 sky130_fd_sc_hd__a211o_1 U1372 (.A1(net606),
    .A2(net217),
    .B1(n1255),
    .C1(n1254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1261));
 sky130_fd_sc_hd__a211o_1 U1373 (.A1(net586),
    .A2(net610),
    .B1(n1482),
    .C1(n1480),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1146));
 sky130_fd_sc_hd__a211o_1 U1374 (.A1(net96),
    .A2(net714),
    .B1(n1142),
    .C1(n1481),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1480));
 sky130_fd_sc_hd__a22o_1 U1375 (.A1(net557),
    .A2(n1422),
    .B1(net350),
    .B2(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1481));
 sky130_fd_sc_hd__a22o_4 U1376 (.A1(n1452),
    .A2(net356),
    .B1(n1422),
    .B2(net559),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1256));
 sky130_fd_sc_hd__a22o_1 U1377 (.A1(net432),
    .A2(n1447),
    .B1(net366),
    .B2(n1403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1482));
 sky130_fd_sc_hd__a22o_2 U1378 (.A1(n1432),
    .A2(net304),
    .B1(n1434),
    .B2(net481),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1263));
 sky130_fd_sc_hd__a22o_1 U1379 (.A1(n1436),
    .A2(net321),
    .B1(n1458),
    .B2(net190),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1262));
 sky130_fd_sc_hd__nor2_1 U1380 (.A(n1263),
    .B(n1262),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1264));
 sky130_fd_sc_hd__or4b_4 U1381 (.A(n1267),
    .B(n1266),
    .C(n1265),
    .D_N(n1264),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1268));
 sky130_fd_sc_hd__or3_4 U1382 (.A(n1270),
    .B(n1268),
    .C(n1269),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net90));
 sky130_fd_sc_hd__a22o_1 U1383 (.A1(net608),
    .A2(net449),
    .B1(n1414),
    .B2(net105),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1274));
 sky130_fd_sc_hd__a22o_4 U1384 (.A1(n1450),
    .A2(net503),
    .B1(n1426),
    .B2(net470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1273));
 sky130_fd_sc_hd__a22o_1 U1385 (.A1(n1401),
    .A2(net461),
    .B1(net720),
    .B2(net297),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1272));
 sky130_fd_sc_hd__a22o_1 U1386 (.A1(n1438),
    .A2(net329),
    .B1(n1443),
    .B2(net262),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1271));
 sky130_fd_sc_hd__a22o_1 U1387 (.A1(n1432),
    .A2(net300),
    .B1(n1434),
    .B2(net487),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1278));
 sky130_fd_sc_hd__a22o_1 U1388 (.A1(n1436),
    .A2(net323),
    .B1(n1463),
    .B2(net222),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1277));
 sky130_fd_sc_hd__a22o_1 U1389 (.A1(n1458),
    .A2(net113),
    .B1(n1460),
    .B2(net227),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1276));
 sky130_fd_sc_hd__a22o_1 U1390 (.A1(n1074),
    .A2(net143),
    .B1(net607),
    .B2(net285),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1275));
 sky130_fd_sc_hd__a22o_1 U1391 (.A1(n1393),
    .A2(net229),
    .B1(n1440),
    .B2(net340),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1319));
 sky130_fd_sc_hd__a22o_1 U1392 (.A1(net612),
    .A2(net527),
    .B1(net615),
    .B2(net382),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1318));
 sky130_fd_sc_hd__nand2_1 U1393 (.A(n1288),
    .B(net60),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1284));
 sky130_fd_sc_hd__or4_1 U1394 (.A(n1367),
    .B(n1366),
    .C(n1486),
    .D(n1363),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1378));
 sky130_fd_sc_hd__or4_1 U1395 (.A(n1337),
    .B(n1336),
    .C(n1487),
    .D(n1333),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1348));
 sky130_fd_sc_hd__inv_2 U1396 (.A(n1280),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1285));
 sky130_fd_sc_hd__nand2_1 U1397 (.A(n1285),
    .B(net54),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1282));
 sky130_fd_sc_hd__a31o_1 U1398 (.A1(n1284),
    .A2(n1283),
    .A3(n1282),
    .B1(n1281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1299));
 sky130_fd_sc_hd__or4_1 U1399 (.A(n1229),
    .B(n1228),
    .C(n1488),
    .D(n1225),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1242));
 sky130_fd_sc_hd__a211o_1 U1400 (.A1(net575),
    .A2(n1424),
    .B1(n1485),
    .C1(n1483),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1260));
 sky130_fd_sc_hd__o21ai_1 U1401 (.A1(n1292),
    .A2(n1291),
    .B1(n1391),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1298));
 sky130_fd_sc_hd__a211o_1 U1402 (.A1(net161),
    .A2(n1418),
    .B1(n1256),
    .C1(n1484),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1483));
 sky130_fd_sc_hd__a22o_1 U1403 (.A1(net252),
    .A2(n1019),
    .B1(net533),
    .B2(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1484));
 sky130_fd_sc_hd__o211ai_4 U1404 (.A1(net9),
    .A2(net61),
    .B1(n1295),
    .C1(n1294),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1296));
 sky130_fd_sc_hd__nand4_1 U1405 (.A(n1299),
    .B(n1298),
    .C(n1297),
    .D(n1296),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1300));
 sky130_fd_sc_hd__a21oi_1 U1406 (.A1(net606),
    .A2(net192),
    .B1(n1300),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1305));
 sky130_fd_sc_hd__inv_2 U1407 (.A(net184),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1301));
 sky130_fd_sc_hd__o2bb2a_1 U1408 (.A1_N(n1418),
    .A2_N(net158),
    .B1(n1302),
    .B2(n1301),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1304));
 sky130_fd_sc_hd__a22oi_2 U1409 (.A1(net613),
    .A2(net125),
    .B1(net611),
    .B2(net408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1303));
 sky130_fd_sc_hd__nand3_2 U1410 (.A(n1305),
    .B(n1304),
    .C(n1303),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1317));
 sky130_fd_sc_hd__a22o_1 U1411 (.A1(n1019),
    .A2(net249),
    .B1(n1424),
    .B2(net566),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1309));
 sky130_fd_sc_hd__a22o_1 U1412 (.A1(n1078),
    .A2(net492),
    .B1(n1447),
    .B2(net427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1308));
 sky130_fd_sc_hd__a22o_1 U1413 (.A1(n1452),
    .A2(net358),
    .B1(n1422),
    .B2(net556),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1307));
 sky130_fd_sc_hd__a22o_1 U1414 (.A1(n1410),
    .A2(net117),
    .B1(net610),
    .B2(net591),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1306));
 sky130_fd_sc_hd__or4_4 U1415 (.A(n1309),
    .B(n1308),
    .C(n1307),
    .D(n1306),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1315));
 sky130_fd_sc_hd__a22o_1 U1416 (.A1(net609),
    .A2(net243),
    .B1(n1412),
    .B2(net546),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1313));
 sky130_fd_sc_hd__a22o_4 U1417 (.A1(n1397),
    .A2(net154),
    .B1(net95),
    .B2(n1416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1312));
 sky130_fd_sc_hd__a22o_1 U1418 (.A1(n1430),
    .A2(net307),
    .B1(n1420),
    .B2(net168),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1311));
 sky130_fd_sc_hd__a22o_1 U1419 (.A1(n1445),
    .A2(net414),
    .B1(n1428),
    .B2(net463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1310));
 sky130_fd_sc_hd__or4_4 U1420 (.A(n1313),
    .B(n1310),
    .C(n1311),
    .D(n1312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1314));
 sky130_fd_sc_hd__or4_4 U1421 (.A(n1319),
    .B(n1318),
    .C(n1316),
    .D(n1317),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1320));
 sky130_fd_sc_hd__or3_4 U1422 (.A(n1322),
    .B(n1320),
    .C(n1321),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net62));
 sky130_fd_sc_hd__a22o_4 U1423 (.A1(n1450),
    .A2(net507),
    .B1(n1414),
    .B2(net110),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1326));
 sky130_fd_sc_hd__a22o_1 U1424 (.A1(n1426),
    .A2(net475),
    .B1(n1443),
    .B2(net258),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1325));
 sky130_fd_sc_hd__a22o_1 U1425 (.A1(n1401),
    .A2(net453),
    .B1(net720),
    .B2(net289),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1324));
 sky130_fd_sc_hd__a22o_2 U1426 (.A1(n1438),
    .A2(net327),
    .B1(n1434),
    .B2(net484),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1323));
 sky130_fd_sc_hd__a22o_1 U1427 (.A1(n1458),
    .A2(net189),
    .B1(n1432),
    .B2(net298),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1330));
 sky130_fd_sc_hd__a22o_1 U1428 (.A1(n1436),
    .A2(net320),
    .B1(n1460),
    .B2(net226),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1329));
 sky130_fd_sc_hd__a22o_1 U1429 (.A1(n1463),
    .A2(net589),
    .B1(net607),
    .B2(net276),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1328));
 sky130_fd_sc_hd__a22o_1 U1430 (.A1(n1074),
    .A2(net153),
    .B1(n1393),
    .B2(net234),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1327));
 sky130_fd_sc_hd__a22o_2 U1431 (.A1(net612),
    .A2(net518),
    .B1(net615),
    .B2(net387),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1337));
 sky130_fd_sc_hd__a22o_1 U1432 (.A1(net606),
    .A2(net214),
    .B1(n1440),
    .B2(net338),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1336));
 sky130_fd_sc_hd__a21o_1 U1433 (.A1(n1418),
    .A2(net165),
    .B1(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1331));
 sky130_fd_sc_hd__a22o_4 U1434 (.A1(net499),
    .A2(n1078),
    .B1(net431),
    .B2(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1485));
 sky130_fd_sc_hd__a22o_1 U1435 (.A1(net613),
    .A2(net135),
    .B1(n1407),
    .B2(net122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1333));
 sky130_fd_sc_hd__a22o_2 U1436 (.A1(n1399),
    .A2(net530),
    .B1(n1424),
    .B2(net574),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1332));
 sky130_fd_sc_hd__a211o_1 U1437 (.A1(net51),
    .A2(n1361),
    .B1(n1362),
    .C1(n1360),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1486));
 sky130_fd_sc_hd__a211o_1 U1438 (.A1(net53),
    .A2(n1361),
    .B1(n1332),
    .C1(n1331),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1487));
 sky130_fd_sc_hd__a22o_1 U1439 (.A1(n1019),
    .A2(net245),
    .B1(n1447),
    .B2(net423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1341));
 sky130_fd_sc_hd__a22o_1 U1440 (.A1(n1078),
    .A2(net495),
    .B1(n1410),
    .B2(net120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1340));
 sky130_fd_sc_hd__a22o_1 U1441 (.A1(n1452),
    .A2(net353),
    .B1(n1412),
    .B2(net549),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1339));
 sky130_fd_sc_hd__a22o_1 U1442 (.A1(net716),
    .A2(net563),
    .B1(n1408),
    .B2(net581),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1338));
 sky130_fd_sc_hd__a22o_1 U1443 (.A1(net609),
    .A2(net361),
    .B1(n1397),
    .B2(net180),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1345));
 sky130_fd_sc_hd__a22o_4 U1444 (.A1(n1445),
    .A2(net410),
    .B1(net714),
    .B2(net101),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1344));
 sky130_fd_sc_hd__a22o_1 U1445 (.A1(n1430),
    .A2(net305),
    .B1(n1420),
    .B2(net176),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1343));
 sky130_fd_sc_hd__a22o_1 U1446 (.A1(net608),
    .A2(net440),
    .B1(n1428),
    .B2(net466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1342));
 sky130_fd_sc_hd__a211o_1 U1447 (.A1(net52),
    .A2(n1361),
    .B1(n1224),
    .C1(n1223),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1488));
 sky130_fd_sc_hd__or3_4 U1448 (.A(n1351),
    .B(n1350),
    .C(n1349),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net87));
 sky130_fd_sc_hd__a22o_4 U1449 (.A1(n1450),
    .A2(net501),
    .B1(n1414),
    .B2(net111),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1355));
 sky130_fd_sc_hd__a22o_1 U1450 (.A1(n1426),
    .A2(net474),
    .B1(n1443),
    .B2(net259),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1354));
 sky130_fd_sc_hd__a22o_1 U1451 (.A1(n1401),
    .A2(net452),
    .B1(net720),
    .B2(net288),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1353));
 sky130_fd_sc_hd__a22o_2 U1452 (.A1(n1438),
    .A2(net328),
    .B1(n1434),
    .B2(net483),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1352));
 sky130_fd_sc_hd__a22o_1 U1453 (.A1(n1458),
    .A2(net188),
    .B1(n1432),
    .B2(net299),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1359));
 sky130_fd_sc_hd__a22o_1 U1454 (.A1(n1436),
    .A2(net319),
    .B1(n1460),
    .B2(net225),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1358));
 sky130_fd_sc_hd__a22o_1 U1455 (.A1(n1463),
    .A2(net588),
    .B1(net607),
    .B2(net275),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1357));
 sky130_fd_sc_hd__a22o_1 U1456 (.A1(n1074),
    .A2(net152),
    .B1(n1393),
    .B2(net233),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1356));
 sky130_fd_sc_hd__a22o_2 U1457 (.A1(net612),
    .A2(net517),
    .B1(net615),
    .B2(net386),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1367));
 sky130_fd_sc_hd__a22o_1 U1458 (.A1(n1466),
    .A2(net209),
    .B1(n1440),
    .B2(net339),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1366));
 sky130_fd_sc_hd__a21o_1 U1459 (.A1(n1418),
    .A2(net164),
    .B1(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1360));
 sky130_fd_sc_hd__a22o_1 U1461 (.A1(net613),
    .A2(net134),
    .B1(n1407),
    .B2(net121),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1363));
 sky130_fd_sc_hd__a22o_4 U1462 (.A1(net611),
    .A2(net529),
    .B1(n1424),
    .B2(net572),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1362));
 sky130_fd_sc_hd__a22o_1 U1465 (.A1(n1019),
    .A2(net246),
    .B1(n1447),
    .B2(net424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1371));
 sky130_fd_sc_hd__a22o_1 U1466 (.A1(n1078),
    .A2(net490),
    .B1(n1410),
    .B2(net119),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1370));
 sky130_fd_sc_hd__a22o_1 U1467 (.A1(n1452),
    .A2(net352),
    .B1(n1412),
    .B2(net548),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1369));
 sky130_fd_sc_hd__a22o_1 U1468 (.A1(n1422),
    .A2(net562),
    .B1(n1408),
    .B2(net580),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1368));
 sky130_fd_sc_hd__a22o_1 U1469 (.A1(net609),
    .A2(net360),
    .B1(n1397),
    .B2(net179),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1375));
 sky130_fd_sc_hd__a22o_4 U1470 (.A1(n1445),
    .A2(net411),
    .B1(net714),
    .B2(net102),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1374));
 sky130_fd_sc_hd__a22o_1 U1471 (.A1(n1430),
    .A2(net306),
    .B1(n1420),
    .B2(net174),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1373));
 sky130_fd_sc_hd__a22o_1 U1472 (.A1(net608),
    .A2(net439),
    .B1(n1428),
    .B2(net467),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1372));
 sky130_fd_sc_hd__or3_4 U1474 (.A(n1381),
    .B(n1379),
    .C(n1380),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net84));
 sky130_fd_sc_hd__a21o_1 U1475 (.A1(net718),
    .A2(net376),
    .B1(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1383));
 sky130_fd_sc_hd__a22o_1 U1476 (.A1(net616),
    .A2(net402),
    .B1(net613),
    .B2(net241),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1382));
 sky130_fd_sc_hd__a211o_4 U1477 (.A1(net606),
    .A2(net206),
    .B1(n1383),
    .C1(n1382),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net71));
 sky130_fd_sc_hd__a21o_1 U1478 (.A1(net718),
    .A2(net592),
    .B1(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1385));
 sky130_fd_sc_hd__a22o_1 U1479 (.A1(net616),
    .A2(net403),
    .B1(net613),
    .B2(net377),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1384));
 sky130_fd_sc_hd__a211o_4 U1480 (.A1(net606),
    .A2(net207),
    .B1(n1385),
    .C1(n1384),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net72));
 sky130_fd_sc_hd__a22o_1 U1481 (.A1(net606),
    .A2(net210),
    .B1(net614),
    .B2(net379),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1386));
 sky130_fd_sc_hd__a211o_1 U1482 (.A1(net615),
    .A2(net405),
    .B1(net619),
    .C1(n1386),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net75));
 sky130_fd_sc_hd__a22o_1 U1483 (.A1(net606),
    .A2(net212),
    .B1(net614),
    .B2(net381),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1387));
 sky130_fd_sc_hd__a211o_1 U1484 (.A1(net615),
    .A2(net407),
    .B1(net619),
    .C1(n1387),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net77));
 sky130_fd_sc_hd__and3_4 U1485 (.A(net17),
    .B(net50),
    .C(net19),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1462));
 sky130_fd_sc_hd__nand2_8 U1486 (.A(n1074),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1388));
 sky130_fd_sc_hd__mux2_1 U1487 (.A0(net658),
    .A1(net149),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n510));
 sky130_fd_sc_hd__mux2_1 U1488 (.A0(net624),
    .A1(net150),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n509));
 sky130_fd_sc_hd__mux2_1 U1489 (.A0(net627),
    .A1(net145),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n508));
 sky130_fd_sc_hd__mux2_1 U1490 (.A0(net630),
    .A1(net144),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n507));
 sky130_fd_sc_hd__mux2_1 U1491 (.A0(net638),
    .A1(net146),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n504));
 sky130_fd_sc_hd__mux2_1 U1492 (.A0(net635),
    .A1(net147),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n505));
 sky130_fd_sc_hd__mux2_1 U1493 (.A0(net633),
    .A1(net148),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n506));
 sky130_fd_sc_hd__mux2_1 U1494 (.A0(net649),
    .A1(net151),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n501));
 sky130_fd_sc_hd__mux2_1 U1495 (.A0(net645),
    .A1(net152),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n502));
 sky130_fd_sc_hd__mux2_1 U1496 (.A0(net641),
    .A1(net153),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n503));
 sky130_fd_sc_hd__mux2_1 U1497 (.A0(net660),
    .A1(net143),
    .S(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n500));
 sky130_fd_sc_hd__nand2_1 U1498 (.A(net615),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1389));
 sky130_fd_sc_hd__mux2_1 U1499 (.A0(net656),
    .A1(net396),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n525));
 sky130_fd_sc_hd__mux2_1 U1500 (.A0(net655),
    .A1(net399),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n526));
 sky130_fd_sc_hd__mux2_1 U1501 (.A0(net654),
    .A1(net400),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n527));
 sky130_fd_sc_hd__mux2_1 U1502 (.A0(net653),
    .A1(net401),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n528));
 sky130_fd_sc_hd__mux2_1 U1503 (.A0(net29),
    .A1(net402),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n529));
 sky130_fd_sc_hd__mux2_1 U1504 (.A0(net30),
    .A1(net403),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n530));
 sky130_fd_sc_hd__mux2_1 U1505 (.A0(net32),
    .A1(net404),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n531));
 sky130_fd_sc_hd__mux2_1 U1506 (.A0(net33),
    .A1(net405),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n532));
 sky130_fd_sc_hd__mux2_1 U1507 (.A0(net34),
    .A1(net406),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n533));
 sky130_fd_sc_hd__mux2_1 U1508 (.A0(net35),
    .A1(net407),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n534));
 sky130_fd_sc_hd__mux2_1 U1509 (.A0(net36),
    .A1(net397),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n535));
 sky130_fd_sc_hd__mux2_1 U1510 (.A0(net37),
    .A1(net398),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n536));
 sky130_fd_sc_hd__mux2_1 U1511 (.A0(net24),
    .A1(net395),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n524));
 sky130_fd_sc_hd__mux2_1 U1512 (.A0(net650),
    .A1(net383),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n512));
 sky130_fd_sc_hd__mux2_1 U1513 (.A0(net645),
    .A1(net386),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n513));
 sky130_fd_sc_hd__mux2_1 U1514 (.A0(net641),
    .A1(net387),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n514));
 sky130_fd_sc_hd__mux2_1 U1515 (.A0(net638),
    .A1(net388),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n515));
 sky130_fd_sc_hd__mux2_1 U1516 (.A0(net635),
    .A1(net389),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n516));
 sky130_fd_sc_hd__mux2_1 U1517 (.A0(net633),
    .A1(net390),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n517));
 sky130_fd_sc_hd__mux2_1 U1518 (.A0(net630),
    .A1(net391),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n518));
 sky130_fd_sc_hd__mux2_1 U1519 (.A0(net627),
    .A1(net392),
    .S(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n519));
 sky130_fd_sc_hd__mux2_1 U1520 (.A0(net624),
    .A1(net393),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n520));
 sky130_fd_sc_hd__mux2_1 U1521 (.A0(net658),
    .A1(net394),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n521));
 sky130_fd_sc_hd__mux2_1 U1522 (.A0(net657),
    .A1(net384),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n522));
 sky130_fd_sc_hd__mux2_1 U1523 (.A0(net23),
    .A1(net385),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n523));
 sky130_fd_sc_hd__mux2_1 U1524 (.A0(net661),
    .A1(net382),
    .S(net604),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n511));
 sky130_fd_sc_hd__and3_1 U1525 (.A(n1462),
    .B(n1391),
    .C(n1390),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1392));
 sky130_fd_sc_hd__mux2_1 U1526 (.A0(net551),
    .A1(net650),
    .S(n1392),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n538));
 sky130_fd_sc_hd__mux2_1 U1527 (.A0(net550),
    .A1(net661),
    .S(n1392),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n537));
 sky130_fd_sc_hd__nand2_8 U1528 (.A(n1393),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1394));
 sky130_fd_sc_hd__mux2_1 U1529 (.A0(net23),
    .A1(net224),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n551));
 sky130_fd_sc_hd__mux2_1 U1530 (.A0(net662),
    .A1(net229),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n539));
 sky130_fd_sc_hd__mux2_1 U1531 (.A0(net651),
    .A1(net232),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n540));
 sky130_fd_sc_hd__mux2_1 U1532 (.A0(net646),
    .A1(net233),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n541));
 sky130_fd_sc_hd__mux2_1 U1533 (.A0(net642),
    .A1(net234),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n542));
 sky130_fd_sc_hd__mux2_1 U1534 (.A0(net639),
    .A1(net235),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n543));
 sky130_fd_sc_hd__mux2_1 U1535 (.A0(net636),
    .A1(net236),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n544));
 sky130_fd_sc_hd__mux2_1 U1536 (.A0(net632),
    .A1(net237),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n545));
 sky130_fd_sc_hd__mux2_1 U1537 (.A0(net628),
    .A1(net238),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n546));
 sky130_fd_sc_hd__mux2_1 U1538 (.A0(net625),
    .A1(net239),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n547));
 sky130_fd_sc_hd__mux2_1 U1539 (.A0(net623),
    .A1(net240),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n548));
 sky130_fd_sc_hd__mux2_1 U1540 (.A0(net658),
    .A1(net230),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n549));
 sky130_fd_sc_hd__mux2_1 U1541 (.A0(net657),
    .A1(net231),
    .S(n1394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n550));
 sky130_fd_sc_hd__nand2_1 U1542 (.A(n1469),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1395));
 sky130_fd_sc_hd__mux2_1 U1543 (.A0(net41),
    .A1(net193),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n581));
 sky130_fd_sc_hd__mux2_1 U1544 (.A0(net37),
    .A1(net194),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n577));
 sky130_fd_sc_hd__mux2_1 U1545 (.A0(net38),
    .A1(net195),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n578));
 sky130_fd_sc_hd__mux2_1 U1546 (.A0(net39),
    .A1(net196),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n579));
 sky130_fd_sc_hd__mux2_1 U1547 (.A0(net40),
    .A1(net197),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n580));
 sky130_fd_sc_hd__mux2_1 U1548 (.A0(net651),
    .A1(net198),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n553));
 sky130_fd_sc_hd__mux2_1 U1549 (.A0(net645),
    .A1(net209),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n554));
 sky130_fd_sc_hd__mux2_1 U1550 (.A0(net641),
    .A1(net214),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n555));
 sky130_fd_sc_hd__mux2_1 U1551 (.A0(net638),
    .A1(net215),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n556));
 sky130_fd_sc_hd__mux2_1 U1552 (.A0(net636),
    .A1(net216),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n557));
 sky130_fd_sc_hd__mux2_1 U1553 (.A0(net632),
    .A1(net217),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n558));
 sky130_fd_sc_hd__mux2_1 U1554 (.A0(net628),
    .A1(net218),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n559));
 sky130_fd_sc_hd__mux2_1 U1555 (.A0(net625),
    .A1(net219),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n560));
 sky130_fd_sc_hd__mux2_1 U1556 (.A0(net623),
    .A1(net220),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n561));
 sky130_fd_sc_hd__mux2_1 U1557 (.A0(net658),
    .A1(net221),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n562));
 sky130_fd_sc_hd__mux2_1 U1558 (.A0(net657),
    .A1(net199),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n563));
 sky130_fd_sc_hd__mux2_1 U1559 (.A0(net23),
    .A1(net200),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n564));
 sky130_fd_sc_hd__mux2_1 U1560 (.A0(net24),
    .A1(net201),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n565));
 sky130_fd_sc_hd__mux2_1 U1561 (.A0(net656),
    .A1(net202),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n566));
 sky130_fd_sc_hd__mux2_1 U1562 (.A0(net655),
    .A1(net203),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n567));
 sky130_fd_sc_hd__mux2_1 U1563 (.A0(net654),
    .A1(net204),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n568));
 sky130_fd_sc_hd__mux2_1 U1564 (.A0(net653),
    .A1(net205),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n569));
 sky130_fd_sc_hd__mux2_1 U1565 (.A0(net29),
    .A1(net206),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n570));
 sky130_fd_sc_hd__mux2_1 U1566 (.A0(net30),
    .A1(net207),
    .S(net602),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n571));
 sky130_fd_sc_hd__mux2_1 U1567 (.A0(net32),
    .A1(net208),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n572));
 sky130_fd_sc_hd__mux2_1 U1568 (.A0(net33),
    .A1(net210),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n573));
 sky130_fd_sc_hd__mux2_1 U1569 (.A0(net34),
    .A1(net211),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n574));
 sky130_fd_sc_hd__mux2_1 U1570 (.A0(net35),
    .A1(net212),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n575));
 sky130_fd_sc_hd__mux2_1 U1571 (.A0(net36),
    .A1(net213),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n576));
 sky130_fd_sc_hd__mux2_1 U1572 (.A0(net661),
    .A1(net192),
    .S(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n552));
 sky130_fd_sc_hd__nand2_1 U1573 (.A(net614),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1396));
 sky130_fd_sc_hd__mux2_1 U1574 (.A0(net36),
    .A1(net242),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n604));
 sky130_fd_sc_hd__mux2_1 U1575 (.A0(net32),
    .A1(net378),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n600));
 sky130_fd_sc_hd__mux2_1 U1576 (.A0(net33),
    .A1(net379),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n601));
 sky130_fd_sc_hd__mux2_1 U1577 (.A0(net34),
    .A1(net380),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n602));
 sky130_fd_sc_hd__mux2_1 U1578 (.A0(net35),
    .A1(net381),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n603));
 sky130_fd_sc_hd__mux2_1 U1579 (.A0(net30),
    .A1(net377),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n599));
 sky130_fd_sc_hd__mux2_1 U1580 (.A0(net29),
    .A1(net241),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n499));
 sky130_fd_sc_hd__mux2_1 U1581 (.A0(net653),
    .A1(net126),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n598));
 sky130_fd_sc_hd__mux2_1 U1582 (.A0(net650),
    .A1(net127),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n582));
 sky130_fd_sc_hd__mux2_1 U1583 (.A0(net648),
    .A1(net134),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n583));
 sky130_fd_sc_hd__mux2_1 U1584 (.A0(net644),
    .A1(net135),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n584));
 sky130_fd_sc_hd__mux2_1 U1585 (.A0(net639),
    .A1(net136),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n585));
 sky130_fd_sc_hd__mux2_1 U1586 (.A0(net636),
    .A1(net137),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n586));
 sky130_fd_sc_hd__mux2_1 U1587 (.A0(net632),
    .A1(net138),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n587));
 sky130_fd_sc_hd__mux2_1 U1588 (.A0(net628),
    .A1(net139),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n588));
 sky130_fd_sc_hd__mux2_1 U1589 (.A0(net625),
    .A1(net140),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n589));
 sky130_fd_sc_hd__mux2_1 U1590 (.A0(net623),
    .A1(net141),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n590));
 sky130_fd_sc_hd__mux2_1 U1591 (.A0(net658),
    .A1(net142),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n591));
 sky130_fd_sc_hd__mux2_1 U1592 (.A0(net657),
    .A1(net128),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n592));
 sky130_fd_sc_hd__mux2_1 U1593 (.A0(net23),
    .A1(net129),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n593));
 sky130_fd_sc_hd__mux2_1 U1594 (.A0(net24),
    .A1(net130),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n594));
 sky130_fd_sc_hd__mux2_1 U1595 (.A0(net656),
    .A1(net131),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n595));
 sky130_fd_sc_hd__mux2_1 U1596 (.A0(net655),
    .A1(net132),
    .S(net600),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n596));
 sky130_fd_sc_hd__mux2_1 U1597 (.A0(net654),
    .A1(net133),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n597));
 sky130_fd_sc_hd__mux2_1 U1598 (.A0(net661),
    .A1(net125),
    .S(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n498));
 sky130_fd_sc_hd__nand2_8 U1599 (.A(n1397),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1398));
 sky130_fd_sc_hd__mux2_1 U1600 (.A0(net658),
    .A1(net553),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n615));
 sky130_fd_sc_hd__mux2_1 U1601 (.A0(net624),
    .A1(net554),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n614));
 sky130_fd_sc_hd__mux2_1 U1602 (.A0(net630),
    .A1(net155),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n612));
 sky130_fd_sc_hd__mux2_1 U1603 (.A0(net627),
    .A1(net156),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n613));
 sky130_fd_sc_hd__mux2_1 U1604 (.A0(net650),
    .A1(net178),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n606));
 sky130_fd_sc_hd__mux2_1 U1605 (.A0(net648),
    .A1(net179),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n607));
 sky130_fd_sc_hd__mux2_1 U1606 (.A0(net644),
    .A1(net180),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n608));
 sky130_fd_sc_hd__mux2_1 U1607 (.A0(net639),
    .A1(net181),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n609));
 sky130_fd_sc_hd__mux2_1 U1608 (.A0(net635),
    .A1(net182),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n610));
 sky130_fd_sc_hd__mux2_1 U1609 (.A0(net633),
    .A1(net183),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n611));
 sky130_fd_sc_hd__mux2_1 U1610 (.A0(net661),
    .A1(net154),
    .S(n1398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n605));
 sky130_fd_sc_hd__nand2_2 U1611 (.A(net611),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1400));
 sky130_fd_sc_hd__mux2_1 U1612 (.A0(net658),
    .A1(net537),
    .S(n1400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n626));
 sky130_fd_sc_hd__mux2_1 U1613 (.A0(net657),
    .A1(net538),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n627));
 sky130_fd_sc_hd__mux2_1 U1614 (.A0(net23),
    .A1(net539),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n628));
 sky130_fd_sc_hd__mux2_1 U1615 (.A0(net24),
    .A1(net540),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n629));
 sky130_fd_sc_hd__mux2_1 U1616 (.A0(net656),
    .A1(net541),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n630));
 sky130_fd_sc_hd__mux2_1 U1617 (.A0(net655),
    .A1(net542),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n631));
 sky130_fd_sc_hd__mux2_1 U1618 (.A0(net654),
    .A1(net543),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n632));
 sky130_fd_sc_hd__mux2_1 U1619 (.A0(net653),
    .A1(net544),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n633));
 sky130_fd_sc_hd__mux2_1 U1620 (.A0(net646),
    .A1(net529),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n618));
 sky130_fd_sc_hd__mux2_1 U1621 (.A0(net642),
    .A1(net530),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n619));
 sky130_fd_sc_hd__mux2_1 U1622 (.A0(net639),
    .A1(net531),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n620));
 sky130_fd_sc_hd__mux2_1 U1623 (.A0(net636),
    .A1(net532),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n621));
 sky130_fd_sc_hd__mux2_1 U1624 (.A0(net632),
    .A1(net533),
    .S(n1400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n622));
 sky130_fd_sc_hd__mux2_1 U1625 (.A0(net628),
    .A1(net534),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n623));
 sky130_fd_sc_hd__mux2_1 U1626 (.A0(net625),
    .A1(net535),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n624));
 sky130_fd_sc_hd__mux2_1 U1627 (.A0(net623),
    .A1(net536),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n625));
 sky130_fd_sc_hd__mux2_1 U1628 (.A0(net651),
    .A1(net489),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n617));
 sky130_fd_sc_hd__mux2_1 U1629 (.A0(net662),
    .A1(net408),
    .S(net599),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n616));
 sky130_fd_sc_hd__nand2_4 U1630 (.A(n1401),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1402));
 sky130_fd_sc_hd__mux2_1 U1631 (.A0(net632),
    .A1(net456),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n640));
 sky130_fd_sc_hd__mux2_1 U1632 (.A0(net628),
    .A1(net457),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n641));
 sky130_fd_sc_hd__mux2_1 U1633 (.A0(net625),
    .A1(net458),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n642));
 sky130_fd_sc_hd__mux2_1 U1634 (.A0(net623),
    .A1(net459),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n643));
 sky130_fd_sc_hd__mux2_1 U1635 (.A0(net658),
    .A1(net460),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n644));
 sky130_fd_sc_hd__mux2_1 U1636 (.A0(net651),
    .A1(net451),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n635));
 sky130_fd_sc_hd__mux2_1 U1637 (.A0(net646),
    .A1(net452),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n636));
 sky130_fd_sc_hd__mux2_1 U1638 (.A0(net642),
    .A1(net453),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n637));
 sky130_fd_sc_hd__mux2_1 U1639 (.A0(net639),
    .A1(net454),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n638));
 sky130_fd_sc_hd__mux2_1 U1640 (.A0(net636),
    .A1(net455),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n639));
 sky130_fd_sc_hd__mux2_1 U1641 (.A0(net662),
    .A1(net461),
    .S(n1402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n634));
 sky130_fd_sc_hd__nand2_2 U1642 (.A(net609),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1404));
 sky130_fd_sc_hd__mux2_1 U1643 (.A0(net658),
    .A1(net368),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n655));
 sky130_fd_sc_hd__mux2_1 U1644 (.A0(net657),
    .A1(net369),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n656));
 sky130_fd_sc_hd__mux2_1 U1645 (.A0(net23),
    .A1(net370),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n657));
 sky130_fd_sc_hd__mux2_1 U1646 (.A0(net24),
    .A1(net371),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n658));
 sky130_fd_sc_hd__mux2_1 U1647 (.A0(net656),
    .A1(net372),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n659));
 sky130_fd_sc_hd__mux2_1 U1648 (.A0(net655),
    .A1(net373),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n660));
 sky130_fd_sc_hd__mux2_1 U1649 (.A0(net654),
    .A1(net374),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n661));
 sky130_fd_sc_hd__mux2_1 U1650 (.A0(net653),
    .A1(net375),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n662));
 sky130_fd_sc_hd__mux2_1 U1651 (.A0(net648),
    .A1(net360),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n647));
 sky130_fd_sc_hd__mux2_1 U1652 (.A0(net644),
    .A1(net361),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n648));
 sky130_fd_sc_hd__mux2_1 U1653 (.A0(net638),
    .A1(net362),
    .S(n1404),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n649));
 sky130_fd_sc_hd__mux2_1 U1654 (.A0(net635),
    .A1(net363),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n650));
 sky130_fd_sc_hd__mux2_1 U1655 (.A0(net633),
    .A1(net364),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n651));
 sky130_fd_sc_hd__mux2_1 U1656 (.A0(net630),
    .A1(net365),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n652));
 sky130_fd_sc_hd__mux2_1 U1657 (.A0(net627),
    .A1(net366),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n653));
 sky130_fd_sc_hd__mux2_1 U1658 (.A0(net624),
    .A1(net367),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n654));
 sky130_fd_sc_hd__mux2_1 U1659 (.A0(net650),
    .A1(net325),
    .S(net598),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n646));
 sky130_fd_sc_hd__mux2_1 U1660 (.A0(net661),
    .A1(net243),
    .S(n1404),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n645));
 sky130_fd_sc_hd__nand2_4 U1661 (.A(net720),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1406));
 sky130_fd_sc_hd__mux2_1 U1662 (.A0(net633),
    .A1(net292),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n669));
 sky130_fd_sc_hd__mux2_1 U1663 (.A0(net630),
    .A1(net293),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n670));
 sky130_fd_sc_hd__mux2_1 U1664 (.A0(net627),
    .A1(net294),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n671));
 sky130_fd_sc_hd__mux2_1 U1665 (.A0(net624),
    .A1(net295),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n672));
 sky130_fd_sc_hd__mux2_1 U1666 (.A0(net658),
    .A1(net296),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n673));
 sky130_fd_sc_hd__mux2_1 U1667 (.A0(net650),
    .A1(net287),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n664));
 sky130_fd_sc_hd__mux2_1 U1668 (.A0(net648),
    .A1(net288),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n665));
 sky130_fd_sc_hd__mux2_1 U1669 (.A0(net644),
    .A1(net289),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n666));
 sky130_fd_sc_hd__mux2_1 U1670 (.A0(net640),
    .A1(net290),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n667));
 sky130_fd_sc_hd__mux2_1 U1671 (.A0(net635),
    .A1(net291),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n668));
 sky130_fd_sc_hd__mux2_1 U1672 (.A0(net661),
    .A1(net297),
    .S(n1406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n663));
 sky130_fd_sc_hd__mux2_1 U1674 (.A0(net637),
    .A1(net124),
    .S(n1470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n679));
 sky130_fd_sc_hd__mux2_1 U1675 (.A0(net645),
    .A1(net121),
    .S(n1470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n676));
 sky130_fd_sc_hd__mux2_1 U1676 (.A0(net641),
    .A1(net122),
    .S(n1470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n677));
 sky130_fd_sc_hd__mux2_1 U1677 (.A0(net650),
    .A1(net186),
    .S(n1470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n675));
 sky130_fd_sc_hd__mux2_1 U1678 (.A0(net661),
    .A1(net184),
    .S(n1470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n674));
 sky130_fd_sc_hd__nand2_8 U1679 (.A(net718),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1409));
 sky130_fd_sc_hd__mux2_1 U1680 (.A0(net32),
    .A1(net593),
    .S(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n700));
 sky130_fd_sc_hd__mux2_1 U1681 (.A0(net30),
    .A1(net592),
    .S(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n699));
 sky130_fd_sc_hd__mux2_1 U1682 (.A0(net29),
    .A1(net376),
    .S(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n698));
 sky130_fd_sc_hd__mux2_1 U1683 (.A0(net653),
    .A1(net545),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n697));
 sky130_fd_sc_hd__mux2_1 U1684 (.A0(net654),
    .A1(net552),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n696));
 sky130_fd_sc_hd__mux2_1 U1685 (.A0(net655),
    .A1(net187),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n695));
 sky130_fd_sc_hd__mux2_1 U1686 (.A0(net656),
    .A1(net185),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n694));
 sky130_fd_sc_hd__mux2_1 U1687 (.A0(net23),
    .A1(net578),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n692));
 sky130_fd_sc_hd__mux2_1 U1688 (.A0(net24),
    .A1(net579),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n693));
 sky130_fd_sc_hd__mux2_1 U1689 (.A0(net658),
    .A1(net576),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n690));
 sky130_fd_sc_hd__mux2_1 U1690 (.A0(net657),
    .A1(net577),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n691));
 sky130_fd_sc_hd__mux2_1 U1691 (.A0(net625),
    .A1(net586),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n688));
 sky130_fd_sc_hd__mux2_1 U1692 (.A0(net623),
    .A1(net587),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n689));
 sky130_fd_sc_hd__mux2_1 U1693 (.A0(net632),
    .A1(net584),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n686));
 sky130_fd_sc_hd__mux2_1 U1694 (.A0(net628),
    .A1(net585),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n687));
 sky130_fd_sc_hd__mux2_1 U1695 (.A0(net639),
    .A1(net582),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n684));
 sky130_fd_sc_hd__mux2_1 U1696 (.A0(net636),
    .A1(net583),
    .S(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n685));
 sky130_fd_sc_hd__mux2_1 U1697 (.A0(net646),
    .A1(net580),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n682));
 sky130_fd_sc_hd__mux2_1 U1698 (.A0(net642),
    .A1(net581),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n683));
 sky130_fd_sc_hd__mux2_1 U1699 (.A0(net651),
    .A1(net590),
    .S(net597),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n681));
 sky130_fd_sc_hd__mux2_1 U1700 (.A0(net662),
    .A1(net591),
    .S(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n680));
 sky130_fd_sc_hd__nand2_2 U1701 (.A(n1410),
    .B(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1411));
 sky130_fd_sc_hd__mux2_1 U1702 (.A0(net648),
    .A1(net119),
    .S(n1411),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n703));
 sky130_fd_sc_hd__mux2_1 U1703 (.A0(net644),
    .A1(net120),
    .S(n1411),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n704));
 sky130_fd_sc_hd__mux2_1 U1704 (.A0(net661),
    .A1(net117),
    .S(n1411),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n701));
 sky130_fd_sc_hd__mux2_1 U1705 (.A0(net650),
    .A1(net118),
    .S(n1411),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n702));
 sky130_fd_sc_hd__nand2_2 U1706 (.A(n1412),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1413));
 sky130_fd_sc_hd__mux2_1 U1707 (.A0(net646),
    .A1(net548),
    .S(n1413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n707));
 sky130_fd_sc_hd__mux2_1 U1708 (.A0(net642),
    .A1(net549),
    .S(n1413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n708));
 sky130_fd_sc_hd__mux2_1 U1709 (.A0(net662),
    .A1(net546),
    .S(n1413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n705));
 sky130_fd_sc_hd__mux2_1 U1710 (.A0(net651),
    .A1(net547),
    .S(n1413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n706));
 sky130_fd_sc_hd__nand2_8 U1711 (.A(n1414),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1415));
 sky130_fd_sc_hd__mux2_1 U1712 (.A0(net628),
    .A1(net106),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n716));
 sky130_fd_sc_hd__mux2_1 U1713 (.A0(net625),
    .A1(net107),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n717));
 sky130_fd_sc_hd__mux2_1 U1714 (.A0(net635),
    .A1(net108),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n714));
 sky130_fd_sc_hd__mux2_1 U1715 (.A0(net633),
    .A1(net109),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n715));
 sky130_fd_sc_hd__mux2_1 U1716 (.A0(net639),
    .A1(net112),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n713));
 sky130_fd_sc_hd__mux2_1 U1717 (.A0(net642),
    .A1(net110),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n712));
 sky130_fd_sc_hd__mux2_1 U1718 (.A0(net646),
    .A1(net111),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n711));
 sky130_fd_sc_hd__mux2_1 U1719 (.A0(net649),
    .A1(net104),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n710));
 sky130_fd_sc_hd__mux2_1 U1720 (.A0(net660),
    .A1(net105),
    .S(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n709));
 sky130_fd_sc_hd__nand2_8 U1721 (.A(net706),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1417));
 sky130_fd_sc_hd__mux2_1 U1722 (.A0(net625),
    .A1(net96),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n726));
 sky130_fd_sc_hd__mux2_1 U1723 (.A0(net623),
    .A1(net97),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n727));
 sky130_fd_sc_hd__mux2_1 U1724 (.A0(net633),
    .A1(net98),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n724));
 sky130_fd_sc_hd__mux2_1 U1725 (.A0(net629),
    .A1(net99),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n725));
 sky130_fd_sc_hd__mux2_1 U1726 (.A0(net636),
    .A1(net103),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n723));
 sky130_fd_sc_hd__mux2_1 U1727 (.A0(net639),
    .A1(net100),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n722));
 sky130_fd_sc_hd__mux2_1 U1728 (.A0(net642),
    .A1(net101),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n721));
 sky130_fd_sc_hd__mux2_1 U1729 (.A0(net646),
    .A1(net102),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n720));
 sky130_fd_sc_hd__mux2_1 U1730 (.A0(net649),
    .A1(net94),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n719));
 sky130_fd_sc_hd__mux2_1 U1731 (.A0(net660),
    .A1(net95),
    .S(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n718));
 sky130_fd_sc_hd__nand2_8 U1732 (.A(n1418),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1419));
 sky130_fd_sc_hd__mux2_1 U1733 (.A0(net625),
    .A1(net159),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n736));
 sky130_fd_sc_hd__mux2_1 U1734 (.A0(net623),
    .A1(net160),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n737));
 sky130_fd_sc_hd__mux2_1 U1735 (.A0(net632),
    .A1(net161),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n734));
 sky130_fd_sc_hd__mux2_1 U1736 (.A0(net628),
    .A1(net162),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n735));
 sky130_fd_sc_hd__mux2_1 U1737 (.A0(net636),
    .A1(net166),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n733));
 sky130_fd_sc_hd__mux2_1 U1738 (.A0(net639),
    .A1(net163),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n732));
 sky130_fd_sc_hd__mux2_1 U1739 (.A0(net642),
    .A1(net165),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n731));
 sky130_fd_sc_hd__mux2_1 U1740 (.A0(net646),
    .A1(net164),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n730));
 sky130_fd_sc_hd__mux2_1 U1741 (.A0(net651),
    .A1(net157),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n729));
 sky130_fd_sc_hd__mux2_1 U1742 (.A0(net662),
    .A1(net158),
    .S(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n728));
 sky130_fd_sc_hd__nand2_8 U1743 (.A(net721),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1421));
 sky130_fd_sc_hd__mux2_1 U1744 (.A0(net623),
    .A1(net169),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n747));
 sky130_fd_sc_hd__mux2_1 U1745 (.A0(net658),
    .A1(net170),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n748));
 sky130_fd_sc_hd__mux2_1 U1746 (.A0(net629),
    .A1(net171),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n745));
 sky130_fd_sc_hd__mux2_1 U1747 (.A0(net626),
    .A1(net172),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n746));
 sky130_fd_sc_hd__mux2_1 U1748 (.A0(net632),
    .A1(net177),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n744));
 sky130_fd_sc_hd__mux2_1 U1749 (.A0(net636),
    .A1(net173),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n743));
 sky130_fd_sc_hd__mux2_1 U1750 (.A0(net639),
    .A1(net175),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n742));
 sky130_fd_sc_hd__mux2_1 U1751 (.A0(net642),
    .A1(net176),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n741));
 sky130_fd_sc_hd__mux2_1 U1752 (.A0(net646),
    .A1(net174),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n740));
 sky130_fd_sc_hd__mux2_1 U1753 (.A0(net651),
    .A1(net167),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n739));
 sky130_fd_sc_hd__mux2_1 U1754 (.A0(net662),
    .A1(net168),
    .S(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n738));
 sky130_fd_sc_hd__nand2_8 U1755 (.A(net716),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1423));
 sky130_fd_sc_hd__mux2_1 U1756 (.A0(net625),
    .A1(net557),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n757));
 sky130_fd_sc_hd__mux2_1 U1757 (.A0(net623),
    .A1(net558),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n758));
 sky130_fd_sc_hd__mux2_1 U1758 (.A0(net633),
    .A1(net559),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n755));
 sky130_fd_sc_hd__mux2_1 U1759 (.A0(net630),
    .A1(net560),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n756));
 sky130_fd_sc_hd__mux2_1 U1760 (.A0(net636),
    .A1(net564),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n754));
 sky130_fd_sc_hd__mux2_1 U1761 (.A0(net639),
    .A1(net561),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n753));
 sky130_fd_sc_hd__mux2_1 U1762 (.A0(net642),
    .A1(net563),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n752));
 sky130_fd_sc_hd__mux2_1 U1763 (.A0(net646),
    .A1(net562),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n751));
 sky130_fd_sc_hd__mux2_1 U1764 (.A0(net651),
    .A1(net555),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n750));
 sky130_fd_sc_hd__mux2_1 U1765 (.A0(net662),
    .A1(net556),
    .S(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n749));
 sky130_fd_sc_hd__nand2_8 U1766 (.A(n1424),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1425));
 sky130_fd_sc_hd__mux2_1 U1767 (.A0(net623),
    .A1(net567),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n768));
 sky130_fd_sc_hd__mux2_1 U1768 (.A0(net658),
    .A1(net568),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n769));
 sky130_fd_sc_hd__mux2_1 U1769 (.A0(net628),
    .A1(net569),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n766));
 sky130_fd_sc_hd__mux2_1 U1770 (.A0(net625),
    .A1(net570),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n767));
 sky130_fd_sc_hd__mux2_1 U1771 (.A0(net632),
    .A1(net575),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n765));
 sky130_fd_sc_hd__mux2_1 U1772 (.A0(net636),
    .A1(net571),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n764));
 sky130_fd_sc_hd__mux2_1 U1773 (.A0(net639),
    .A1(net573),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n763));
 sky130_fd_sc_hd__mux2_1 U1774 (.A0(net642),
    .A1(net574),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n762));
 sky130_fd_sc_hd__mux2_1 U1775 (.A0(net646),
    .A1(net572),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n761));
 sky130_fd_sc_hd__mux2_1 U1776 (.A0(net651),
    .A1(net565),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n760));
 sky130_fd_sc_hd__mux2_1 U1777 (.A0(net662),
    .A1(net566),
    .S(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n759));
 sky130_fd_sc_hd__nand2_4 U1778 (.A(n1426),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1427));
 sky130_fd_sc_hd__mux2_1 U1779 (.A0(net632),
    .A1(net471),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n776));
 sky130_fd_sc_hd__mux2_1 U1780 (.A0(net628),
    .A1(net472),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n777));
 sky130_fd_sc_hd__mux2_1 U1781 (.A0(net636),
    .A1(net476),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n775));
 sky130_fd_sc_hd__mux2_1 U1782 (.A0(net639),
    .A1(net473),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n774));
 sky130_fd_sc_hd__mux2_1 U1783 (.A0(net642),
    .A1(net475),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n773));
 sky130_fd_sc_hd__mux2_1 U1784 (.A0(net646),
    .A1(net474),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n772));
 sky130_fd_sc_hd__mux2_1 U1785 (.A0(net651),
    .A1(net469),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n771));
 sky130_fd_sc_hd__mux2_1 U1786 (.A0(net662),
    .A1(net470),
    .S(n1427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n770));
 sky130_fd_sc_hd__nand2_4 U1787 (.A(n1428),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1429));
 sky130_fd_sc_hd__mux2_1 U1788 (.A0(net636),
    .A1(net464),
    .S(n1429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n783));
 sky130_fd_sc_hd__mux2_1 U1789 (.A0(net632),
    .A1(net465),
    .S(n1429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n784));
 sky130_fd_sc_hd__mux2_1 U1790 (.A0(net639),
    .A1(net468),
    .S(n1429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n782));
 sky130_fd_sc_hd__mux2_1 U1791 (.A0(net642),
    .A1(net466),
    .S(n1429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n781));
 sky130_fd_sc_hd__mux2_1 U1792 (.A0(net646),
    .A1(net467),
    .S(n1429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n780));
 sky130_fd_sc_hd__mux2_1 U1793 (.A0(net651),
    .A1(net462),
    .S(n1429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n779));
 sky130_fd_sc_hd__mux2_1 U1794 (.A0(net662),
    .A1(net463),
    .S(n1429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n778));
 sky130_fd_sc_hd__nand2_8 U1795 (.A(n1430),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1431));
 sky130_fd_sc_hd__mux2_1 U1796 (.A0(net628),
    .A1(net312),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n792));
 sky130_fd_sc_hd__mux2_1 U1797 (.A0(net632),
    .A1(net309),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n791));
 sky130_fd_sc_hd__mux2_1 U1798 (.A0(net636),
    .A1(net311),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n790));
 sky130_fd_sc_hd__mux2_1 U1799 (.A0(net639),
    .A1(net310),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n789));
 sky130_fd_sc_hd__mux2_1 U1800 (.A0(net641),
    .A1(net305),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n788));
 sky130_fd_sc_hd__mux2_1 U1801 (.A0(net645),
    .A1(net306),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n787));
 sky130_fd_sc_hd__mux2_1 U1802 (.A0(net660),
    .A1(net307),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n785));
 sky130_fd_sc_hd__mux2_1 U1803 (.A0(net649),
    .A1(net308),
    .S(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n786));
 sky130_fd_sc_hd__nand2_8 U1804 (.A(n1432),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1433));
 sky130_fd_sc_hd__mux2_1 U1805 (.A0(net632),
    .A1(net304),
    .S(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n799));
 sky130_fd_sc_hd__mux2_1 U1806 (.A0(net636),
    .A1(net302),
    .S(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n798));
 sky130_fd_sc_hd__mux2_1 U1807 (.A0(net639),
    .A1(net303),
    .S(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n797));
 sky130_fd_sc_hd__mux2_1 U1808 (.A0(net641),
    .A1(net298),
    .S(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n796));
 sky130_fd_sc_hd__mux2_1 U1809 (.A0(net645),
    .A1(net299),
    .S(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n795));
 sky130_fd_sc_hd__mux2_1 U1810 (.A0(net660),
    .A1(net300),
    .S(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n793));
 sky130_fd_sc_hd__mux2_1 U1811 (.A0(net649),
    .A1(net301),
    .S(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n794));
 sky130_fd_sc_hd__nand2_8 U1812 (.A(n1434),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1435));
 sky130_fd_sc_hd__mux2_1 U1813 (.A0(net659),
    .A1(net485),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n810));
 sky130_fd_sc_hd__mux2_1 U1814 (.A0(net657),
    .A1(net486),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n811));
 sky130_fd_sc_hd__mux2_1 U1815 (.A0(net625),
    .A1(net479),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n808));
 sky130_fd_sc_hd__mux2_1 U1816 (.A0(net623),
    .A1(net480),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n809));
 sky130_fd_sc_hd__mux2_1 U1817 (.A0(net632),
    .A1(net481),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n806));
 sky130_fd_sc_hd__mux2_1 U1818 (.A0(net628),
    .A1(net482),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n807));
 sky130_fd_sc_hd__mux2_1 U1819 (.A0(net638),
    .A1(net477),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n804));
 sky130_fd_sc_hd__mux2_1 U1820 (.A0(net635),
    .A1(net478),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n805));
 sky130_fd_sc_hd__mux2_1 U1821 (.A0(net645),
    .A1(net483),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n802));
 sky130_fd_sc_hd__mux2_1 U1822 (.A0(net641),
    .A1(net484),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n803));
 sky130_fd_sc_hd__mux2_1 U1823 (.A0(net660),
    .A1(net487),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n800));
 sky130_fd_sc_hd__mux2_1 U1824 (.A0(net649),
    .A1(net488),
    .S(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n801));
 sky130_fd_sc_hd__nand2_8 U1825 (.A(n1436),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1437));
 sky130_fd_sc_hd__mux2_1 U1826 (.A0(net658),
    .A1(net315),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n822));
 sky130_fd_sc_hd__mux2_1 U1827 (.A0(net657),
    .A1(net316),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n823));
 sky130_fd_sc_hd__mux2_1 U1828 (.A0(net626),
    .A1(net317),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n820));
 sky130_fd_sc_hd__mux2_1 U1829 (.A0(net624),
    .A1(net318),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n821));
 sky130_fd_sc_hd__mux2_1 U1830 (.A0(net633),
    .A1(net321),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n818));
 sky130_fd_sc_hd__mux2_1 U1831 (.A0(net629),
    .A1(net322),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n819));
 sky130_fd_sc_hd__mux2_1 U1832 (.A0(net638),
    .A1(net313),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n816));
 sky130_fd_sc_hd__mux2_1 U1833 (.A0(net635),
    .A1(net314),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n817));
 sky130_fd_sc_hd__mux2_1 U1834 (.A0(net645),
    .A1(net319),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n814));
 sky130_fd_sc_hd__mux2_1 U1835 (.A0(net641),
    .A1(net320),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n815));
 sky130_fd_sc_hd__mux2_1 U1836 (.A0(net660),
    .A1(net323),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n812));
 sky130_fd_sc_hd__mux2_1 U1837 (.A0(net649),
    .A1(net324),
    .S(n1437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n813));
 sky130_fd_sc_hd__nand2_8 U1838 (.A(n1438),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1439));
 sky130_fd_sc_hd__mux2_1 U1839 (.A0(net659),
    .A1(net336),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n834));
 sky130_fd_sc_hd__mux2_1 U1840 (.A0(net623),
    .A1(net333),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n833));
 sky130_fd_sc_hd__mux2_1 U1841 (.A0(net625),
    .A1(net335),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n832));
 sky130_fd_sc_hd__mux2_1 U1842 (.A0(net628),
    .A1(net334),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n831));
 sky130_fd_sc_hd__mux2_1 U1843 (.A0(net633),
    .A1(net332),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n830));
 sky130_fd_sc_hd__mux2_1 U1844 (.A0(net637),
    .A1(net331),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n829));
 sky130_fd_sc_hd__mux2_1 U1845 (.A0(net638),
    .A1(net326),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n828));
 sky130_fd_sc_hd__mux2_1 U1846 (.A0(net641),
    .A1(net327),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n827));
 sky130_fd_sc_hd__mux2_1 U1847 (.A0(net645),
    .A1(net328),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n826));
 sky130_fd_sc_hd__mux2_1 U1848 (.A0(net660),
    .A1(net329),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n824));
 sky130_fd_sc_hd__mux2_1 U1849 (.A0(net649),
    .A1(net330),
    .S(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n825));
 sky130_fd_sc_hd__nand2_8 U1850 (.A(n1440),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1441));
 sky130_fd_sc_hd__mux2_1 U1851 (.A0(net625),
    .A1(net345),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n843));
 sky130_fd_sc_hd__mux2_1 U1852 (.A0(net628),
    .A1(net342),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n842));
 sky130_fd_sc_hd__mux2_1 U1853 (.A0(net632),
    .A1(net344),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n841));
 sky130_fd_sc_hd__mux2_1 U1854 (.A0(net635),
    .A1(net343),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n840));
 sky130_fd_sc_hd__mux2_1 U1855 (.A0(net638),
    .A1(net337),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n839));
 sky130_fd_sc_hd__mux2_1 U1856 (.A0(net641),
    .A1(net338),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n838));
 sky130_fd_sc_hd__mux2_1 U1857 (.A0(net645),
    .A1(net339),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n837));
 sky130_fd_sc_hd__mux2_1 U1858 (.A0(net660),
    .A1(net340),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n835));
 sky130_fd_sc_hd__mux2_1 U1859 (.A0(net649),
    .A1(net341),
    .S(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n836));
 sky130_fd_sc_hd__nand2_8 U1860 (.A(n1019),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1442));
 sky130_fd_sc_hd__mux2_1 U1861 (.A0(net657),
    .A1(net247),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n855));
 sky130_fd_sc_hd__mux2_1 U1862 (.A0(net23),
    .A1(net248),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n856));
 sky130_fd_sc_hd__mux2_1 U1863 (.A0(net659),
    .A1(net256),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n854));
 sky130_fd_sc_hd__mux2_1 U1864 (.A0(net623),
    .A1(net253),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n853));
 sky130_fd_sc_hd__mux2_1 U1865 (.A0(net625),
    .A1(net255),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n852));
 sky130_fd_sc_hd__mux2_1 U1866 (.A0(net628),
    .A1(net254),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n851));
 sky130_fd_sc_hd__mux2_1 U1867 (.A0(net633),
    .A1(net252),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n850));
 sky130_fd_sc_hd__mux2_1 U1868 (.A0(net635),
    .A1(net251),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n849));
 sky130_fd_sc_hd__mux2_1 U1869 (.A0(net638),
    .A1(net244),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n848));
 sky130_fd_sc_hd__mux2_1 U1870 (.A0(net641),
    .A1(net245),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n847));
 sky130_fd_sc_hd__mux2_1 U1871 (.A0(net645),
    .A1(net246),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n846));
 sky130_fd_sc_hd__mux2_1 U1872 (.A0(net660),
    .A1(net249),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n844));
 sky130_fd_sc_hd__mux2_1 U1873 (.A0(net649),
    .A1(net250),
    .S(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n845));
 sky130_fd_sc_hd__nand2_8 U1874 (.A(n1443),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1444));
 sky130_fd_sc_hd__mux2_1 U1875 (.A0(net659),
    .A1(net260),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n867));
 sky130_fd_sc_hd__mux2_1 U1876 (.A0(net657),
    .A1(net261),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n868));
 sky130_fd_sc_hd__mux2_1 U1877 (.A0(net623),
    .A1(net268),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n866));
 sky130_fd_sc_hd__mux2_1 U1878 (.A0(net625),
    .A1(net264),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n865));
 sky130_fd_sc_hd__mux2_1 U1879 (.A0(net628),
    .A1(net267),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n864));
 sky130_fd_sc_hd__mux2_1 U1880 (.A0(net632),
    .A1(net266),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n863));
 sky130_fd_sc_hd__mux2_1 U1881 (.A0(net635),
    .A1(net265),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n862));
 sky130_fd_sc_hd__mux2_1 U1882 (.A0(net638),
    .A1(net257),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n861));
 sky130_fd_sc_hd__mux2_1 U1883 (.A0(net641),
    .A1(net258),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n860));
 sky130_fd_sc_hd__mux2_1 U1884 (.A0(net645),
    .A1(net259),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n859));
 sky130_fd_sc_hd__mux2_1 U1885 (.A0(net660),
    .A1(net262),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n857));
 sky130_fd_sc_hd__mux2_1 U1886 (.A0(net649),
    .A1(net263),
    .S(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n858));
 sky130_fd_sc_hd__nand2_8 U1887 (.A(n1445),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1446));
 sky130_fd_sc_hd__mux2_1 U1888 (.A0(net657),
    .A1(net412),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n880));
 sky130_fd_sc_hd__mux2_1 U1889 (.A0(net23),
    .A1(net413),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n881));
 sky130_fd_sc_hd__mux2_1 U1890 (.A0(net659),
    .A1(net421),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n879));
 sky130_fd_sc_hd__mux2_1 U1891 (.A0(net623),
    .A1(net418),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n878));
 sky130_fd_sc_hd__mux2_1 U1892 (.A0(net627),
    .A1(net420),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n877));
 sky130_fd_sc_hd__mux2_1 U1893 (.A0(net631),
    .A1(net419),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n876));
 sky130_fd_sc_hd__mux2_1 U1894 (.A0(net634),
    .A1(net417),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n875));
 sky130_fd_sc_hd__mux2_1 U1895 (.A0(net636),
    .A1(net416),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n874));
 sky130_fd_sc_hd__mux2_1 U1896 (.A0(net640),
    .A1(net409),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n873));
 sky130_fd_sc_hd__mux2_1 U1897 (.A0(net642),
    .A1(net410),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n872));
 sky130_fd_sc_hd__mux2_1 U1898 (.A0(net646),
    .A1(net411),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n871));
 sky130_fd_sc_hd__mux2_1 U1899 (.A0(net662),
    .A1(net414),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n869));
 sky130_fd_sc_hd__mux2_1 U1900 (.A0(net651),
    .A1(net415),
    .S(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n870));
 sky130_fd_sc_hd__nand2_8 U1901 (.A(n1447),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1448));
 sky130_fd_sc_hd__mux2_1 U1902 (.A0(net624),
    .A1(net425),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n891));
 sky130_fd_sc_hd__mux2_1 U1903 (.A0(net659),
    .A1(net426),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n892));
 sky130_fd_sc_hd__mux2_1 U1904 (.A0(net627),
    .A1(net432),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n890));
 sky130_fd_sc_hd__mux2_1 U1905 (.A0(net631),
    .A1(net429),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n889));
 sky130_fd_sc_hd__mux2_1 U1906 (.A0(net634),
    .A1(net431),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n888));
 sky130_fd_sc_hd__mux2_1 U1907 (.A0(net637),
    .A1(net430),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n887));
 sky130_fd_sc_hd__mux2_1 U1908 (.A0(net640),
    .A1(net422),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n886));
 sky130_fd_sc_hd__mux2_1 U1909 (.A0(net642),
    .A1(net423),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n885));
 sky130_fd_sc_hd__mux2_1 U1910 (.A0(net646),
    .A1(net424),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n884));
 sky130_fd_sc_hd__mux2_1 U1911 (.A0(net662),
    .A1(net427),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n882));
 sky130_fd_sc_hd__mux2_1 U1912 (.A0(net651),
    .A1(net428),
    .S(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n883));
 sky130_fd_sc_hd__nand2_4 U1913 (.A(n1078),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1449));
 sky130_fd_sc_hd__mux2_1 U1914 (.A0(net624),
    .A1(net493),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n902));
 sky130_fd_sc_hd__mux2_1 U1915 (.A0(net659),
    .A1(net494),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n903));
 sky130_fd_sc_hd__mux2_1 U1916 (.A0(net627),
    .A1(net500),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n901));
 sky130_fd_sc_hd__mux2_1 U1917 (.A0(net631),
    .A1(net497),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n900));
 sky130_fd_sc_hd__mux2_1 U1918 (.A0(net634),
    .A1(net499),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n899));
 sky130_fd_sc_hd__mux2_1 U1919 (.A0(net637),
    .A1(net498),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n898));
 sky130_fd_sc_hd__mux2_1 U1920 (.A0(net640),
    .A1(net496),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n897));
 sky130_fd_sc_hd__mux2_1 U1921 (.A0(net642),
    .A1(net495),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n896));
 sky130_fd_sc_hd__mux2_1 U1922 (.A0(net646),
    .A1(net490),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n895));
 sky130_fd_sc_hd__mux2_1 U1923 (.A0(net651),
    .A1(net491),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n894));
 sky130_fd_sc_hd__mux2_1 U1924 (.A0(net662),
    .A1(net492),
    .S(n1449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n893));
 sky130_fd_sc_hd__nand2_4 U1925 (.A(n1450),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1451));
 sky130_fd_sc_hd__mux2_1 U1926 (.A0(net627),
    .A1(net504),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n912));
 sky130_fd_sc_hd__mux2_1 U1927 (.A0(net624),
    .A1(net505),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n913));
 sky130_fd_sc_hd__mux2_1 U1928 (.A0(net630),
    .A1(net510),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n911));
 sky130_fd_sc_hd__mux2_1 U1929 (.A0(net634),
    .A1(net506),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n910));
 sky130_fd_sc_hd__mux2_1 U1930 (.A0(net637),
    .A1(net509),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n909));
 sky130_fd_sc_hd__mux2_1 U1931 (.A0(net640),
    .A1(net508),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n908));
 sky130_fd_sc_hd__mux2_1 U1932 (.A0(net644),
    .A1(net507),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n907));
 sky130_fd_sc_hd__mux2_1 U1933 (.A0(net648),
    .A1(net501),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n906));
 sky130_fd_sc_hd__mux2_1 U1934 (.A0(net651),
    .A1(net502),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n905));
 sky130_fd_sc_hd__mux2_1 U1935 (.A0(net662),
    .A1(net503),
    .S(n1451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n904));
 sky130_fd_sc_hd__nand2_8 U1936 (.A(net717),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1453));
 sky130_fd_sc_hd__mux2_1 U1937 (.A0(net23),
    .A1(net354),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n926));
 sky130_fd_sc_hd__mux2_1 U1938 (.A0(net24),
    .A1(net355),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n927));
 sky130_fd_sc_hd__mux2_1 U1939 (.A0(net658),
    .A1(net348),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n924));
 sky130_fd_sc_hd__mux2_1 U1940 (.A0(net657),
    .A1(net349),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n925));
 sky130_fd_sc_hd__mux2_1 U1941 (.A0(net627),
    .A1(net350),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n922));
 sky130_fd_sc_hd__mux2_1 U1942 (.A0(net624),
    .A1(net351),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n923));
 sky130_fd_sc_hd__mux2_1 U1943 (.A0(net633),
    .A1(net356),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n920));
 sky130_fd_sc_hd__mux2_1 U1944 (.A0(net629),
    .A1(net357),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n921));
 sky130_fd_sc_hd__mux2_1 U1945 (.A0(net638),
    .A1(net346),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n918));
 sky130_fd_sc_hd__mux2_1 U1946 (.A0(net635),
    .A1(net347),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n919));
 sky130_fd_sc_hd__mux2_1 U1947 (.A0(net645),
    .A1(net352),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n916));
 sky130_fd_sc_hd__mux2_1 U1948 (.A0(net641),
    .A1(net353),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n917));
 sky130_fd_sc_hd__mux2_1 U1949 (.A0(net660),
    .A1(net358),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n914));
 sky130_fd_sc_hd__mux2_1 U1950 (.A0(net649),
    .A1(net359),
    .S(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n915));
 sky130_fd_sc_hd__nand2_2 U1951 (.A(net607),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1454));
 sky130_fd_sc_hd__mux2_1 U1952 (.A0(net654),
    .A1(net277),
    .S(n1454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n944));
 sky130_fd_sc_hd__mux2_1 U1953 (.A0(net653),
    .A1(net278),
    .S(n1454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n945));
 sky130_fd_sc_hd__mux2_1 U1954 (.A0(net656),
    .A1(net279),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n942));
 sky130_fd_sc_hd__mux2_1 U1955 (.A0(net655),
    .A1(net280),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n943));
 sky130_fd_sc_hd__mux2_1 U1956 (.A0(net23),
    .A1(net271),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n940));
 sky130_fd_sc_hd__mux2_1 U1957 (.A0(net24),
    .A1(net272),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n941));
 sky130_fd_sc_hd__mux2_1 U1958 (.A0(net658),
    .A1(net273),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n938));
 sky130_fd_sc_hd__mux2_1 U1959 (.A0(net657),
    .A1(net274),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n939));
 sky130_fd_sc_hd__mux2_1 U1960 (.A0(net626),
    .A1(net281),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n936));
 sky130_fd_sc_hd__mux2_1 U1961 (.A0(net624),
    .A1(net282),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n937));
 sky130_fd_sc_hd__mux2_1 U1962 (.A0(net633),
    .A1(net283),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n934));
 sky130_fd_sc_hd__mux2_1 U1963 (.A0(net629),
    .A1(net284),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n935));
 sky130_fd_sc_hd__mux2_1 U1964 (.A0(net638),
    .A1(net269),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n932));
 sky130_fd_sc_hd__mux2_1 U1965 (.A0(net635),
    .A1(net270),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n933));
 sky130_fd_sc_hd__mux2_1 U1966 (.A0(net645),
    .A1(net275),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n930));
 sky130_fd_sc_hd__mux2_1 U1967 (.A0(net641),
    .A1(net276),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n931));
 sky130_fd_sc_hd__mux2_1 U1968 (.A0(net660),
    .A1(net285),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n928));
 sky130_fd_sc_hd__mux2_1 U1969 (.A0(net649),
    .A1(net286),
    .S(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n929));
 sky130_fd_sc_hd__nand2_2 U1970 (.A(n1455),
    .B(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1456));
 sky130_fd_sc_hd__mux2_1 U1971 (.A0(net654),
    .A1(net441),
    .S(n1456),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n962));
 sky130_fd_sc_hd__mux2_1 U1972 (.A0(net653),
    .A1(net442),
    .S(n1456),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n963));
 sky130_fd_sc_hd__mux2_1 U1973 (.A0(net656),
    .A1(net443),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n960));
 sky130_fd_sc_hd__mux2_1 U1974 (.A0(net655),
    .A1(net444),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n961));
 sky130_fd_sc_hd__mux2_1 U1975 (.A0(net23),
    .A1(net435),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n958));
 sky130_fd_sc_hd__mux2_1 U1976 (.A0(net24),
    .A1(net436),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n959));
 sky130_fd_sc_hd__mux2_1 U1977 (.A0(net659),
    .A1(net437),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n956));
 sky130_fd_sc_hd__mux2_1 U1978 (.A0(net657),
    .A1(net438),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n957));
 sky130_fd_sc_hd__mux2_1 U1979 (.A0(net626),
    .A1(net445),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n954));
 sky130_fd_sc_hd__mux2_1 U1980 (.A0(net624),
    .A1(net446),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n955));
 sky130_fd_sc_hd__mux2_1 U1981 (.A0(net633),
    .A1(net447),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n952));
 sky130_fd_sc_hd__mux2_1 U1982 (.A0(net629),
    .A1(net448),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n953));
 sky130_fd_sc_hd__mux2_1 U1983 (.A0(net638),
    .A1(net433),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n950));
 sky130_fd_sc_hd__mux2_1 U1984 (.A0(net635),
    .A1(net434),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n951));
 sky130_fd_sc_hd__mux2_1 U1985 (.A0(net645),
    .A1(net439),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n948));
 sky130_fd_sc_hd__mux2_1 U1986 (.A0(net641),
    .A1(net440),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n949));
 sky130_fd_sc_hd__mux2_1 U1987 (.A0(net660),
    .A1(net449),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n946));
 sky130_fd_sc_hd__mux2_1 U1988 (.A0(net649),
    .A1(net450),
    .S(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n947));
 sky130_fd_sc_hd__nand2_8 U1989 (.A(net612),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1457));
 sky130_fd_sc_hd__mux2_1 U1990 (.A0(net654),
    .A1(net519),
    .S(n1457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n980));
 sky130_fd_sc_hd__mux2_1 U1991 (.A0(net653),
    .A1(net520),
    .S(n1457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n981));
 sky130_fd_sc_hd__mux2_1 U1992 (.A0(net656),
    .A1(net521),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n978));
 sky130_fd_sc_hd__mux2_1 U1993 (.A0(net655),
    .A1(net522),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n979));
 sky130_fd_sc_hd__mux2_1 U1994 (.A0(net23),
    .A1(net513),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n976));
 sky130_fd_sc_hd__mux2_1 U1995 (.A0(net24),
    .A1(net514),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n977));
 sky130_fd_sc_hd__mux2_1 U1996 (.A0(net659),
    .A1(net515),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n974));
 sky130_fd_sc_hd__mux2_1 U1997 (.A0(net657),
    .A1(net516),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n975));
 sky130_fd_sc_hd__mux2_1 U1998 (.A0(net626),
    .A1(net523),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n972));
 sky130_fd_sc_hd__mux2_1 U1999 (.A0(net624),
    .A1(net524),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n973));
 sky130_fd_sc_hd__mux2_1 U2000 (.A0(net633),
    .A1(net525),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n970));
 sky130_fd_sc_hd__mux2_1 U2001 (.A0(net629),
    .A1(net526),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n971));
 sky130_fd_sc_hd__mux2_1 U2002 (.A0(net638),
    .A1(net511),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n968));
 sky130_fd_sc_hd__mux2_1 U2003 (.A0(net635),
    .A1(net512),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n969));
 sky130_fd_sc_hd__mux2_1 U2004 (.A0(net645),
    .A1(net517),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n966));
 sky130_fd_sc_hd__mux2_1 U2005 (.A0(net641),
    .A1(net518),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n967));
 sky130_fd_sc_hd__mux2_1 U2006 (.A0(net660),
    .A1(net527),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n964));
 sky130_fd_sc_hd__mux2_1 U2007 (.A0(net649),
    .A1(net528),
    .S(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n965));
 sky130_fd_sc_hd__nand2_8 U2008 (.A(n1458),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1459));
 sky130_fd_sc_hd__mux2_1 U2009 (.A0(net634),
    .A1(net190),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n988));
 sky130_fd_sc_hd__mux2_1 U2010 (.A0(net630),
    .A1(net191),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n989));
 sky130_fd_sc_hd__mux2_1 U2011 (.A0(net638),
    .A1(net115),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n986));
 sky130_fd_sc_hd__mux2_1 U2012 (.A0(net635),
    .A1(net116),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n987));
 sky130_fd_sc_hd__mux2_1 U2013 (.A0(net648),
    .A1(net188),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n984));
 sky130_fd_sc_hd__mux2_1 U2014 (.A0(net644),
    .A1(net189),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n985));
 sky130_fd_sc_hd__mux2_1 U2015 (.A0(net660),
    .A1(net113),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n982));
 sky130_fd_sc_hd__mux2_1 U2016 (.A0(net649),
    .A1(net114),
    .S(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n983));
 sky130_fd_sc_hd__nand2_8 U2017 (.A(n1460),
    .B(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1461));
 sky130_fd_sc_hd__mux2_1 U2018 (.A0(net648),
    .A1(net225),
    .S(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n992));
 sky130_fd_sc_hd__mux2_1 U2019 (.A0(net644),
    .A1(net226),
    .S(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n993));
 sky130_fd_sc_hd__mux2_1 U2020 (.A0(net662),
    .A1(net227),
    .S(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n990));
 sky130_fd_sc_hd__mux2_1 U2021 (.A0(net652),
    .A1(net228),
    .S(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n991));
 sky130_fd_sc_hd__nand2_2 U2022 (.A(n1463),
    .B(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(n1464));
 sky130_fd_sc_hd__mux2_1 U2023 (.A0(net648),
    .A1(net588),
    .S(n1464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n996));
 sky130_fd_sc_hd__mux2_1 U2024 (.A0(net644),
    .A1(net589),
    .S(n1464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n997));
 sky130_fd_sc_hd__mux2_1 U2025 (.A0(net663),
    .A1(net222),
    .S(n1464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n994));
 sky130_fd_sc_hd__mux2_1 U2026 (.A0(net652),
    .A1(net223),
    .S(n1464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n995));
 sky130_fd_sc_hd__a22o_1 U2027 (.A1(net606),
    .A2(net211),
    .B1(net614),
    .B2(net380),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1465));
 sky130_fd_sc_hd__a21o_1 U2028 (.A1(net615),
    .A2(net406),
    .B1(n1465),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net76));
 sky130_fd_sc_hd__a22o_1 U2029 (.A1(net606),
    .A2(net213),
    .B1(net614),
    .B2(net242),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(n1467));
 sky130_fd_sc_hd__a21o_1 U2030 (.A1(net615),
    .A2(net397),
    .B1(n1467),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net78));
 sky130_fd_sc_hd__a21o_1 U2033 (.A1(n1469),
    .A2(net195),
    .B1(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net80));
 sky130_fd_sc_hd__a21o_1 U2034 (.A1(n1469),
    .A2(net196),
    .B1(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net81));
 sky130_fd_sc_hd__a21o_1 U2035 (.A1(n1469),
    .A2(net197),
    .B1(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net82));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc0_in_REG_reg_0_ (.CLK(clknet_leaf_3_PCLK),
    .D(n718),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net95));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc0_in_REG_reg_1_ (.CLK(clknet_leaf_3_PCLK),
    .D(n719),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net94));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_adc0_in_REG_reg_2_ (.CLK(clknet_leaf_7_PCLK),
    .D(n720),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net102));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_adc0_in_REG_reg_3_ (.CLK(clknet_leaf_8_PCLK),
    .D(n721),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net101));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_adc0_in_REG_reg_4_ (.CLK(clknet_leaf_7_PCLK),
    .D(n722),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net100));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc0_in_REG_reg_5_ (.CLK(clknet_leaf_10_PCLK),
    .D(n723),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net103));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc0_in_REG_reg_6_ (.CLK(clknet_leaf_2_PCLK),
    .D(n724),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net98));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc0_in_REG_reg_7_ (.CLK(clknet_leaf_2_PCLK),
    .D(n725),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net99));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc0_in_REG_reg_8_ (.CLK(clknet_leaf_7_PCLK),
    .D(n726),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net96));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc0_in_REG_reg_9_ (.CLK(clknet_leaf_9_PCLK),
    .D(n727),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net97));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_adc1_in_REG_reg_0_ (.CLK(clknet_leaf_0_PCLK),
    .D(n709),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net105));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc1_in_REG_reg_1_ (.CLK(clknet_leaf_0_PCLK),
    .D(n710),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net104));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_adc1_in_REG_reg_2_ (.CLK(clknet_leaf_11_PCLK),
    .D(n711),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net111));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_adc1_in_REG_reg_3_ (.CLK(clknet_leaf_10_PCLK),
    .D(n712),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net110));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc1_in_REG_reg_4_ (.CLK(clknet_leaf_12_PCLK),
    .D(n713),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net112));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc1_in_REG_reg_5_ (.CLK(clknet_leaf_2_PCLK),
    .D(n714),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net108));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc1_in_REG_reg_6_ (.CLK(clknet_leaf_2_PCLK),
    .D(n715),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net109));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc1_in_REG_reg_7_ (.CLK(clknet_leaf_12_PCLK),
    .D(n716),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net106));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_adc1_in_REG_reg_8_ (.CLK(clknet_leaf_12_PCLK),
    .D(n717),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net107));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inn_REG_reg_0_ (.CLK(clknet_leaf_1_PCLK),
    .D(n824),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net329));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp0_inn_REG_reg_10_ (.CLK(clknet_leaf_11_PCLK),
    .D(n834),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net336));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inn_REG_reg_1_ (.CLK(clknet_leaf_2_PCLK),
    .D(n825),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net330));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp0_inn_REG_reg_2_ (.CLK(clknet_leaf_1_PCLK),
    .D(n826),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net328));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp0_inn_REG_reg_3_ (.CLK(clknet_leaf_1_PCLK),
    .D(n827),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net327));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp0_inn_REG_reg_4_ (.CLK(clknet_leaf_2_PCLK),
    .D(n828),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net326));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inn_REG_reg_5_ (.CLK(clknet_leaf_19_PCLK),
    .D(n829),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net331));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inn_REG_reg_6_ (.CLK(clknet_leaf_19_PCLK),
    .D(n830),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net332));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inn_REG_reg_7_ (.CLK(clknet_leaf_7_PCLK),
    .D(n831),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net334));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inn_REG_reg_8_ (.CLK(clknet_leaf_10_PCLK),
    .D(n832),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net335));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inn_REG_reg_9_ (.CLK(clknet_leaf_10_PCLK),
    .D(n833),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net333));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inp_REG_reg_0_ (.CLK(clknet_leaf_1_PCLK),
    .D(n835),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net340));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inp_REG_reg_1_ (.CLK(clknet_leaf_2_PCLK),
    .D(n836),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net341));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inp_REG_reg_2_ (.CLK(clknet_leaf_1_PCLK),
    .D(n837),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net339));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inp_REG_reg_3_ (.CLK(clknet_leaf_19_PCLK),
    .D(n838),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net338));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp0_inp_REG_reg_4_ (.CLK(clknet_leaf_0_PCLK),
    .D(n839),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net337));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp0_inp_REG_reg_5_ (.CLK(clknet_leaf_0_PCLK),
    .D(n840),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net343));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inp_REG_reg_6_ (.CLK(clknet_leaf_13_PCLK),
    .D(n841),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net344));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inp_REG_reg_7_ (.CLK(clknet_leaf_14_PCLK),
    .D(n842),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net342));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_inp_REG_reg_8_ (.CLK(clknet_leaf_14_PCLK),
    .D(n843),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net345));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_0_ (.CLK(clknet_leaf_3_PCLK),
    .D(n914),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net358));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_10_ (.CLK(clknet_leaf_1_PCLK),
    .D(n924),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net348));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_11_ (.CLK(clknet_leaf_0_PCLK),
    .D(n925),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net349));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_12_ (.CLK(clknet_leaf_14_PCLK),
    .D(n926),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net354));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_13_ (.CLK(clknet_leaf_14_PCLK),
    .D(n927),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net355));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_1_ (.CLK(clknet_leaf_4_PCLK),
    .D(n915),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net359));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_2_ (.CLK(clknet_leaf_1_PCLK),
    .D(n916),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net352));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_3_ (.CLK(clknet_leaf_0_PCLK),
    .D(n917),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net353));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_4_ (.CLK(clknet_leaf_3_PCLK),
    .D(n918),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net346));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_5_ (.CLK(clknet_leaf_3_PCLK),
    .D(n919),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net347));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_6_ (.CLK(clknet_leaf_3_PCLK),
    .D(n920),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net356));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_7_ (.CLK(clknet_leaf_3_PCLK),
    .D(n921),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net357));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_8_ (.CLK(clknet_leaf_3_PCLK),
    .D(n922),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net350));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp0_out_REG_reg_9_ (.CLK(clknet_leaf_1_PCLK),
    .D(n923),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net351));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_0_ (.CLK(clknet_leaf_2_PCLK),
    .D(n844),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net249));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp1_inn_REG_reg_10_ (.CLK(clknet_leaf_10_PCLK),
    .D(n854),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net256));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_11_ (.CLK(clknet_leaf_12_PCLK),
    .D(n855),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net247));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_12_ (.CLK(clknet_leaf_11_PCLK),
    .D(n856),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net248));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_1_ (.CLK(clknet_leaf_3_PCLK),
    .D(n845),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net250));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_2_ (.CLK(clknet_leaf_3_PCLK),
    .D(n846),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net246));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_3_ (.CLK(clknet_leaf_0_PCLK),
    .D(n847),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net245));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_4_ (.CLK(clknet_leaf_4_PCLK),
    .D(n848),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net244));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_5_ (.CLK(clknet_leaf_4_PCLK),
    .D(n849),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net251));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_6_ (.CLK(clknet_leaf_3_PCLK),
    .D(n850),
    .RESET_B(net672),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net252));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_7_ (.CLK(clknet_leaf_7_PCLK),
    .D(n851),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net254));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_8_ (.CLK(clknet_leaf_8_PCLK),
    .D(n852),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net255));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inn_REG_reg_9_ (.CLK(clknet_leaf_9_PCLK),
    .D(n853),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net253));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_0_ (.CLK(clknet_leaf_19_PCLK),
    .D(n857),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net262));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_10_ (.CLK(clknet_leaf_13_PCLK),
    .D(n867),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net260));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_11_ (.CLK(clknet_leaf_14_PCLK),
    .D(n868),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net261));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_1_ (.CLK(clknet_leaf_19_PCLK),
    .D(n858),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net263));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_2_ (.CLK(clknet_leaf_19_PCLK),
    .D(n859),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net259));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_3_ (.CLK(clknet_leaf_0_PCLK),
    .D(n860),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net258));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_4_ (.CLK(clknet_leaf_0_PCLK),
    .D(n861),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net257));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_5_ (.CLK(clknet_leaf_19_PCLK),
    .D(n862),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net265));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_6_ (.CLK(clknet_leaf_11_PCLK),
    .D(n863),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net266));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_inp_REG_reg_7_ (.CLK(clknet_leaf_11_PCLK),
    .D(n864),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net267));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp1_inp_REG_reg_8_ (.CLK(clknet_leaf_12_PCLK),
    .D(n865),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net264));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp1_inp_REG_reg_9_ (.CLK(clknet_leaf_12_PCLK),
    .D(n866),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net268));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp1_out_REG_reg_0_ (.CLK(clknet_leaf_3_PCLK),
    .D(n928),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net285));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_10_ (.CLK(clknet_leaf_1_PCLK),
    .D(n938),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net273));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_11_ (.CLK(clknet_leaf_19_PCLK),
    .D(n939),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net274));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_12_ (.CLK(clknet_leaf_19_PCLK),
    .D(n940),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net271));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_13_ (.CLK(clknet_leaf_19_PCLK),
    .D(n941),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net272));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp1_out_REG_reg_14_ (.CLK(clknet_leaf_12_PCLK),
    .D(n942),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net279));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp1_out_REG_reg_15_ (.CLK(clknet_leaf_10_PCLK),
    .D(n943),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net280));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp1_out_REG_reg_16_ (.CLK(clknet_leaf_12_PCLK),
    .D(n944),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net277));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp1_out_REG_reg_17_ (.CLK(clknet_leaf_12_PCLK),
    .D(n945),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net278));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp1_out_REG_reg_1_ (.CLK(clknet_leaf_4_PCLK),
    .D(n929),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net286));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_2_ (.CLK(clknet_leaf_1_PCLK),
    .D(n930),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net275));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_3_ (.CLK(clknet_leaf_4_PCLK),
    .D(n931),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net276));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_4_ (.CLK(clknet_leaf_4_PCLK),
    .D(n932),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net269));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp1_out_REG_reg_5_ (.CLK(clknet_leaf_3_PCLK),
    .D(n933),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net270));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_6_ (.CLK(clknet_leaf_2_PCLK),
    .D(n934),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net283));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_7_ (.CLK(clknet_leaf_3_PCLK),
    .D(n935),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net284));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_8_ (.CLK(clknet_leaf_1_PCLK),
    .D(n936),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net281));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp1_out_REG_reg_9_ (.CLK(clknet_leaf_1_PCLK),
    .D(n937),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net282));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_0_ (.CLK(clknet_leaf_11_PCLK),
    .D(n869),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net414));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_10_ (.CLK(clknet_leaf_12_PCLK),
    .D(n879),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net421));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_11_ (.CLK(clknet_leaf_13_PCLK),
    .D(n880),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net412));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_12_ (.CLK(clknet_leaf_13_PCLK),
    .D(n881),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net413));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_1_ (.CLK(clknet_leaf_11_PCLK),
    .D(n870),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net415));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_2_ (.CLK(clknet_leaf_10_PCLK),
    .D(n871),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net411));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_3_ (.CLK(clknet_leaf_10_PCLK),
    .D(n872),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net410));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_4_ (.CLK(clknet_leaf_12_PCLK),
    .D(n873),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net409));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_5_ (.CLK(clknet_leaf_13_PCLK),
    .D(n874),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net416));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_6_ (.CLK(clknet_leaf_13_PCLK),
    .D(n875),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net417));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_7_ (.CLK(clknet_leaf_13_PCLK),
    .D(n876),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net419));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_8_ (.CLK(clknet_leaf_13_PCLK),
    .D(n877),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net420));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inn_REG_reg_9_ (.CLK(clknet_leaf_13_PCLK),
    .D(n878),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net418));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_0_ (.CLK(clknet_leaf_7_PCLK),
    .D(n882),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net427));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_10_ (.CLK(clknet_leaf_9_PCLK),
    .D(n892),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net426));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_1_ (.CLK(clknet_leaf_7_PCLK),
    .D(n883),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net428));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_2_ (.CLK(clknet_leaf_8_PCLK),
    .D(n884),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net424));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_3_ (.CLK(clknet_leaf_8_PCLK),
    .D(n885),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net423));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_4_ (.CLK(clknet_leaf_9_PCLK),
    .D(n886),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net422));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_5_ (.CLK(clknet_leaf_8_PCLK),
    .D(n887),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net430));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp2_inp_REG_reg_6_ (.CLK(clknet_leaf_8_PCLK),
    .D(n888),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net431));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_7_ (.CLK(clknet_leaf_8_PCLK),
    .D(n889),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net429));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_8_ (.CLK(clknet_leaf_9_PCLK),
    .D(n890),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net432));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_inp_REG_reg_9_ (.CLK(clknet_leaf_9_PCLK),
    .D(n891),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net425));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_0_ (.CLK(clknet_leaf_19_PCLK),
    .D(n946),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net449));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp2_out_REG_reg_10_ (.CLK(clknet_leaf_13_PCLK),
    .D(n956),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net437));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_11_ (.CLK(clknet_leaf_13_PCLK),
    .D(n957),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net438));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_12_ (.CLK(clknet_leaf_13_PCLK),
    .D(n958),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net435));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_13_ (.CLK(clknet_leaf_13_PCLK),
    .D(n959),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net436));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp2_out_REG_reg_14_ (.CLK(clknet_leaf_13_PCLK),
    .D(n960),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net443));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_15_ (.CLK(clknet_leaf_13_PCLK),
    .D(n961),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net444));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_16_ (.CLK(clknet_leaf_13_PCLK),
    .D(n962),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net441));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp2_out_REG_reg_17_ (.CLK(clknet_leaf_12_PCLK),
    .D(n963),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net442));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_1_ (.CLK(clknet_leaf_19_PCLK),
    .D(n947),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net450));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_2_ (.CLK(clknet_leaf_19_PCLK),
    .D(n948),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net439));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_3_ (.CLK(clknet_leaf_19_PCLK),
    .D(n949),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net440));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_4_ (.CLK(clknet_leaf_19_PCLK),
    .D(n950),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net433));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_5_ (.CLK(clknet_leaf_18_PCLK),
    .D(n951),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net434));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_6_ (.CLK(clknet_leaf_19_PCLK),
    .D(n952),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net447));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_7_ (.CLK(clknet_leaf_1_PCLK),
    .D(n953),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net448));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_8_ (.CLK(clknet_leaf_19_PCLK),
    .D(n954),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net445));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp2_out_REG_reg_9_ (.CLK(clknet_leaf_19_PCLK),
    .D(n955),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net446));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_0_ (.CLK(clknet_leaf_8_PCLK),
    .D(n893),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net492));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_10_ (.CLK(clknet_leaf_10_PCLK),
    .D(n903),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net494));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_1_ (.CLK(clknet_leaf_7_PCLK),
    .D(n894),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net491));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_2_ (.CLK(clknet_leaf_9_PCLK),
    .D(n895),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net490));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_3_ (.CLK(clknet_leaf_9_PCLK),
    .D(n896),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net495));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_4_ (.CLK(clknet_leaf_8_PCLK),
    .D(n897),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net496));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_5_ (.CLK(clknet_leaf_8_PCLK),
    .D(n898),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net498));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp3_inn_REG_reg_6_ (.CLK(clknet_leaf_8_PCLK),
    .D(n899),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net499));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_7_ (.CLK(clknet_leaf_10_PCLK),
    .D(n900),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net497));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_8_ (.CLK(clknet_leaf_9_PCLK),
    .D(n901),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net500));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inn_REG_reg_9_ (.CLK(clknet_leaf_9_PCLK),
    .D(n902),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net493));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp3_inp_REG_reg_0_ (.CLK(clknet_leaf_12_PCLK),
    .D(n904),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net503));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inp_REG_reg_1_ (.CLK(clknet_leaf_12_PCLK),
    .D(n905),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net502));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp3_inp_REG_reg_2_ (.CLK(clknet_leaf_12_PCLK),
    .D(n906),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net501));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp3_inp_REG_reg_3_ (.CLK(clknet_leaf_11_PCLK),
    .D(n907),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net507));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp3_inp_REG_reg_4_ (.CLK(clknet_leaf_13_PCLK),
    .D(n908),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net508));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inp_REG_reg_5_ (.CLK(clknet_leaf_13_PCLK),
    .D(n909),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net509));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp3_inp_REG_reg_6_ (.CLK(clknet_leaf_13_PCLK),
    .D(n910),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net506));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_amp3_inp_REG_reg_7_ (.CLK(clknet_leaf_13_PCLK),
    .D(n911),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net510));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inp_REG_reg_8_ (.CLK(clknet_leaf_13_PCLK),
    .D(n912),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net504));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_inp_REG_reg_9_ (.CLK(clknet_leaf_13_PCLK),
    .D(n913),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net505));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_0_ (.CLK(clknet_leaf_19_PCLK),
    .D(n964),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net527));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_10_ (.CLK(clknet_leaf_9_PCLK),
    .D(n974),
    .RESET_B(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net515));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_11_ (.CLK(clknet_leaf_12_PCLK),
    .D(n975),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net516));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_12_ (.CLK(clknet_leaf_14_PCLK),
    .D(n976),
    .RESET_B(net694),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net513));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp3_out_REG_reg_13_ (.CLK(clknet_leaf_14_PCLK),
    .D(n977),
    .RESET_B(net695),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net514));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_14_ (.CLK(clknet_leaf_13_PCLK),
    .D(n978),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net521));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp3_out_REG_reg_15_ (.CLK(clknet_leaf_12_PCLK),
    .D(n979),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net522));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_amp3_out_REG_reg_16_ (.CLK(clknet_leaf_13_PCLK),
    .D(n980),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net519));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_17_ (.CLK(clknet_leaf_12_PCLK),
    .D(n981),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net520));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_1_ (.CLK(clknet_leaf_3_PCLK),
    .D(n965),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net528));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_2_ (.CLK(clknet_leaf_2_PCLK),
    .D(n966),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net517));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_3_ (.CLK(clknet_leaf_19_PCLK),
    .D(n967),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net518));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_4_ (.CLK(clknet_leaf_2_PCLK),
    .D(n968),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net511));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_5_ (.CLK(clknet_leaf_3_PCLK),
    .D(n969),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net512));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_6_ (.CLK(clknet_leaf_2_PCLK),
    .D(n970),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net525));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_7_ (.CLK(clknet_leaf_2_PCLK),
    .D(n971),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net526));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_8_ (.CLK(clknet_leaf_2_PCLK),
    .D(n972),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net523));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_amp3_out_REG_reg_9_ (.CLK(clknet_leaf_1_PCLK),
    .D(n973),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net524));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_0_ (.CLK(clknet_leaf_11_PCLK),
    .D(n728),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net158));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_1_ (.CLK(clknet_leaf_10_PCLK),
    .D(n729),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net157));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_2_ (.CLK(clknet_leaf_7_PCLK),
    .D(n730),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net164));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_3_ (.CLK(clknet_leaf_7_PCLK),
    .D(n731),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net165));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_4_ (.CLK(clknet_leaf_11_PCLK),
    .D(n732),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net163));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_5_ (.CLK(clknet_leaf_11_PCLK),
    .D(n733),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net166));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_6_ (.CLK(clknet_leaf_6_PCLK),
    .D(n734),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net161));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_7_ (.CLK(clknet_leaf_6_PCLK),
    .D(n735),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net162));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_8_ (.CLK(clknet_leaf_7_PCLK),
    .D(n736),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net159));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inn_REG_reg_9_ (.CLK(clknet_leaf_11_PCLK),
    .D(n737),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net160));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_comp0_inp_REG_reg_0_ (.CLK(clknet_leaf_10_PCLK),
    .D(n738),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net168));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inp_REG_reg_10_ (.CLK(clknet_leaf_12_PCLK),
    .D(n748),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net170));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp0_inp_REG_reg_1_ (.CLK(clknet_leaf_14_PCLK),
    .D(n739),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net167));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inp_REG_reg_2_ (.CLK(clknet_leaf_14_PCLK),
    .D(n740),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net174));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inp_REG_reg_3_ (.CLK(clknet_leaf_14_PCLK),
    .D(n741),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net176));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp0_inp_REG_reg_4_ (.CLK(clknet_leaf_14_PCLK),
    .D(n742),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net175));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp0_inp_REG_reg_5_ (.CLK(clknet_leaf_13_PCLK),
    .D(n743),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net173));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inp_REG_reg_6_ (.CLK(clknet_leaf_14_PCLK),
    .D(n744),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net177));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inp_REG_reg_7_ (.CLK(clknet_leaf_1_PCLK),
    .D(n745),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net171));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inp_REG_reg_8_ (.CLK(clknet_leaf_2_PCLK),
    .D(n746),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net172));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp0_inp_REG_reg_9_ (.CLK(clknet_leaf_12_PCLK),
    .D(n747),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net169));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_comp1_inn_REG_reg_0_ (.CLK(clknet_leaf_7_PCLK),
    .D(n749),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net556));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inn_REG_reg_1_ (.CLK(clknet_leaf_10_PCLK),
    .D(n750),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net555));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp1_inn_REG_reg_2_ (.CLK(clknet_leaf_10_PCLK),
    .D(n751),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net562));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp1_inn_REG_reg_3_ (.CLK(clknet_leaf_9_PCLK),
    .D(n752),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net563));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_comp1_inn_REG_reg_4_ (.CLK(clknet_leaf_9_PCLK),
    .D(n753),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net561));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp1_inn_REG_reg_5_ (.CLK(clknet_leaf_7_PCLK),
    .D(n754),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net564));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inn_REG_reg_6_ (.CLK(clknet_leaf_5_PCLK),
    .D(n755),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net559));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inn_REG_reg_7_ (.CLK(clknet_leaf_5_PCLK),
    .D(n756),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net560));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inn_REG_reg_8_ (.CLK(clknet_leaf_7_PCLK),
    .D(n757),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net557));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inn_REG_reg_9_ (.CLK(clknet_leaf_9_PCLK),
    .D(n758),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net558));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_comp1_inp_REG_reg_0_ (.CLK(clknet_leaf_7_PCLK),
    .D(n759),
    .RESET_B(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net566));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_10_ (.CLK(clknet_leaf_10_PCLK),
    .D(n769),
    .RESET_B(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net568));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_1_ (.CLK(clknet_leaf_7_PCLK),
    .D(n760),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net565));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp1_inp_REG_reg_2_ (.CLK(clknet_leaf_7_PCLK),
    .D(n761),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net572));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_comp1_inp_REG_reg_3_ (.CLK(clknet_leaf_7_PCLK),
    .D(n762),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net574));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_4_ (.CLK(clknet_leaf_7_PCLK),
    .D(n763),
    .RESET_B(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net573));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_5_ (.CLK(clknet_leaf_10_PCLK),
    .D(n764),
    .RESET_B(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net571));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_6_ (.CLK(clknet_leaf_7_PCLK),
    .D(n765),
    .RESET_B(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net575));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_7_ (.CLK(clknet_leaf_6_PCLK),
    .D(n766),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net569));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_8_ (.CLK(clknet_leaf_6_PCLK),
    .D(n767),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net570));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_comp1_inp_REG_reg_9_ (.CLK(clknet_leaf_7_PCLK),
    .D(n768),
    .RESET_B(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net567));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_dac_out_REG_reg_0_ (.CLK(clknet_leaf_0_PCLK),
    .D(n674),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net184));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_dac_out_REG_reg_1_ (.CLK(clknet_leaf_0_PCLK),
    .D(n675),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net186));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_dac_out_REG_reg_2_ (.CLK(clknet_leaf_4_PCLK),
    .D(n676),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net121));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_dac_out_REG_reg_3_ (.CLK(clknet_leaf_3_PCLK),
    .D(n677),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net122));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_dac_out_REG_reg_4_ (.CLK(clknet_leaf_4_PCLK),
    .D(n678),
    .RESET_B(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net123));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_dac_out_REG_reg_5_ (.CLK(clknet_leaf_1_PCLK),
    .D(n679),
    .RESET_B(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net124));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_idac_REG_reg_0_ (.CLK(clknet_leaf_8_PCLK),
    .D(n990),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net227));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_idac_REG_reg_1_ (.CLK(clknet_leaf_8_PCLK),
    .D(n991),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net228));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_idac_REG_reg_2_ (.CLK(clknet_leaf_8_PCLK),
    .D(n992),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net225));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_idac_REG_reg_3_ (.CLK(clknet_leaf_8_PCLK),
    .D(n993),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net226));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inn_REG_reg_0_ (.CLK(clknet_leaf_2_PCLK),
    .D(n793),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net300));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inn_REG_reg_1_ (.CLK(clknet_leaf_3_PCLK),
    .D(n794),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net301));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inn_REG_reg_2_ (.CLK(clknet_leaf_2_PCLK),
    .D(n795),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net299));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inn_REG_reg_3_ (.CLK(clknet_leaf_3_PCLK),
    .D(n796),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net298));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inn_REG_reg_4_ (.CLK(clknet_leaf_10_PCLK),
    .D(n797),
    .RESET_B(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net303));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inn_REG_reg_5_ (.CLK(clknet_leaf_11_PCLK),
    .D(n798),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net302));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_preamp0_inn_REG_reg_6_ (.CLK(clknet_leaf_10_PCLK),
    .D(n799),
    .RESET_B(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net304));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inp_REG_reg_0_ (.CLK(clknet_leaf_2_PCLK),
    .D(n785),
    .RESET_B(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net307));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inp_REG_reg_1_ (.CLK(clknet_leaf_1_PCLK),
    .D(n786),
    .RESET_B(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net308));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inp_REG_reg_2_ (.CLK(clknet_leaf_19_PCLK),
    .D(n787),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net306));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inp_REG_reg_3_ (.CLK(clknet_leaf_19_PCLK),
    .D(n788),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net305));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inp_REG_reg_4_ (.CLK(clknet_leaf_14_PCLK),
    .D(n789),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net310));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_preamp0_inp_REG_reg_5_ (.CLK(clknet_leaf_14_PCLK),
    .D(n790),
    .RESET_B(net691),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net311));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_preamp0_inp_REG_reg_6_ (.CLK(clknet_leaf_14_PCLK),
    .D(n791),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net309));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_inp_REG_reg_7_ (.CLK(clknet_leaf_12_PCLK),
    .D(n792),
    .RESET_B(net692),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net312));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_0_ (.CLK(clknet_leaf_1_PCLK),
    .D(n812),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net323));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_10_ (.CLK(clknet_leaf_1_PCLK),
    .D(n822),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net315));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_11_ (.CLK(clknet_leaf_19_PCLK),
    .D(n823),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net316));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_preamp0_out_REG_reg_1_ (.CLK(clknet_leaf_3_PCLK),
    .D(n813),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net324));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_2_ (.CLK(clknet_leaf_2_PCLK),
    .D(n814),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net319));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_3_ (.CLK(clknet_leaf_2_PCLK),
    .D(n815),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net320));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_4_ (.CLK(clknet_leaf_1_PCLK),
    .D(n816),
    .RESET_B(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net313));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_preamp0_out_REG_reg_5_ (.CLK(clknet_leaf_2_PCLK),
    .D(n817),
    .RESET_B(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net314));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_6_ (.CLK(clknet_leaf_2_PCLK),
    .D(n818),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net321));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_7_ (.CLK(clknet_leaf_2_PCLK),
    .D(n819),
    .RESET_B(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net322));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_8_ (.CLK(clknet_leaf_1_PCLK),
    .D(n820),
    .RESET_B(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net317));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp0_out_REG_reg_9_ (.CLK(clknet_leaf_1_PCLK),
    .D(n821),
    .RESET_B(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net318));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inn_REG_reg_0_ (.CLK(clknet_leaf_8_PCLK),
    .D(n778),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net463));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inn_REG_reg_1_ (.CLK(clknet_leaf_8_PCLK),
    .D(n779),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net462));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inn_REG_reg_2_ (.CLK(clknet_leaf_9_PCLK),
    .D(n780),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net467));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inn_REG_reg_3_ (.CLK(clknet_leaf_8_PCLK),
    .D(n781),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net466));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inn_REG_reg_4_ (.CLK(clknet_leaf_9_PCLK),
    .D(n782),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net468));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inn_REG_reg_5_ (.CLK(clknet_leaf_9_PCLK),
    .D(n783),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net464));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inn_REG_reg_6_ (.CLK(clknet_leaf_8_PCLK),
    .D(n784),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net465));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_0_ (.CLK(clknet_leaf_10_PCLK),
    .D(n770),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net470));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_1_ (.CLK(clknet_leaf_9_PCLK),
    .D(n771),
    .RESET_B(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net469));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_2_ (.CLK(clknet_leaf_10_PCLK),
    .D(n772),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net474));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_3_ (.CLK(clknet_leaf_9_PCLK),
    .D(n773),
    .RESET_B(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net475));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_4_ (.CLK(clknet_leaf_10_PCLK),
    .D(n774),
    .RESET_B(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net473));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_5_ (.CLK(clknet_leaf_12_PCLK),
    .D(n775),
    .RESET_B(net700),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net476));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_6_ (.CLK(clknet_leaf_9_PCLK),
    .D(n776),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net471));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_inp_REG_reg_7_ (.CLK(clknet_leaf_9_PCLK),
    .D(n777),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net472));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_preamp1_out_REG_reg_0_ (.CLK(clknet_leaf_3_PCLK),
    .D(n800),
    .RESET_B(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net487));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_out_REG_reg_10_ (.CLK(clknet_leaf_12_PCLK),
    .D(n810),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net485));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_out_REG_reg_11_ (.CLK(clknet_leaf_12_PCLK),
    .D(n811),
    .RESET_B(net697),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net486));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_preamp1_out_REG_reg_1_ (.CLK(clknet_leaf_3_PCLK),
    .D(n801),
    .RESET_B(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net488));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_preamp1_out_REG_reg_2_ (.CLK(clknet_leaf_1_PCLK),
    .D(n802),
    .RESET_B(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net483));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_preamp1_out_REG_reg_3_ (.CLK(clknet_leaf_1_PCLK),
    .D(n803),
    .RESET_B(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net484));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_out_REG_reg_4_ (.CLK(clknet_leaf_1_PCLK),
    .D(n804),
    .RESET_B(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net477));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_preamp1_out_REG_reg_5_ (.CLK(clknet_leaf_3_PCLK),
    .D(n805),
    .RESET_B(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net478));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_out_REG_reg_6_ (.CLK(clknet_leaf_8_PCLK),
    .D(n806),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net481));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_out_REG_reg_7_ (.CLK(clknet_leaf_8_PCLK),
    .D(n807),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net482));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_out_REG_reg_8_ (.CLK(clknet_leaf_12_PCLK),
    .D(n808),
    .RESET_B(net698),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net479));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_preamp1_out_REG_reg_9_ (.CLK(clknet_leaf_10_PCLK),
    .D(n809),
    .RESET_B(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net480));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_0_ (.CLK(clknet_leaf_3_PCLK),
    .D(n982),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net113));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_1_ (.CLK(clknet_leaf_2_PCLK),
    .D(n983),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net114));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_2_ (.CLK(clknet_leaf_8_PCLK),
    .D(n984),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net188));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_3_ (.CLK(clknet_leaf_8_PCLK),
    .D(n985),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net189));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_4_ (.CLK(clknet_leaf_2_PCLK),
    .D(n986),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net115));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_5_ (.CLK(clknet_leaf_3_PCLK),
    .D(n987),
    .RESET_B(net664),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net116));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_6_ (.CLK(clknet_leaf_8_PCLK),
    .D(n988),
    .RESET_B(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net190));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_ref_REG_reg_7_ (.CLK(clknet_leaf_8_PCLK),
    .D(n989),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net191));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_sio_ana_REG_reg_0_ (.CLK(clknet_leaf_17_PCLK),
    .D(n701),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net117));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_sio_ana_REG_reg_1_ (.CLK(clknet_leaf_16_PCLK),
    .D(n702),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net118));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_sio_ana_REG_reg_2_ (.CLK(clknet_leaf_17_PCLK),
    .D(n703),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net119));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_sio_ana_REG_reg_3_ (.CLK(clknet_leaf_17_PCLK),
    .D(n704),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net120));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_sio_iso_REG_reg_0_ (.CLK(clknet_leaf_11_PCLK),
    .D(n705),
    .RESET_B(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net546));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_sio_iso_REG_reg_1_ (.CLK(clknet_leaf_11_PCLK),
    .D(n706),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net547));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_sio_iso_REG_reg_2_ (.CLK(clknet_leaf_11_PCLK),
    .D(n707),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net548));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_sio_iso_REG_reg_3_ (.CLK(clknet_leaf_14_PCLK),
    .D(n708),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net549));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_test_REG_reg_0_ (.CLK(clknet_leaf_9_PCLK),
    .D(n994),
    .RESET_B(net701),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net222));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_test_REG_reg_1_ (.CLK(clknet_leaf_9_PCLK),
    .D(n995),
    .RESET_B(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net223));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_test_REG_reg_2_ (.CLK(clknet_leaf_9_PCLK),
    .D(n996),
    .RESET_B(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net588));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_test_REG_reg_3_ (.CLK(clknet_leaf_9_PCLK),
    .D(n997),
    .RESET_B(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net589));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_0_ (.CLK(clknet_leaf_7_PCLK),
    .D(n680),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net591));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_10_ (.CLK(clknet_leaf_11_PCLK),
    .D(n690),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net576));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_uproj_REG_reg_11_ (.CLK(clknet_leaf_14_PCLK),
    .D(n691),
    .RESET_B(net689),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net577));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_uproj_REG_reg_12_ (.CLK(clknet_leaf_14_PCLK),
    .D(n692),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net578));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_uproj_REG_reg_13_ (.CLK(clknet_leaf_14_PCLK),
    .D(n693),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net579));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_uproj_REG_reg_14_ (.CLK(clknet_leaf_14_PCLK),
    .D(n694),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net185));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_uproj_REG_reg_15_ (.CLK(clknet_leaf_15_PCLK),
    .D(n695),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net187));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_uproj_REG_reg_16_ (.CLK(clknet_leaf_14_PCLK),
    .D(n696),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net552));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_uproj_REG_reg_17_ (.CLK(clknet_leaf_14_PCLK),
    .D(n697),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net545));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_uproj_REG_reg_18_ (.CLK(clknet_leaf_15_PCLK),
    .D(n698),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net376));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_uproj_REG_reg_19_ (.CLK(clknet_leaf_15_PCLK),
    .D(n699),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net592));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_1_ (.CLK(clknet_leaf_10_PCLK),
    .D(n681),
    .RESET_B(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net590));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_uproj_REG_reg_20_ (.CLK(clknet_leaf_15_PCLK),
    .D(n700),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net593));
 sky130_fd_sc_hd__dfrtp_2 reg_ana_uproj_REG_reg_2_ (.CLK(clknet_leaf_14_PCLK),
    .D(n682),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net580));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_3_ (.CLK(clknet_leaf_11_PCLK),
    .D(n683),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net581));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_4_ (.CLK(clknet_leaf_7_PCLK),
    .D(n684),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net582));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_5_ (.CLK(clknet_leaf_7_PCLK),
    .D(n685),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net583));
 sky130_fd_sc_hd__dfrtp_4 reg_ana_uproj_REG_reg_6_ (.CLK(clknet_leaf_14_PCLK),
    .D(n686),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net584));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_7_ (.CLK(clknet_leaf_11_PCLK),
    .D(n687),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net585));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_8_ (.CLK(clknet_leaf_11_PCLK),
    .D(n688),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net586));
 sky130_fd_sc_hd__dfrtp_1 reg_ana_uproj_REG_reg_9_ (.CLK(clknet_leaf_11_PCLK),
    .D(n689),
    .RESET_B(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net587));
 sky130_fd_sc_hd__dfstp_1 reg_bandgap_ctrl_REG_reg_0_ (.CLK(clknet_leaf_16_PCLK),
    .D(n498),
    .SET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net125));
 sky130_fd_sc_hd__dfrtp_1 reg_bandgap_ctrl_REG_reg_10_ (.CLK(clknet_leaf_5_PCLK),
    .D(n591),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net142));
 sky130_fd_sc_hd__dfrtp_2 reg_bandgap_ctrl_REG_reg_11_ (.CLK(clknet_leaf_16_PCLK),
    .D(n592),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net128));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_12_ (.CLK(clknet_leaf_16_PCLK),
    .D(n593),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net129));
 sky130_fd_sc_hd__dfrtp_2 reg_bandgap_ctrl_REG_reg_13_ (.CLK(clknet_leaf_17_PCLK),
    .D(n594),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net130));
 sky130_fd_sc_hd__dfrtp_2 reg_bandgap_ctrl_REG_reg_14_ (.CLK(clknet_leaf_17_PCLK),
    .D(n595),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net131));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_15_ (.CLK(clknet_leaf_16_PCLK),
    .D(n596),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net132));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_16_ (.CLK(clknet_leaf_17_PCLK),
    .D(n597),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net133));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_17_ (.CLK(clknet_leaf_17_PCLK),
    .D(n598),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net126));
 sky130_fd_sc_hd__dfstp_1 reg_bandgap_ctrl_REG_reg_18_ (.CLK(clknet_leaf_17_PCLK),
    .D(n499),
    .SET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net241));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_19_ (.CLK(clknet_leaf_15_PCLK),
    .D(n599),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net377));
 sky130_fd_sc_hd__dfrtp_2 reg_bandgap_ctrl_REG_reg_1_ (.CLK(clknet_leaf_5_PCLK),
    .D(n582),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net127));
 sky130_fd_sc_hd__dfrtp_2 reg_bandgap_ctrl_REG_reg_20_ (.CLK(clknet_leaf_15_PCLK),
    .D(n600),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net378));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_21_ (.CLK(clknet_leaf_18_PCLK),
    .D(n601),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net379));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_22_ (.CLK(clknet_leaf_18_PCLK),
    .D(n602),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net380));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_23_ (.CLK(clknet_leaf_18_PCLK),
    .D(n603),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net381));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_24_ (.CLK(clknet_leaf_18_PCLK),
    .D(n604),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net242));
 sky130_fd_sc_hd__dfrtp_1 reg_bandgap_ctrl_REG_reg_2_ (.CLK(clknet_leaf_5_PCLK),
    .D(n583),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net134));
 sky130_fd_sc_hd__dfrtp_2 reg_bandgap_ctrl_REG_reg_3_ (.CLK(clknet_leaf_17_PCLK),
    .D(n584),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net135));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_4_ (.CLK(clknet_leaf_6_PCLK),
    .D(n585),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net136));
 sky130_fd_sc_hd__dfrtp_1 reg_bandgap_ctrl_REG_reg_5_ (.CLK(clknet_leaf_5_PCLK),
    .D(n586),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net137));
 sky130_fd_sc_hd__dfrtp_2 reg_bandgap_ctrl_REG_reg_6_ (.CLK(clknet_leaf_17_PCLK),
    .D(n587),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net138));
 sky130_fd_sc_hd__dfrtp_1 reg_bandgap_ctrl_REG_reg_7_ (.CLK(clknet_leaf_6_PCLK),
    .D(n588),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net139));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_8_ (.CLK(clknet_leaf_6_PCLK),
    .D(n589),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net140));
 sky130_fd_sc_hd__dfrtp_4 reg_bandgap_ctrl_REG_reg_9_ (.CLK(clknet_leaf_6_PCLK),
    .D(n590),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net141));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_0_ (.CLK(clknet_leaf_4_PCLK),
    .D(n500),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net143));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_10_ (.CLK(clknet_leaf_0_PCLK),
    .D(n510),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net149));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_1_ (.CLK(clknet_leaf_4_PCLK),
    .D(n501),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net151));
 sky130_fd_sc_hd__dfrtp_1 reg_brownout_ctrl_REG_reg_2_ (.CLK(clknet_leaf_5_PCLK),
    .D(n502),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net152));
 sky130_fd_sc_hd__dfrtp_1 reg_brownout_ctrl_REG_reg_3_ (.CLK(clknet_leaf_4_PCLK),
    .D(n503),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net153));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_4_ (.CLK(clknet_leaf_4_PCLK),
    .D(n504),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net146));
 sky130_fd_sc_hd__dfrtp_1 reg_brownout_ctrl_REG_reg_5_ (.CLK(clknet_leaf_5_PCLK),
    .D(n505),
    .RESET_B(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net147));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_6_ (.CLK(clknet_leaf_5_PCLK),
    .D(n506),
    .RESET_B(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net148));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_7_ (.CLK(clknet_leaf_5_PCLK),
    .D(n507),
    .RESET_B(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net144));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_8_ (.CLK(clknet_leaf_5_PCLK),
    .D(n508),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net145));
 sky130_fd_sc_hd__dfrtp_4 reg_brownout_ctrl_REG_reg_9_ (.CLK(clknet_leaf_4_PCLK),
    .D(n509),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net150));
 sky130_fd_sc_hd__dfrtp_1 reg_comparator_ctrl_REG_reg_0_ (.CLK(clknet_leaf_5_PCLK),
    .D(n605),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net154));
 sky130_fd_sc_hd__dfrtp_4 reg_comparator_ctrl_REG_reg_10_ (.CLK(clknet_leaf_5_PCLK),
    .D(n615),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net553));
 sky130_fd_sc_hd__dfrtp_2 reg_comparator_ctrl_REG_reg_1_ (.CLK(clknet_leaf_17_PCLK),
    .D(n606),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net178));
 sky130_fd_sc_hd__dfrtp_1 reg_comparator_ctrl_REG_reg_2_ (.CLK(clknet_leaf_16_PCLK),
    .D(n607),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net179));
 sky130_fd_sc_hd__dfrtp_1 reg_comparator_ctrl_REG_reg_3_ (.CLK(clknet_leaf_5_PCLK),
    .D(n608),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net180));
 sky130_fd_sc_hd__dfrtp_4 reg_comparator_ctrl_REG_reg_4_ (.CLK(clknet_leaf_5_PCLK),
    .D(n609),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net181));
 sky130_fd_sc_hd__dfrtp_4 reg_comparator_ctrl_REG_reg_5_ (.CLK(clknet_leaf_16_PCLK),
    .D(n610),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net182));
 sky130_fd_sc_hd__dfrtp_1 reg_comparator_ctrl_REG_reg_6_ (.CLK(clknet_leaf_16_PCLK),
    .D(n611),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net183));
 sky130_fd_sc_hd__dfrtp_1 reg_comparator_ctrl_REG_reg_7_ (.CLK(clknet_leaf_5_PCLK),
    .D(n612),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net155));
 sky130_fd_sc_hd__dfrtp_1 reg_comparator_ctrl_REG_reg_8_ (.CLK(clknet_leaf_5_PCLK),
    .D(n613),
    .RESET_B(net679),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net156));
 sky130_fd_sc_hd__dfrtp_4 reg_comparator_ctrl_REG_reg_9_ (.CLK(clknet_leaf_16_PCLK),
    .D(n614),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net554));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_0_ (.CLK(clknet_leaf_17_PCLK),
    .D(n552),
    .RESET_B(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net192));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_10_ (.CLK(clknet_leaf_6_PCLK),
    .D(n562),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net221));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_11_ (.CLK(clknet_leaf_16_PCLK),
    .D(n563),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net199));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_12_ (.CLK(clknet_leaf_16_PCLK),
    .D(n564),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net200));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_13_ (.CLK(clknet_leaf_16_PCLK),
    .D(n565),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net201));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_14_ (.CLK(clknet_leaf_15_PCLK),
    .D(n566),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net202));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_15_ (.CLK(clknet_leaf_5_PCLK),
    .D(n567),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net203));
 sky130_fd_sc_hd__dfrtp_2 reg_ibias_ctrl_REG_reg_16_ (.CLK(clknet_leaf_15_PCLK),
    .D(n568),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net204));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_17_ (.CLK(clknet_leaf_16_PCLK),
    .D(n569),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net205));
 sky130_fd_sc_hd__dfrtp_2 reg_ibias_ctrl_REG_reg_18_ (.CLK(clknet_leaf_15_PCLK),
    .D(n570),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net206));
 sky130_fd_sc_hd__dfrtp_2 reg_ibias_ctrl_REG_reg_19_ (.CLK(clknet_leaf_15_PCLK),
    .D(n571),
    .RESET_B(net683),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net207));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_1_ (.CLK(clknet_leaf_6_PCLK),
    .D(n553),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net198));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_20_ (.CLK(clknet_leaf_18_PCLK),
    .D(n572),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net208));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_21_ (.CLK(clknet_leaf_18_PCLK),
    .D(n573),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net210));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_22_ (.CLK(clknet_leaf_19_PCLK),
    .D(n574),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net211));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_23_ (.CLK(clknet_leaf_18_PCLK),
    .D(n575),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net212));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_24_ (.CLK(clknet_leaf_18_PCLK),
    .D(n576),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net213));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_25_ (.CLK(clknet_leaf_18_PCLK),
    .D(n577),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net194));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_26_ (.CLK(clknet_leaf_18_PCLK),
    .D(n578),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net195));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_27_ (.CLK(clknet_leaf_18_PCLK),
    .D(n579),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net196));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_28_ (.CLK(clknet_leaf_19_PCLK),
    .D(n580),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net197));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_29_ (.CLK(clknet_leaf_18_PCLK),
    .D(n581),
    .RESET_B(net665),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net193));
 sky130_fd_sc_hd__dfrtp_2 reg_ibias_ctrl_REG_reg_2_ (.CLK(clknet_leaf_5_PCLK),
    .D(n554),
    .RESET_B(net680),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net209));
 sky130_fd_sc_hd__dfrtp_2 reg_ibias_ctrl_REG_reg_3_ (.CLK(clknet_leaf_6_PCLK),
    .D(n555),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net214));
 sky130_fd_sc_hd__dfrtp_4 reg_ibias_ctrl_REG_reg_4_ (.CLK(clknet_leaf_18_PCLK),
    .D(n556),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net215));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_5_ (.CLK(clknet_leaf_15_PCLK),
    .D(n557),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net216));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_6_ (.CLK(clknet_leaf_6_PCLK),
    .D(n558),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net217));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_7_ (.CLK(clknet_leaf_6_PCLK),
    .D(n559),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net218));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_8_ (.CLK(clknet_leaf_6_PCLK),
    .D(n560),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net219));
 sky130_fd_sc_hd__dfrtp_1 reg_ibias_ctrl_REG_reg_9_ (.CLK(clknet_leaf_16_PCLK),
    .D(n561),
    .RESET_B(net684),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net220));
 sky130_fd_sc_hd__dfrtp_4 reg_idac_ctrl_REG_reg_0_ (.CLK(clknet_leaf_16_PCLK),
    .D(n539),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net229));
 sky130_fd_sc_hd__dfrtp_4 reg_idac_ctrl_REG_reg_10_ (.CLK(clknet_leaf_15_PCLK),
    .D(n549),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net230));
 sky130_fd_sc_hd__dfrtp_1 reg_idac_ctrl_REG_reg_11_ (.CLK(clknet_leaf_16_PCLK),
    .D(n550),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net231));
 sky130_fd_sc_hd__dfrtp_1 reg_idac_ctrl_REG_reg_12_ (.CLK(clknet_leaf_16_PCLK),
    .D(n551),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net224));
 sky130_fd_sc_hd__dfrtp_4 reg_idac_ctrl_REG_reg_1_ (.CLK(clknet_leaf_6_PCLK),
    .D(n540),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net232));
 sky130_fd_sc_hd__dfrtp_4 reg_idac_ctrl_REG_reg_2_ (.CLK(clknet_leaf_15_PCLK),
    .D(n541),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net233));
 sky130_fd_sc_hd__dfrtp_4 reg_idac_ctrl_REG_reg_3_ (.CLK(clknet_leaf_6_PCLK),
    .D(n542),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net234));
 sky130_fd_sc_hd__dfrtp_4 reg_idac_ctrl_REG_reg_4_ (.CLK(clknet_leaf_15_PCLK),
    .D(n543),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net235));
 sky130_fd_sc_hd__dfrtp_4 reg_idac_ctrl_REG_reg_5_ (.CLK(clknet_leaf_6_PCLK),
    .D(n544),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net236));
 sky130_fd_sc_hd__dfrtp_1 reg_idac_ctrl_REG_reg_6_ (.CLK(clknet_leaf_6_PCLK),
    .D(n545),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net237));
 sky130_fd_sc_hd__dfrtp_1 reg_idac_ctrl_REG_reg_7_ (.CLK(clknet_leaf_6_PCLK),
    .D(n546),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net238));
 sky130_fd_sc_hd__dfrtp_1 reg_idac_ctrl_REG_reg_8_ (.CLK(clknet_leaf_6_PCLK),
    .D(n547),
    .RESET_B(net685),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net239));
 sky130_fd_sc_hd__dfrtp_2 reg_idac_ctrl_REG_reg_9_ (.CLK(clknet_leaf_15_PCLK),
    .D(n548),
    .RESET_B(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net240));
 sky130_fd_sc_hd__dfrtp_1 reg_left_instramp_ctrl_REG_reg_0_ (.CLK(clknet_leaf_4_PCLK),
    .D(n663),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net297));
 sky130_fd_sc_hd__dfrtp_4 reg_left_instramp_ctrl_REG_reg_10_ (.CLK(clknet_leaf_0_PCLK),
    .D(n673),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net296));
 sky130_fd_sc_hd__dfrtp_1 reg_left_instramp_ctrl_REG_reg_1_ (.CLK(clknet_leaf_4_PCLK),
    .D(n664),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net287));
 sky130_fd_sc_hd__dfrtp_1 reg_left_instramp_ctrl_REG_reg_2_ (.CLK(clknet_leaf_5_PCLK),
    .D(n665),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net288));
 sky130_fd_sc_hd__dfrtp_1 reg_left_instramp_ctrl_REG_reg_3_ (.CLK(clknet_leaf_4_PCLK),
    .D(n666),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net289));
 sky130_fd_sc_hd__dfrtp_1 reg_left_instramp_ctrl_REG_reg_4_ (.CLK(clknet_leaf_5_PCLK),
    .D(n667),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net290));
 sky130_fd_sc_hd__dfrtp_1 reg_left_instramp_ctrl_REG_reg_5_ (.CLK(clknet_leaf_4_PCLK),
    .D(n668),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net291));
 sky130_fd_sc_hd__dfrtp_4 reg_left_instramp_ctrl_REG_reg_6_ (.CLK(clknet_leaf_4_PCLK),
    .D(n669),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net292));
 sky130_fd_sc_hd__dfrtp_4 reg_left_instramp_ctrl_REG_reg_7_ (.CLK(clknet_leaf_4_PCLK),
    .D(n670),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net293));
 sky130_fd_sc_hd__dfrtp_4 reg_left_instramp_ctrl_REG_reg_8_ (.CLK(clknet_leaf_5_PCLK),
    .D(n671),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net294));
 sky130_fd_sc_hd__dfrtp_4 reg_left_instramp_ctrl_REG_reg_9_ (.CLK(clknet_leaf_0_PCLK),
    .D(n672),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net295));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_0_ (.CLK(clknet_leaf_4_PCLK),
    .D(n645),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net243));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_10_ (.CLK(clknet_leaf_0_PCLK),
    .D(n655),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net368));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_11_ (.CLK(clknet_leaf_17_PCLK),
    .D(n656),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net369));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_12_ (.CLK(clknet_leaf_17_PCLK),
    .D(n657),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net370));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_13_ (.CLK(clknet_leaf_17_PCLK),
    .D(n658),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net371));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_14_ (.CLK(clknet_leaf_17_PCLK),
    .D(n659),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net372));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_15_ (.CLK(clknet_leaf_16_PCLK),
    .D(n660),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net373));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_16_ (.CLK(clknet_leaf_17_PCLK),
    .D(n661),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net374));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_17_ (.CLK(clknet_leaf_17_PCLK),
    .D(n662),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net375));
 sky130_fd_sc_hd__dfrtp_1 reg_left_opamp_ctrl_REG_reg_1_ (.CLK(clknet_leaf_5_PCLK),
    .D(n646),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net325));
 sky130_fd_sc_hd__dfrtp_2 reg_left_opamp_ctrl_REG_reg_2_ (.CLK(clknet_leaf_0_PCLK),
    .D(n647),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net360));
 sky130_fd_sc_hd__dfrtp_2 reg_left_opamp_ctrl_REG_reg_3_ (.CLK(clknet_leaf_4_PCLK),
    .D(n648),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net361));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_4_ (.CLK(clknet_leaf_5_PCLK),
    .D(n649),
    .RESET_B(net678),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net362));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_5_ (.CLK(clknet_leaf_0_PCLK),
    .D(n650),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net363));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_6_ (.CLK(clknet_leaf_17_PCLK),
    .D(n651),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net364));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_7_ (.CLK(clknet_leaf_5_PCLK),
    .D(n652),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net365));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_8_ (.CLK(clknet_leaf_4_PCLK),
    .D(n653),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net366));
 sky130_fd_sc_hd__dfrtp_4 reg_left_opamp_ctrl_REG_reg_9_ (.CLK(clknet_leaf_0_PCLK),
    .D(n654),
    .RESET_B(net677),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net367));
 sky130_fd_sc_hd__dfrtp_1 reg_rdac_ctrl_REG_reg_0_ (.CLK(clknet_leaf_0_PCLK),
    .D(n511),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net382));
 sky130_fd_sc_hd__dfrtp_1 reg_rdac_ctrl_REG_reg_10_ (.CLK(clknet_leaf_0_PCLK),
    .D(n521),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net394));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_11_ (.CLK(clknet_leaf_17_PCLK),
    .D(n522),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net384));
 sky130_fd_sc_hd__dfrtp_2 reg_rdac_ctrl_REG_reg_12_ (.CLK(clknet_leaf_17_PCLK),
    .D(n523),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net385));
 sky130_fd_sc_hd__dfrtp_2 reg_rdac_ctrl_REG_reg_13_ (.CLK(clknet_leaf_18_PCLK),
    .D(n524),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net395));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_14_ (.CLK(clknet_leaf_17_PCLK),
    .D(n525),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net396));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_15_ (.CLK(clknet_leaf_0_PCLK),
    .D(n526),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net399));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_16_ (.CLK(clknet_leaf_17_PCLK),
    .D(n527),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net400));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_17_ (.CLK(clknet_leaf_0_PCLK),
    .D(n528),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net401));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_18_ (.CLK(clknet_leaf_18_PCLK),
    .D(n529),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net402));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_19_ (.CLK(clknet_leaf_17_PCLK),
    .D(n530),
    .RESET_B(net676),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net403));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_1_ (.CLK(clknet_leaf_4_PCLK),
    .D(n512),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net383));
 sky130_fd_sc_hd__dfrtp_2 reg_rdac_ctrl_REG_reg_20_ (.CLK(clknet_leaf_18_PCLK),
    .D(n531),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net404));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_21_ (.CLK(clknet_leaf_18_PCLK),
    .D(n532),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net405));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_22_ (.CLK(clknet_leaf_18_PCLK),
    .D(n533),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net406));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_23_ (.CLK(clknet_leaf_18_PCLK),
    .D(n534),
    .RESET_B(net671),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net407));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_24_ (.CLK(clknet_leaf_18_PCLK),
    .D(n535),
    .RESET_B(net673),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net397));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_25_ (.CLK(clknet_leaf_18_PCLK),
    .D(n536),
    .RESET_B(net668),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net398));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_2_ (.CLK(clknet_leaf_18_PCLK),
    .D(n513),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net386));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_3_ (.CLK(clknet_leaf_18_PCLK),
    .D(n514),
    .RESET_B(net669),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net387));
 sky130_fd_sc_hd__dfrtp_1 reg_rdac_ctrl_REG_reg_4_ (.CLK(clknet_leaf_0_PCLK),
    .D(n515),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net388));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_5_ (.CLK(clknet_leaf_0_PCLK),
    .D(n516),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net389));
 sky130_fd_sc_hd__dfrtp_1 reg_rdac_ctrl_REG_reg_6_ (.CLK(clknet_leaf_0_PCLK),
    .D(n517),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net390));
 sky130_fd_sc_hd__dfrtp_2 reg_rdac_ctrl_REG_reg_7_ (.CLK(clknet_leaf_18_PCLK),
    .D(n518),
    .RESET_B(net674),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net391));
 sky130_fd_sc_hd__dfrtp_4 reg_rdac_ctrl_REG_reg_8_ (.CLK(clknet_leaf_4_PCLK),
    .D(n519),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net392));
 sky130_fd_sc_hd__dfrtp_1 reg_rdac_ctrl_REG_reg_9_ (.CLK(clknet_leaf_4_PCLK),
    .D(n520),
    .RESET_B(net675),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net393));
 sky130_fd_sc_hd__dfrtp_4 reg_right_instramp_ctrl_REG_reg_0_ (.CLK(clknet_leaf_11_PCLK),
    .D(n634),
    .RESET_B(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net461));
 sky130_fd_sc_hd__dfrtp_2 reg_right_instramp_ctrl_REG_reg_10_ (.CLK(clknet_leaf_15_PCLK),
    .D(n644),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net460));
 sky130_fd_sc_hd__dfrtp_2 reg_right_instramp_ctrl_REG_reg_1_ (.CLK(clknet_leaf_16_PCLK),
    .D(n635),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net451));
 sky130_fd_sc_hd__dfrtp_4 reg_right_instramp_ctrl_REG_reg_2_ (.CLK(clknet_leaf_15_PCLK),
    .D(n636),
    .RESET_B(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net452));
 sky130_fd_sc_hd__dfrtp_4 reg_right_instramp_ctrl_REG_reg_3_ (.CLK(clknet_leaf_15_PCLK),
    .D(n637),
    .RESET_B(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net453));
 sky130_fd_sc_hd__dfrtp_4 reg_right_instramp_ctrl_REG_reg_4_ (.CLK(clknet_leaf_11_PCLK),
    .D(n638),
    .RESET_B(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net454));
 sky130_fd_sc_hd__dfrtp_2 reg_right_instramp_ctrl_REG_reg_5_ (.CLK(clknet_leaf_15_PCLK),
    .D(n639),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net455));
 sky130_fd_sc_hd__dfrtp_2 reg_right_instramp_ctrl_REG_reg_6_ (.CLK(clknet_leaf_16_PCLK),
    .D(n640),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net456));
 sky130_fd_sc_hd__dfrtp_2 reg_right_instramp_ctrl_REG_reg_7_ (.CLK(clknet_leaf_15_PCLK),
    .D(n641),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net457));
 sky130_fd_sc_hd__dfrtp_1 reg_right_instramp_ctrl_REG_reg_8_ (.CLK(clknet_leaf_16_PCLK),
    .D(n642),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net458));
 sky130_fd_sc_hd__dfrtp_1 reg_right_instramp_ctrl_REG_reg_9_ (.CLK(clknet_leaf_15_PCLK),
    .D(n643),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net459));
 sky130_fd_sc_hd__dfrtp_4 reg_right_opamp_ctrl_REG_reg_0_ (.CLK(clknet_leaf_16_PCLK),
    .D(n616),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net408));
 sky130_fd_sc_hd__dfrtp_2 reg_right_opamp_ctrl_REG_reg_10_ (.CLK(clknet_leaf_11_PCLK),
    .D(n626),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net537));
 sky130_fd_sc_hd__dfrtp_2 reg_right_opamp_ctrl_REG_reg_11_ (.CLK(clknet_leaf_15_PCLK),
    .D(n627),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net538));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_12_ (.CLK(clknet_leaf_16_PCLK),
    .D(n628),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net539));
 sky130_fd_sc_hd__dfrtp_4 reg_right_opamp_ctrl_REG_reg_13_ (.CLK(clknet_leaf_14_PCLK),
    .D(n629),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net540));
 sky130_fd_sc_hd__dfrtp_4 reg_right_opamp_ctrl_REG_reg_14_ (.CLK(clknet_leaf_15_PCLK),
    .D(n630),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net541));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_15_ (.CLK(clknet_leaf_15_PCLK),
    .D(n631),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net542));
 sky130_fd_sc_hd__dfrtp_2 reg_right_opamp_ctrl_REG_reg_16_ (.CLK(clknet_leaf_15_PCLK),
    .D(n632),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net543));
 sky130_fd_sc_hd__dfrtp_4 reg_right_opamp_ctrl_REG_reg_17_ (.CLK(clknet_leaf_16_PCLK),
    .D(n633),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net544));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_1_ (.CLK(clknet_leaf_6_PCLK),
    .D(n617),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net489));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_2_ (.CLK(clknet_leaf_6_PCLK),
    .D(n618),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net529));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_3_ (.CLK(clknet_leaf_6_PCLK),
    .D(n619),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net530));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_4_ (.CLK(clknet_leaf_10_PCLK),
    .D(n620),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net531));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_5_ (.CLK(clknet_leaf_7_PCLK),
    .D(n621),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net532));
 sky130_fd_sc_hd__dfrtp_2 reg_right_opamp_ctrl_REG_reg_6_ (.CLK(clknet_leaf_6_PCLK),
    .D(n622),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net533));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_7_ (.CLK(clknet_leaf_6_PCLK),
    .D(n623),
    .RESET_B(net687),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net534));
 sky130_fd_sc_hd__dfrtp_1 reg_right_opamp_ctrl_REG_reg_8_ (.CLK(clknet_leaf_10_PCLK),
    .D(n624),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net535));
 sky130_fd_sc_hd__dfrtp_2 reg_right_opamp_ctrl_REG_reg_9_ (.CLK(clknet_leaf_11_PCLK),
    .D(n625),
    .RESET_B(net688),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net536));
 sky130_fd_sc_hd__dfrtp_4 reg_tempsense_ctrl_REG_reg_0_ (.CLK(clknet_leaf_16_PCLK),
    .D(n537),
    .RESET_B(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net550));
 sky130_fd_sc_hd__dfrtp_1 reg_tempsense_ctrl_REG_reg_1_ (.CLK(clknet_leaf_17_PCLK),
    .D(n538),
    .RESET_B(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Q(net551));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_34 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_35 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_36 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_37 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_38 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_39 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_40 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_41 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_42 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_43 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_44 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_45 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_46 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_47 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_48 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_49 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_50 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_52 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_53 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_54 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_56 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_57 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_58 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_59 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_60 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_61 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_62 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_63 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_64 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_65 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_66 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_67 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_68 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_69 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_70 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_71 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_72 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_73 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_74 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_75 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_76 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_77 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_89 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_90 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_91 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_92 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_93 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_94 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_95 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_96 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_97 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_98 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_99 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_100 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_101 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_102 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_103 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_104 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_105 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_106 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_107 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_108 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_109 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_110 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_111 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_112 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_113 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_114 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_115 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_116 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_117 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_118 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_119 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_120 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_121 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_122 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_123 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_124 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_125 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_126 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_127 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_128 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_129 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_130 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_131 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_132 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_133 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_134 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_135 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_136 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_137 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_138 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_139 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_140 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_141 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_142 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_143 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_144 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_145 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_146 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_147 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_148 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_149 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_150 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_151 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_152 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_153 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_154 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_155 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_156 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_157 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_158 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_159 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_160 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_161 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_178 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_179 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_180 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_181 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_182 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_183 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_184 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_185 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_186 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_187 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_188 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_189 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_190 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_191 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_192 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_193 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_194 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_195 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_196 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_197 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_198 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_199 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_200 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_201 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_202 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_203 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_204 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_205 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_206 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_207 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_208 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_209 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_210 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_211 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_212 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_213 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_214 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_215 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_216 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_217 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_218 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_219 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_220 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_221 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_222 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_223 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_224 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_225 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_226 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_227 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_228 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_229 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_230 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_231 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_232 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_233 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_234 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_235 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_236 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_237 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_238 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_239 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_240 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_241 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_242 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_243 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_244 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_245 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_246 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_247 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_248 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_249 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_250 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_251 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_252 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_253 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_254 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_255 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_256 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_257 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_258 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_259 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_260 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_261 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_262 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_263 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_264 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_265 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_266 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_267 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_268 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_269 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_270 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_271 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_272 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_273 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_274 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_275 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_276 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_277 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_278 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_279 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_280 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_281 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_282 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_283 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_284 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_285 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_286 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_287 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_288 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_289 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_290 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_291 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_292 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_293 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_294 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_295 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_296 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_297 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_298 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_299 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_300 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_301 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_302 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_303 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_304 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_305 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_306 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_307 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_308 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_309 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_310 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_311 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_312 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_313 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_314 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_315 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_316 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_317 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_318 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_319 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_320 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_321 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_322 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_323 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_324 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_325 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_326 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_327 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_328 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_329 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_330 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_331 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_332 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_333 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_334 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_335 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_336 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_337 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_338 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_339 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_340 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_341 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_342 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_343 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_344 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_345 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_346 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_347 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_348 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_349 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_350 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_351 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_352 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_353 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_354 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_355 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_356 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_357 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_358 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_359 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_360 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_361 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_362 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_363 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_364 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_365 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_366 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_367 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_368 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_369 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_370 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_371 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_372 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_373 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_374 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_375 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_376 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_377 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_378 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_379 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_380 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_381 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_382 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_383 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_384 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_385 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_386 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_387 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_388 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_389 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_390 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_391 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_392 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_393 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_394 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_395 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_396 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_397 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_398 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_399 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_400 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_401 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_402 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_403 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_404 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_405 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_406 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_407 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_408 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_409 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_410 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_411 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_412 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_413 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_414 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_415 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_416 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_417 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_418 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_419 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_420 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_421 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_422 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_423 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_424 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_425 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_426 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_427 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_428 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_429 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_430 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_431 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_432 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_433 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_434 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_435 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_436 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_437 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_438 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_439 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_440 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_441 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_442 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_443 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_444 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_445 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_446 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_447 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_448 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_449 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_450 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_451 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_452 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_453 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_454 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_455 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_456 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_457 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_458 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_459 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_460 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_461 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_462 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_463 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_464 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_465 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_466 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_467 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_468 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_469 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_470 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_471 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_472 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_473 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_474 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_475 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_476 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_477 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_478 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_479 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_480 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_481 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_482 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_483 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_484 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_485 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_486 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_487 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_488 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_489 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_490 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_491 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_492 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_493 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_494 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_495 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_496 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_497 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_498 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_499 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_500 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_501 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_502 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_503 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_504 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_505 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_506 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_507 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_508 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_509 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_510 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_511 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_512 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_513 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_514 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_515 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_516 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_517 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_518 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_519 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_520 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_521 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_522 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_523 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_524 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_525 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_526 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_527 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_528 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_529 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_530 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_531 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_532 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_533 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_534 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_535 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_536 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_537 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_538 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_539 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_540 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_541 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_542 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_543 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_544 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_545 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_546 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_547 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_548 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_549 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_550 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_551 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_552 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_553 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_554 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_555 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_556 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_557 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_558 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_559 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_560 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_561 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_562 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_563 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_564 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_565 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_566 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_567 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_568 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_569 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_570 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_571 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_572 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_573 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_574 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_575 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_576 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_577 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_578 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_579 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_580 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_581 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_582 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_583 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_584 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_585 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_586 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_587 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_588 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_589 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_590 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_591 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_592 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_593 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_594 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_595 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_596 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_597 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_598 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_599 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_600 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_601 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_602 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_603 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_604 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_605 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_606 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_607 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_608 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_609 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_610 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_611 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_612 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_613 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_614 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_615 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_616 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_617 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_618 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_619 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_620 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_621 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_622 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_623 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_624 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_625 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_626 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_627 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_628 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_629 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_630 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_631 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_632 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_633 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_634 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_635 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_636 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_637 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_638 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_639 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_640 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_641 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_642 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_643 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_644 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_645 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_646 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_647 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_648 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_649 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_650 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_651 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_652 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_653 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_654 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_655 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_656 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_657 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_658 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_659 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_660 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_661 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_662 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_663 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_664 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_665 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_666 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_667 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_668 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_669 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_670 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_671 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_672 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_673 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_674 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_675 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_676 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_677 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_678 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_679 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_680 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_681 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_682 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_683 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_684 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_685 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_686 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_687 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_688 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_689 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_690 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_691 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_692 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_693 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_694 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_695 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_696 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_697 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_698 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_699 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_700 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_701 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_702 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_703 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_704 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_705 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_706 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_707 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_708 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_709 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_710 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_711 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_712 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_713 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_714 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_715 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_716 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_717 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_718 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_719 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_720 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_721 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_722 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_723 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_724 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_725 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_726 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_727 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_728 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_729 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_730 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_731 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_732 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_733 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_734 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_735 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_736 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_737 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_738 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_739 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_740 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_741 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_742 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_743 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_744 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_745 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_746 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_747 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_748 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_749 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_750 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_751 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_752 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_753 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_754 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_755 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_756 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_757 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_758 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_759 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_760 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_761 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_762 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_763 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_764 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_765 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_766 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_767 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_768 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_769 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_770 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_771 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_772 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_773 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_774 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_775 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_776 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_777 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_778 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_779 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_780 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_781 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_782 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_783 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_784 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_785 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_786 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_787 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_788 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_789 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_790 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_791 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_792 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_793 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_794 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_795 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_796 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_797 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_798 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_799 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_800 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_801 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_802 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_803 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_804 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_805 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_806 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_807 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_808 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_809 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_810 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_811 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_812 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_813 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_814 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_815 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_816 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_817 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_818 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_819 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_820 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_821 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_822 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_823 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_824 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_825 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_826 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_827 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_828 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_829 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_830 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_831 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_832 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_833 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_834 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_835 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_836 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_837 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_838 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_839 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_840 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_841 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_842 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_843 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_844 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_845 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_846 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_847 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_848 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_849 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_850 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_851 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_852 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_853 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_854 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_855 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_856 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_857 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_858 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_859 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_860 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_861 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_862 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_863 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_864 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_865 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_866 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_867 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_868 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_869 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_870 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_871 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_872 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_873 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_874 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_875 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_876 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_877 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_878 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_879 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_880 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_881 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_882 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_883 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_884 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_885 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_886 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_887 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_888 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_889 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_890 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_891 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_892 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_893 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_894 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_895 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_896 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_897 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_898 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_899 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_900 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_901 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_902 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_903 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_904 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_905 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_906 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_907 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_908 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_909 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_910 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_911 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_912 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_913 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_914 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_915 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_916 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_917 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_918 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_919 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_920 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_921 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_922 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_923 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_924 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_925 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_926 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_927 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_928 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_929 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_930 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_931 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_932 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_933 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_934 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_935 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_936 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_937 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_938 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_939 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_940 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_941 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_942 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_943 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_944 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_945 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_946 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_947 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_948 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_949 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_950 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_951 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_952 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_953 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_954 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_955 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_956 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_957 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_958 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_959 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_960 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_961 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_962 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_963 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_964 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_965 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_966 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_967 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_968 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_969 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_970 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_971 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_972 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_973 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_974 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_975 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_976 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_977 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_978 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_979 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_980 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_981 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_982 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_983 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_984 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_985 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_986 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_987 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_988 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_989 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_990 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_991 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_992 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_993 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_994 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_995 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_996 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_997 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_998 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_999 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1000 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1001 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1002 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1003 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1004 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1005 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1006 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1007 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1008 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1009 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1010 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1011 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1012 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1013 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1014 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1015 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1016 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1017 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1018 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1019 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1020 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1021 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1022 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1023 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1024 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1025 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1026 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1027 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1028 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1029 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1030 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1031 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1032 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1033 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1034 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1035 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1036 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1037 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1038 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1039 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1040 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1041 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1042 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1043 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1044 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1045 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1046 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1047 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1048 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1049 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1050 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_1051 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1052 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1053 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1054 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1055 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1056 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1057 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1058 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1059 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1060 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1061 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1062 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1063 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1064 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1065 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1066 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1067 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1068 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1069 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1070 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1071 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1072 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1073 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1074 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1075 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1076 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1077 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1078 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1079 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1080 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1081 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1082 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1083 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1084 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1085 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1086 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1087 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1088 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1089 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1090 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1091 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1092 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1093 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1094 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1095 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1096 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1097 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1098 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1099 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1100 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1101 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1102 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1103 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1104 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1105 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1106 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1107 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1108 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1109 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1110 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1111 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_1112 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1113 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1114 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1115 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1116 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1117 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1118 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1119 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1120 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1121 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1122 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1123 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1124 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1125 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1126 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1127 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1128 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1129 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1130 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1131 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1132 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1133 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1134 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1135 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1136 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1137 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1138 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1139 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1140 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1141 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1142 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1143 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1144 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1145 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1146 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1147 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1148 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1149 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1150 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1151 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1152 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1153 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1154 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1155 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1156 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1157 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1158 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1159 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1160 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1161 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1162 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1163 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1164 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1165 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1166 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1167 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1168 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1169 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1170 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1171 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1172 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1173 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_1174 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1175 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1176 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1177 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1178 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1179 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1180 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1181 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1182 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1183 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1184 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1185 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1186 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1187 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1188 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1189 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1190 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1191 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1192 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1193 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1194 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1195 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1196 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1197 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1198 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1199 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1200 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1201 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1202 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1203 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1204 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1205 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1206 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1207 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1208 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1209 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1210 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1211 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1212 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1213 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1214 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1215 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1216 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1217 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1218 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1219 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1220 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1221 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1222 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1223 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1224 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1225 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1226 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1227 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1228 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1229 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1230 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1231 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1232 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1233 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1234 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_1235 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1236 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1237 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1238 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1239 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1240 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1241 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1242 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1243 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1244 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1245 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1246 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1247 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1248 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1249 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1250 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1251 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1252 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1253 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1254 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1255 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1256 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1257 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1258 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1259 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1260 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1261 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1262 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1263 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1264 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1265 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1266 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1267 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1268 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1269 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1270 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1271 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1272 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1273 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1274 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1275 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1276 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1277 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1278 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1279 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1280 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1281 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1282 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1283 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1284 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1285 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1286 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1287 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1288 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1289 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1290 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1291 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1292 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1293 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1294 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1295 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1296 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_1297 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1298 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1299 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1300 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1301 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1302 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1303 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1304 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1305 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1306 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1307 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1308 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1309 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1310 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1311 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1312 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1313 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1314 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1315 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1316 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1317 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1318 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1319 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1320 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1321 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1322 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1323 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1324 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1325 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1326 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1327 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1328 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1329 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1330 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1331 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1332 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1333 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1334 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1335 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1336 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1337 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1338 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1339 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1340 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1341 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1342 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1343 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1344 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1345 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1346 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1347 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1348 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1349 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1350 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1351 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1352 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1353 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1354 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1355 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1356 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1357 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_1358 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1359 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1360 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1361 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1362 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1363 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1364 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1365 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1366 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1367 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1368 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1369 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1370 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1371 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1372 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1373 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1374 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1375 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1376 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1377 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1378 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1379 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1380 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1381 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1382 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1383 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1384 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1385 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1386 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1387 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1388 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1389 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1390 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1391 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1392 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1393 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1394 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1395 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1396 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1397 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1398 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1399 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1400 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1401 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1402 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1403 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1404 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1405 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1406 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1407 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1408 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1409 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1410 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1411 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1412 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1413 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1414 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1415 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1416 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1417 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1418 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1419 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_1420 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1421 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1422 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1423 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1424 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1425 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1426 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1427 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1428 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1429 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1430 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1431 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1432 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1433 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1434 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1435 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1436 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1437 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1438 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1439 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1440 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1441 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1442 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1443 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1444 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1445 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1446 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1447 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1448 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1449 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1450 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1451 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1452 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1453 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1454 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1455 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1456 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1457 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1458 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1459 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1460 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1461 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1462 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1463 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1464 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1465 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1466 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1467 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1468 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1469 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1470 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1471 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1472 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1473 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1474 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1475 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1476 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1477 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1478 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1479 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1480 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_1481 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1482 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1483 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1484 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1485 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1486 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1487 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1488 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1489 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1490 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1491 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1492 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1493 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1494 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1495 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1496 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1497 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1498 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1499 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1500 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1501 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1502 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1503 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1504 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1505 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1506 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1507 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1508 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1509 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1510 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1511 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1512 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1513 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1514 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1515 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1516 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1517 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1518 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1519 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1520 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1521 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1522 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1523 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1524 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1525 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1526 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1527 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1528 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1529 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1530 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1531 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1532 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1533 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1534 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1535 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1536 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1537 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1538 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1539 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1540 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1541 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1542 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_1543 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1544 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1545 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1546 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1547 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1548 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1549 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1550 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1551 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1552 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1553 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1554 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1555 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1556 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1557 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1558 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1559 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1560 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1561 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1562 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1563 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1564 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1565 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1566 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1567 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1568 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1569 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1570 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1571 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1572 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1573 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1574 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1575 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1576 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1577 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1578 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1579 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1580 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1581 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1582 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1583 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1584 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1585 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1586 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1587 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1588 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1589 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1590 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1591 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1592 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1593 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1594 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1595 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1596 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1597 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1598 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1599 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1600 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1601 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1602 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1603 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_1604 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1605 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1606 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1607 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1608 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1609 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1610 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1611 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1612 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1613 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1614 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1615 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1616 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1617 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1618 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1619 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1620 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1621 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1622 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1623 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1624 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1625 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1626 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1627 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1628 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1629 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1630 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1631 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1632 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1633 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1634 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1635 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1636 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1637 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1638 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1639 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1640 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1641 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1642 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1643 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1644 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1645 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1646 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1647 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1648 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1649 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1650 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1651 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1652 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1653 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1654 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1655 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1656 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1657 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1658 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1659 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1660 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1661 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1662 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1663 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1664 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1665 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_1666 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1667 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1668 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1669 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1670 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1671 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1672 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1673 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1674 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1675 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1676 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1677 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1678 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1679 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1680 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1681 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1682 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1683 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1684 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1685 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1686 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1687 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1688 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1689 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1690 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1691 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1692 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1693 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1694 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1695 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1696 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1697 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1698 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1699 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1700 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1701 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1702 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1703 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1704 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1705 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1706 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1707 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1708 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1709 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1710 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1711 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1712 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1713 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1714 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1715 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1716 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1717 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1718 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1719 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1720 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1721 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1722 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1723 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1724 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1725 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1726 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_1727 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1728 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1729 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1730 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1731 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1732 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1733 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1734 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1735 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1736 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1737 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1738 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1739 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1740 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1741 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1742 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1743 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1744 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1745 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1746 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1747 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1748 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1749 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1750 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1751 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1752 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1753 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1754 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1755 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1756 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1757 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1758 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1759 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1760 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1761 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1762 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1763 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1764 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1765 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1766 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1767 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1768 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1769 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1770 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1771 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1772 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1773 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1774 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1775 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1776 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1777 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1778 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1779 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1780 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1781 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1782 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1783 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1784 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1785 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1786 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1787 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1788 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_1789 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1790 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1791 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1792 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1793 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1794 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1795 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1796 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1797 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1798 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1799 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1800 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1801 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1802 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1803 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1804 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1805 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1806 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1807 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1808 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1809 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1810 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1811 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1812 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1813 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1814 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1815 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1816 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1817 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1818 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1819 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1820 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1821 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1822 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1823 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1824 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1825 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1826 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1827 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1828 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1829 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1830 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1831 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1832 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1833 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1834 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1835 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1836 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1837 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1838 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1839 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1840 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1841 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1842 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1843 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1844 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1845 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1846 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1847 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1848 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1849 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_1850 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1851 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1852 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1853 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1854 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1855 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1856 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1857 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1858 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1859 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1860 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1861 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1862 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1863 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1864 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1865 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1866 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1867 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1868 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1869 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1870 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1871 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1872 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1873 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1874 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1875 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1876 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1877 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1878 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1879 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1880 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1881 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1882 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1883 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1884 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1885 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1886 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1887 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1888 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1889 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1890 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1891 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1892 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1893 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1894 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1895 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1896 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1897 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1898 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1899 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1900 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1901 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1902 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1903 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1904 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1905 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1906 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1907 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1908 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1909 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1910 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1911 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_1912 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1913 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1914 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1915 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1916 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1917 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1918 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1919 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1920 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1921 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1922 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1923 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1924 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1925 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1926 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1927 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1928 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1929 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1930 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1931 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1932 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1933 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1934 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1935 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1936 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1937 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1938 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1939 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1940 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1941 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1942 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1943 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1944 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1945 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1946 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1947 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1948 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1949 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1950 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1951 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1952 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1953 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1954 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1955 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1956 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1957 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1958 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1959 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1960 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1961 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1962 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1963 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1964 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1965 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1966 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1967 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1968 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1969 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1970 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1971 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1972 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_1973 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1974 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1975 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1976 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1977 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1978 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1979 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1980 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1981 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1982 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1983 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1984 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1985 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1986 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1987 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1988 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1989 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1990 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1991 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1992 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1993 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1994 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1995 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1996 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1997 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1998 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_1999 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2000 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2001 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2002 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2003 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2004 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2005 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2006 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2007 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2008 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2009 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2010 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2011 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2012 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2013 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2014 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2015 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2016 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2017 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2018 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2019 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2020 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2021 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2022 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2023 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2024 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2025 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2026 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2027 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2028 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2029 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2030 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2031 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2032 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2033 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2034 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_2035 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2036 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2037 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2038 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2039 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2040 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2041 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2042 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2043 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2044 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2045 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2046 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2047 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2048 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2049 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2050 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2051 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2052 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2053 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2054 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2055 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2056 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2057 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2058 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2059 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2060 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2061 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2062 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2063 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2064 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2065 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2066 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2067 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2068 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2069 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2070 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2071 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2072 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2073 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2074 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2075 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2076 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2077 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2078 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2079 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2080 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2081 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2082 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2083 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2084 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2085 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2086 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2087 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2088 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2089 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2090 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2091 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2092 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2093 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2094 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2095 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_2096 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2097 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2098 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2099 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2100 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2101 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2102 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2103 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2104 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2105 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2106 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2107 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2108 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2109 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2110 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2111 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2112 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2113 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2114 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2115 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2116 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2117 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2118 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2119 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2120 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2121 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2122 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2123 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2124 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2125 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2126 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2127 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2128 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2129 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2130 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2131 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2132 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2133 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2134 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2135 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2136 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2137 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2138 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2139 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2140 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2141 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2142 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2143 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2144 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2145 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2146 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2147 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2148 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2149 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2150 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2151 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2152 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2153 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2154 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2155 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2156 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2157 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_2158 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2159 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2160 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2161 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2162 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2163 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2164 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2165 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2166 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2167 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2168 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2169 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2170 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2171 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2172 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2173 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2174 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2175 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2176 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2177 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2178 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2179 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2180 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2181 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2182 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2183 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2184 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2185 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2186 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2187 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2188 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2189 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2190 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2191 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2192 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2193 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2194 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2195 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2196 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2197 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2198 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2199 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2200 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2201 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2202 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2203 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2204 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2205 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2206 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2207 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2208 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2209 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2210 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2211 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2212 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2213 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2214 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2215 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2216 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2217 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2218 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2219 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2220 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2221 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2222 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2223 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2224 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2225 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2226 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2227 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2228 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2229 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2230 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2231 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2232 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2233 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2234 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2235 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2236 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2237 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2238 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2239 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2240 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2241 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2242 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2243 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2244 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2245 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2246 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2247 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2248 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2249 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2250 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2251 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2252 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2253 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2254 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2255 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2256 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2257 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2258 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2259 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2260 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2261 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2262 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2263 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2264 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2265 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2266 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2267 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2268 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2269 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2270 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2271 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2272 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2273 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2274 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2275 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2276 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2277 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2278 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2279 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2280 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_2281 (.VGND(vssd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__buf_6 input1 (.A(PADDR[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(PADDR[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(PADDR[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(PADDR[12]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(PADDR[13]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(PADDR[14]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(PADDR[15]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net7));
 sky130_fd_sc_hd__buf_6 input8 (.A(PADDR[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net8));
 sky130_fd_sc_hd__buf_6 input9 (.A(PADDR[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net9));
 sky130_fd_sc_hd__buf_12 input10 (.A(PADDR[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_8 input11 (.A(PADDR[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net11));
 sky130_fd_sc_hd__buf_12 input12 (.A(PADDR[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net12));
 sky130_fd_sc_hd__buf_6 input13 (.A(PADDR[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(PADDR[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net14));
 sky130_fd_sc_hd__buf_6 input15 (.A(PADDR[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net15));
 sky130_fd_sc_hd__buf_6 input16 (.A(PADDR[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(PENABLE),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net17));
 sky130_fd_sc_hd__buf_6 input18 (.A(PRESETn),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(PSEL),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net19));
 sky130_fd_sc_hd__buf_6 input20 (.A(PWDATA[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net20));
 sky130_fd_sc_hd__buf_8 input21 (.A(PWDATA[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net21));
 sky130_fd_sc_hd__buf_6 input22 (.A(PWDATA[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_16 input23 (.A(PWDATA[12]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_16 input24 (.A(PWDATA[13]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net24));
 sky130_fd_sc_hd__buf_6 input25 (.A(PWDATA[14]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(PWDATA[15]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net26));
 sky130_fd_sc_hd__buf_6 input27 (.A(PWDATA[16]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(PWDATA[17]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(PWDATA[18]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net29));
 sky130_fd_sc_hd__buf_4 input30 (.A(PWDATA[19]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net30));
 sky130_fd_sc_hd__buf_6 input31 (.A(PWDATA[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_8 input32 (.A(PWDATA[20]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(PWDATA[21]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net33));
 sky130_fd_sc_hd__buf_2 input34 (.A(PWDATA[22]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_2 input35 (.A(PWDATA[23]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net35));
 sky130_fd_sc_hd__buf_2 input36 (.A(PWDATA[24]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net36));
 sky130_fd_sc_hd__dlymetal6s2s_1 input37 (.A(PWDATA[25]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net37));
 sky130_fd_sc_hd__buf_1 input38 (.A(PWDATA[26]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net38));
 sky130_fd_sc_hd__buf_1 input39 (.A(PWDATA[27]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net39));
 sky130_fd_sc_hd__buf_1 input40 (.A(PWDATA[28]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net40));
 sky130_fd_sc_hd__buf_1 input41 (.A(PWDATA[29]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(PWDATA[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(PWDATA[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net43));
 sky130_fd_sc_hd__buf_6 input44 (.A(PWDATA[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net44));
 sky130_fd_sc_hd__buf_6 input45 (.A(PWDATA[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net45));
 sky130_fd_sc_hd__buf_8 input46 (.A(PWDATA[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net46));
 sky130_fd_sc_hd__buf_6 input47 (.A(PWDATA[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(PWDATA[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_2 input49 (.A(PWDATA[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 input50 (.A(PWRITE),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net50));
 sky130_fd_sc_hd__buf_1 input51 (.A(brownout_filt),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(brownout_timeout),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(brownout_unfilt),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(brownout_vunder),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net54));
 sky130_fd_sc_hd__buf_1 input55 (.A(comp_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net55));
 sky130_fd_sc_hd__buf_1 input56 (.A(overvoltage_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net56));
 sky130_fd_sc_hd__buf_1 input57 (.A(ulpcomp_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_2 input58 (.A(vccd1_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(vccd2_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_2 input60 (.A(vdda1_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net60));
 sky130_fd_sc_hd__dlymetal6s2s_1 input61 (.A(vdda2_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net61));
 sky130_fd_sc_hd__buf_12 output62 (.A(net62),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[0]));
 sky130_fd_sc_hd__clkbuf_8 output63 (.A(net63),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[10]));
 sky130_fd_sc_hd__clkbuf_8 output64 (.A(net64),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[11]));
 sky130_fd_sc_hd__clkbuf_8 output65 (.A(net65),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[12]));
 sky130_fd_sc_hd__clkbuf_8 output66 (.A(net66),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[13]));
 sky130_fd_sc_hd__clkbuf_8 output67 (.A(net67),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[14]));
 sky130_fd_sc_hd__clkbuf_8 output68 (.A(net68),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[15]));
 sky130_fd_sc_hd__clkbuf_8 output69 (.A(net69),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[16]));
 sky130_fd_sc_hd__clkbuf_8 output70 (.A(net70),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[17]));
 sky130_fd_sc_hd__clkbuf_8 output71 (.A(net71),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[18]));
 sky130_fd_sc_hd__clkbuf_8 output72 (.A(net72),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[19]));
 sky130_fd_sc_hd__clkbuf_8 output73 (.A(net73),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[1]));
 sky130_fd_sc_hd__clkbuf_8 output74 (.A(net74),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[20]));
 sky130_fd_sc_hd__clkbuf_8 output75 (.A(net75),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[21]));
 sky130_fd_sc_hd__clkbuf_8 output76 (.A(net76),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[22]));
 sky130_fd_sc_hd__clkbuf_8 output77 (.A(net77),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[23]));
 sky130_fd_sc_hd__clkbuf_8 output78 (.A(net78),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[24]));
 sky130_fd_sc_hd__clkbuf_8 output79 (.A(net79),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[25]));
 sky130_fd_sc_hd__clkbuf_8 output80 (.A(net80),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[26]));
 sky130_fd_sc_hd__clkbuf_8 output81 (.A(net81),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[27]));
 sky130_fd_sc_hd__clkbuf_8 output82 (.A(net82),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[28]));
 sky130_fd_sc_hd__clkbuf_8 output83 (.A(net83),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[29]));
 sky130_fd_sc_hd__buf_12 output84 (.A(net84),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[2]));
 sky130_fd_sc_hd__clkbuf_8 output85 (.A(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[30]));
 sky130_fd_sc_hd__clkbuf_8 output86 (.A(net86),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[31]));
 sky130_fd_sc_hd__buf_8 output87 (.A(net87),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[3]));
 sky130_fd_sc_hd__clkbuf_8 output88 (.A(net88),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[4]));
 sky130_fd_sc_hd__buf_12 output89 (.A(net89),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[5]));
 sky130_fd_sc_hd__buf_12 output90 (.A(net90),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[6]));
 sky130_fd_sc_hd__buf_12 output91 (.A(net91),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[7]));
 sky130_fd_sc_hd__clkbuf_8 output92 (.A(net92),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[8]));
 sky130_fd_sc_hd__clkbuf_8 output93 (.A(net93),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(PRDATA[9]));
 sky130_fd_sc_hd__clkbuf_8 output94 (.A(net94),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output95 (.A(net95),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_dac0));
 sky130_fd_sc_hd__clkbuf_8 output96 (.A(net96),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_gpio1_3[0]));
 sky130_fd_sc_hd__clkbuf_8 output97 (.A(net97),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_gpio1_3[1]));
 sky130_fd_sc_hd__clkbuf_8 output98 (.A(net98),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_gpio6_4[0]));
 sky130_fd_sc_hd__clkbuf_8 output99 (.A(net99),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_gpio6_4[1]));
 sky130_fd_sc_hd__clkbuf_8 output100 (.A(net100),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output101 (.A(net101),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_tempsense));
 sky130_fd_sc_hd__clkbuf_8 output102 (.A(net102),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_vbgtc));
 sky130_fd_sc_hd__clkbuf_8 output103 (.A(net103),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc0_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output104 (.A(net104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output105 (.A(net105),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_dac1));
 sky130_fd_sc_hd__clkbuf_8 output106 (.A(net106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_gpio1_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output107 (.A(net107),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_gpio1_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output108 (.A(net108),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_gpio6_5[0]));
 sky130_fd_sc_hd__clkbuf_8 output109 (.A(net109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_gpio6_5[1]));
 sky130_fd_sc_hd__clkbuf_8 output110 (.A(net110),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output111 (.A(net111),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_vbgsc));
 sky130_fd_sc_hd__clkbuf_8 output112 (.A(net112),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc1_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output113 (.A(net113),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc_refh_to_gpio6_6[0]));
 sky130_fd_sc_hd__clkbuf_8 output114 (.A(net114),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc_refh_to_gpio6_6[1]));
 sky130_fd_sc_hd__clkbuf_8 output115 (.A(net115),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc_refl_to_gpio6_7[0]));
 sky130_fd_sc_hd__clkbuf_8 output116 (.A(net116),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(adc_refl_to_gpio6_7[1]));
 sky130_fd_sc_hd__clkbuf_8 output117 (.A(net117),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(analog0_connect[0]));
 sky130_fd_sc_hd__clkbuf_8 output118 (.A(net118),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(analog0_connect[1]));
 sky130_fd_sc_hd__clkbuf_8 output119 (.A(net119),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(analog1_connect[0]));
 sky130_fd_sc_hd__clkbuf_8 output120 (.A(net120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(analog1_connect[1]));
 sky130_fd_sc_hd__clkbuf_8 output121 (.A(net121),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(audiodac_out_to_analog1[0]));
 sky130_fd_sc_hd__clkbuf_8 output122 (.A(net122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(audiodac_out_to_analog1[1]));
 sky130_fd_sc_hd__clkbuf_8 output123 (.A(net123),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(audiodac_outb_to_analog0[0]));
 sky130_fd_sc_hd__clkbuf_8 output124 (.A(net124),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(audiodac_outb_to_analog0[1]));
 sky130_fd_sc_hd__clkbuf_8 output125 (.A(net125),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_ena));
 sky130_fd_sc_hd__clkbuf_8 output126 (.A(net126),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_sel));
 sky130_fd_sc_hd__clkbuf_8 output127 (.A(net127),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[0]));
 sky130_fd_sc_hd__clkbuf_8 output128 (.A(net128),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[10]));
 sky130_fd_sc_hd__clkbuf_8 output129 (.A(net129),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[11]));
 sky130_fd_sc_hd__clkbuf_8 output130 (.A(net130),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[12]));
 sky130_fd_sc_hd__clkbuf_8 output131 (.A(net131),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[13]));
 sky130_fd_sc_hd__clkbuf_8 output132 (.A(net132),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[14]));
 sky130_fd_sc_hd__clkbuf_8 output133 (.A(net133),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[15]));
 sky130_fd_sc_hd__clkbuf_8 output134 (.A(net134),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[1]));
 sky130_fd_sc_hd__clkbuf_8 output135 (.A(net135),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[2]));
 sky130_fd_sc_hd__clkbuf_8 output136 (.A(net136),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[3]));
 sky130_fd_sc_hd__clkbuf_8 output137 (.A(net137),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[4]));
 sky130_fd_sc_hd__clkbuf_8 output138 (.A(net138),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[5]));
 sky130_fd_sc_hd__clkbuf_8 output139 (.A(net139),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[6]));
 sky130_fd_sc_hd__clkbuf_8 output140 (.A(net140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[7]));
 sky130_fd_sc_hd__clkbuf_8 output141 (.A(net141),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[8]));
 sky130_fd_sc_hd__clkbuf_8 output142 (.A(net142),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(bandgap_trim[9]));
 sky130_fd_sc_hd__clkbuf_8 output143 (.A(net143),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_ena));
 sky130_fd_sc_hd__clkbuf_8 output144 (.A(net144),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_isrc_sel));
 sky130_fd_sc_hd__clkbuf_8 output145 (.A(net145),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_oneshot));
 sky130_fd_sc_hd__clkbuf_8 output146 (.A(net146),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_otrip[0]));
 sky130_fd_sc_hd__clkbuf_8 output147 (.A(net147),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_otrip[1]));
 sky130_fd_sc_hd__clkbuf_8 output148 (.A(net148),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_otrip[2]));
 sky130_fd_sc_hd__clkbuf_8 output149 (.A(net149),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_rc_dis));
 sky130_fd_sc_hd__clkbuf_8 output150 (.A(net150),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_rc_ena));
 sky130_fd_sc_hd__clkbuf_8 output151 (.A(net151),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_vtrip[0]));
 sky130_fd_sc_hd__clkbuf_8 output152 (.A(net152),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_vtrip[1]));
 sky130_fd_sc_hd__clkbuf_8 output153 (.A(net153),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(brownout_vtrip[2]));
 sky130_fd_sc_hd__clkbuf_8 output154 (.A(net154),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_ena));
 sky130_fd_sc_hd__clkbuf_8 output155 (.A(net155),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_hyst[0]));
 sky130_fd_sc_hd__clkbuf_8 output156 (.A(net156),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_hyst[1]));
 sky130_fd_sc_hd__clkbuf_8 output157 (.A(net157),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output158 (.A(net158),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_dac1));
 sky130_fd_sc_hd__clkbuf_8 output159 (.A(net159),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_gpio1_4[0]));
 sky130_fd_sc_hd__clkbuf_8 output160 (.A(net160),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_gpio1_4[1]));
 sky130_fd_sc_hd__clkbuf_8 output161 (.A(net161),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_gpio6_3[0]));
 sky130_fd_sc_hd__clkbuf_8 output162 (.A(net162),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_gpio6_3[1]));
 sky130_fd_sc_hd__clkbuf_8 output163 (.A(net163),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output164 (.A(net164),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output165 (.A(net165),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_vbgsc));
 sky130_fd_sc_hd__clkbuf_8 output166 (.A(net166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output167 (.A(net167),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output168 (.A(net168),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_dac0));
 sky130_fd_sc_hd__clkbuf_8 output169 (.A(net169),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_gpio1_5[0]));
 sky130_fd_sc_hd__clkbuf_8 output170 (.A(net170),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_gpio1_5[1]));
 sky130_fd_sc_hd__clkbuf_8 output171 (.A(net171),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_gpio6_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output172 (.A(net172),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_gpio6_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output173 (.A(net173),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output174 (.A(net174),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output175 (.A(net175),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_tempsense));
 sky130_fd_sc_hd__clkbuf_8 output176 (.A(net176),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_vbgtc));
 sky130_fd_sc_hd__clkbuf_8 output177 (.A(net177),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output178 (.A(net178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_trim[0]));
 sky130_fd_sc_hd__clkbuf_8 output179 (.A(net179),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_trim[1]));
 sky130_fd_sc_hd__clkbuf_8 output180 (.A(net180),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_trim[2]));
 sky130_fd_sc_hd__clkbuf_8 output181 (.A(net181),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_trim[3]));
 sky130_fd_sc_hd__clkbuf_8 output182 (.A(net182),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_trim[4]));
 sky130_fd_sc_hd__clkbuf_8 output183 (.A(net183),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(comp_trim[5]));
 sky130_fd_sc_hd__clkbuf_8 output184 (.A(net184),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac0_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output185 (.A(net185),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac0_to_user));
 sky130_fd_sc_hd__clkbuf_8 output186 (.A(net186),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac1_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output187 (.A(net187),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac1_to_user));
 sky130_fd_sc_hd__clkbuf_8 output188 (.A(net188),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac_refh_to_gpio1_1[0]));
 sky130_fd_sc_hd__clkbuf_8 output189 (.A(net189),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac_refh_to_gpio1_1[1]));
 sky130_fd_sc_hd__clkbuf_8 output190 (.A(net190),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac_refl_to_gpio1_0[0]));
 sky130_fd_sc_hd__clkbuf_8 output191 (.A(net191),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(dac_refl_to_gpio1_0[1]));
 sky130_fd_sc_hd__clkbuf_8 output192 (.A(net192),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_ena));
 sky130_fd_sc_hd__clkbuf_8 output193 (.A(net193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_ref_select));
 sky130_fd_sc_hd__clkbuf_8 output194 (.A(net194),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_snk_ena[0]));
 sky130_fd_sc_hd__clkbuf_8 output195 (.A(net195),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_snk_ena[1]));
 sky130_fd_sc_hd__clkbuf_8 output196 (.A(net196),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_snk_ena[2]));
 sky130_fd_sc_hd__clkbuf_8 output197 (.A(net197),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_snk_ena[3]));
 sky130_fd_sc_hd__clkbuf_8 output198 (.A(net198),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[0]));
 sky130_fd_sc_hd__clkbuf_8 output199 (.A(net199),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[10]));
 sky130_fd_sc_hd__clkbuf_8 output200 (.A(net200),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[11]));
 sky130_fd_sc_hd__clkbuf_8 output201 (.A(net201),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[12]));
 sky130_fd_sc_hd__clkbuf_8 output202 (.A(net202),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[13]));
 sky130_fd_sc_hd__clkbuf_8 output203 (.A(net203),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[14]));
 sky130_fd_sc_hd__clkbuf_8 output204 (.A(net204),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[15]));
 sky130_fd_sc_hd__clkbuf_8 output205 (.A(net205),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[16]));
 sky130_fd_sc_hd__clkbuf_8 output206 (.A(net206),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[17]));
 sky130_fd_sc_hd__clkbuf_8 output207 (.A(net207),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[18]));
 sky130_fd_sc_hd__clkbuf_8 output208 (.A(net208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[19]));
 sky130_fd_sc_hd__clkbuf_8 output209 (.A(net209),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[1]));
 sky130_fd_sc_hd__clkbuf_8 output210 (.A(net210),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[20]));
 sky130_fd_sc_hd__clkbuf_8 output211 (.A(net211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[21]));
 sky130_fd_sc_hd__clkbuf_8 output212 (.A(net212),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[22]));
 sky130_fd_sc_hd__clkbuf_8 output213 (.A(net213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[23]));
 sky130_fd_sc_hd__clkbuf_8 output214 (.A(net214),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[2]));
 sky130_fd_sc_hd__clkbuf_8 output215 (.A(net215),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[3]));
 sky130_fd_sc_hd__clkbuf_8 output216 (.A(net216),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[4]));
 sky130_fd_sc_hd__clkbuf_8 output217 (.A(net217),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[5]));
 sky130_fd_sc_hd__clkbuf_8 output218 (.A(net218),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[6]));
 sky130_fd_sc_hd__clkbuf_8 output219 (.A(net219),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[7]));
 sky130_fd_sc_hd__clkbuf_8 output220 (.A(net220),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[8]));
 sky130_fd_sc_hd__clkbuf_8 output221 (.A(net221),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_src_ena[9]));
 sky130_fd_sc_hd__clkbuf_8 output222 (.A(net222),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_test_to_gpio1_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output223 (.A(net223),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ibias_test_to_gpio1_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output224 (.A(net224),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_ena));
 sky130_fd_sc_hd__clkbuf_8 output225 (.A(net225),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_to_gpio1_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output226 (.A(net226),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_to_gpio1_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output227 (.A(net227),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_to_gpio1_3[0]));
 sky130_fd_sc_hd__clkbuf_8 output228 (.A(net228),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_to_gpio1_3[1]));
 sky130_fd_sc_hd__clkbuf_8 output229 (.A(net229),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[0]));
 sky130_fd_sc_hd__clkbuf_8 output230 (.A(net230),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[10]));
 sky130_fd_sc_hd__clkbuf_8 output231 (.A(net231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[11]));
 sky130_fd_sc_hd__clkbuf_8 output232 (.A(net232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[1]));
 sky130_fd_sc_hd__clkbuf_8 output233 (.A(net233),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[2]));
 sky130_fd_sc_hd__clkbuf_8 output234 (.A(net234),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[3]));
 sky130_fd_sc_hd__clkbuf_8 output235 (.A(net235),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[4]));
 sky130_fd_sc_hd__clkbuf_8 output236 (.A(net236),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[5]));
 sky130_fd_sc_hd__clkbuf_8 output237 (.A(net237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[6]));
 sky130_fd_sc_hd__clkbuf_8 output238 (.A(net238),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[7]));
 sky130_fd_sc_hd__clkbuf_8 output239 (.A(net239),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[8]));
 sky130_fd_sc_hd__clkbuf_8 output240 (.A(net240),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(idac_value[9]));
 sky130_fd_sc_hd__clkbuf_8 output241 (.A(net241),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ldo_ena));
 sky130_fd_sc_hd__clkbuf_8 output242 (.A(net242),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ldo_ref_sel));
 sky130_fd_sc_hd__clkbuf_8 output243 (.A(net243),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_ena));
 sky130_fd_sc_hd__clkbuf_8 output244 (.A(net244),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_amuxbusB));
 sky130_fd_sc_hd__clkbuf_8 output245 (.A(net245),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output246 (.A(net246),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_dac1));
 sky130_fd_sc_hd__clkbuf_8 output247 (.A(net247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_gpio2_0[0]));
 sky130_fd_sc_hd__clkbuf_8 output248 (.A(net248),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_gpio2_0[1]));
 sky130_fd_sc_hd__clkbuf_8 output249 (.A(net249),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_gpio5_3[0]));
 sky130_fd_sc_hd__clkbuf_8 output250 (.A(net250),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_gpio5_3[1]));
 sky130_fd_sc_hd__clkbuf_8 output251 (.A(net251),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output252 (.A(net252),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_rheostat_tap));
 sky130_fd_sc_hd__clkbuf_8 output253 (.A(net253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output254 (.A(net254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output255 (.A(net255),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_vbgtc));
 sky130_fd_sc_hd__clkbuf_8 output256 (.A(net256),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output257 (.A(net257),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_amuxbusA));
 sky130_fd_sc_hd__clkbuf_8 output258 (.A(net258),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output259 (.A(net259),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_dac0));
 sky130_fd_sc_hd__clkbuf_8 output260 (.A(net260),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_gpio2_1[0]));
 sky130_fd_sc_hd__clkbuf_8 output261 (.A(net261),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_gpio2_1[1]));
 sky130_fd_sc_hd__clkbuf_8 output262 (.A(net262),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_gpio5_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output263 (.A(net263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_gpio5_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output264 (.A(net264),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output265 (.A(net265),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output266 (.A(net266),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output267 (.A(net267),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_tempsense));
 sky130_fd_sc_hd__clkbuf_8 output268 (.A(net268),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output269 (.A(net269),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_adc0[0]));
 sky130_fd_sc_hd__clkbuf_8 output270 (.A(net270),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_adc0[1]));
 sky130_fd_sc_hd__clkbuf_8 output271 (.A(net271),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_amuxbusB[0]));
 sky130_fd_sc_hd__clkbuf_8 output272 (.A(net272),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_amuxbusB[1]));
 sky130_fd_sc_hd__clkbuf_8 output273 (.A(net273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_analog1[0]));
 sky130_fd_sc_hd__clkbuf_8 output274 (.A(net274),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_analog1[1]));
 sky130_fd_sc_hd__clkbuf_8 output275 (.A(net275),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_comp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output276 (.A(net276),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_comp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output277 (.A(net277),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio3_1[0]));
 sky130_fd_sc_hd__clkbuf_8 output278 (.A(net278),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio3_1[1]));
 sky130_fd_sc_hd__clkbuf_8 output279 (.A(net279),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio3_5[0]));
 sky130_fd_sc_hd__clkbuf_8 output280 (.A(net280),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio3_5[1]));
 sky130_fd_sc_hd__clkbuf_8 output281 (.A(net281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio4_1[0]));
 sky130_fd_sc_hd__clkbuf_8 output282 (.A(net282),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio4_1[1]));
 sky130_fd_sc_hd__clkbuf_8 output283 (.A(net283),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio4_5[0]));
 sky130_fd_sc_hd__clkbuf_8 output284 (.A(net284),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_gpio4_5[1]));
 sky130_fd_sc_hd__clkbuf_8 output285 (.A(net285),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_ulpcomp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output286 (.A(net286),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_hgbw_opamp_to_ulpcomp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output287 (.A(net287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G1[0]));
 sky130_fd_sc_hd__clkbuf_8 output288 (.A(net288),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G1[1]));
 sky130_fd_sc_hd__clkbuf_8 output289 (.A(net289),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G1[2]));
 sky130_fd_sc_hd__clkbuf_8 output290 (.A(net290),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G1[3]));
 sky130_fd_sc_hd__clkbuf_8 output291 (.A(net291),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G1[4]));
 sky130_fd_sc_hd__clkbuf_8 output292 (.A(net292),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G2[0]));
 sky130_fd_sc_hd__clkbuf_8 output293 (.A(net293),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G2[1]));
 sky130_fd_sc_hd__clkbuf_8 output294 (.A(net294),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G2[2]));
 sky130_fd_sc_hd__clkbuf_8 output295 (.A(net295),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G2[3]));
 sky130_fd_sc_hd__clkbuf_8 output296 (.A(net296),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_G2[4]));
 sky130_fd_sc_hd__clkbuf_8 output297 (.A(net297),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_ena));
 sky130_fd_sc_hd__clkbuf_8 output298 (.A(net298),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_n_to_amuxbusB));
 sky130_fd_sc_hd__clkbuf_8 output299 (.A(net299),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_n_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output300 (.A(net300),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_n_to_gpio5_7[0]));
 sky130_fd_sc_hd__clkbuf_8 output301 (.A(net301),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_n_to_gpio5_7[1]));
 sky130_fd_sc_hd__clkbuf_8 output302 (.A(net302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output303 (.A(net303),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output304 (.A(net304),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output305 (.A(net305),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_amuxbusA));
 sky130_fd_sc_hd__clkbuf_8 output306 (.A(net306),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output307 (.A(net307),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_gpio5_6[0]));
 sky130_fd_sc_hd__clkbuf_8 output308 (.A(net308),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_gpio5_6[1]));
 sky130_fd_sc_hd__clkbuf_8 output309 (.A(net309),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output310 (.A(net310),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output311 (.A(net311),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_tempsense));
 sky130_fd_sc_hd__clkbuf_8 output312 (.A(net312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output313 (.A(net313),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_adc0[0]));
 sky130_fd_sc_hd__clkbuf_8 output314 (.A(net314),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_adc0[1]));
 sky130_fd_sc_hd__clkbuf_8 output315 (.A(net315),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_amuxbusB[0]));
 sky130_fd_sc_hd__clkbuf_8 output316 (.A(net316),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_amuxbusB[1]));
 sky130_fd_sc_hd__clkbuf_8 output317 (.A(net317),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_analog1[0]));
 sky130_fd_sc_hd__clkbuf_8 output318 (.A(net318),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_analog1[1]));
 sky130_fd_sc_hd__clkbuf_8 output319 (.A(net319),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_comp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output320 (.A(net320),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_comp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output321 (.A(net321),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_gpio4_4[0]));
 sky130_fd_sc_hd__clkbuf_8 output322 (.A(net322),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_gpio4_4[1]));
 sky130_fd_sc_hd__clkbuf_8 output323 (.A(net323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_ulpcomp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output324 (.A(net324),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_instramp_to_ulpcomp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output325 (.A(net325),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_ena));
 sky130_fd_sc_hd__clkbuf_8 output326 (.A(net326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_amuxbusB));
 sky130_fd_sc_hd__clkbuf_8 output327 (.A(net327),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output328 (.A(net328),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_dac1));
 sky130_fd_sc_hd__clkbuf_8 output329 (.A(net329),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_gpio5_5[0]));
 sky130_fd_sc_hd__clkbuf_8 output330 (.A(net330),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_gpio5_5[1]));
 sky130_fd_sc_hd__clkbuf_8 output331 (.A(net331),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output332 (.A(net332),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_rheostat_tap));
 sky130_fd_sc_hd__clkbuf_8 output333 (.A(net333),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output334 (.A(net334),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output335 (.A(net335),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_vbgsc));
 sky130_fd_sc_hd__clkbuf_8 output336 (.A(net336),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output337 (.A(net337),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_amuxbusA));
 sky130_fd_sc_hd__clkbuf_8 output338 (.A(net338),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output339 (.A(net339),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_dac0));
 sky130_fd_sc_hd__clkbuf_8 output340 (.A(net340),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_gpio5_4[0]));
 sky130_fd_sc_hd__clkbuf_8 output341 (.A(net341),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_gpio5_4[1]));
 sky130_fd_sc_hd__clkbuf_8 output342 (.A(net342),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output343 (.A(net343),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output344 (.A(net344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output345 (.A(net345),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output346 (.A(net346),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_adc1[0]));
 sky130_fd_sc_hd__clkbuf_8 output347 (.A(net347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_adc1[1]));
 sky130_fd_sc_hd__clkbuf_8 output348 (.A(net348),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_amuxbusA[0]));
 sky130_fd_sc_hd__clkbuf_8 output349 (.A(net349),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_amuxbusA[1]));
 sky130_fd_sc_hd__clkbuf_8 output350 (.A(net350),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_analog0[0]));
 sky130_fd_sc_hd__clkbuf_8 output351 (.A(net351),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_analog0[1]));
 sky130_fd_sc_hd__clkbuf_8 output352 (.A(net352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_comp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output353 (.A(net353),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_comp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output354 (.A(net354),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_gpio3_4[0]));
 sky130_fd_sc_hd__clkbuf_8 output355 (.A(net355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_gpio3_4[1]));
 sky130_fd_sc_hd__clkbuf_8 output356 (.A(net356),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_gpio4_0[0]));
 sky130_fd_sc_hd__clkbuf_8 output357 (.A(net357),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_gpio4_0[1]));
 sky130_fd_sc_hd__clkbuf_8 output358 (.A(net358),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_ulpcomp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output359 (.A(net359),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_lp_opamp_to_ulpcomp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output360 (.A(net360),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[0]));
 sky130_fd_sc_hd__clkbuf_8 output361 (.A(net361),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[1]));
 sky130_fd_sc_hd__clkbuf_8 output362 (.A(net362),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[2]));
 sky130_fd_sc_hd__clkbuf_8 output363 (.A(net363),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[3]));
 sky130_fd_sc_hd__clkbuf_8 output364 (.A(net364),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[4]));
 sky130_fd_sc_hd__clkbuf_8 output365 (.A(net365),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[5]));
 sky130_fd_sc_hd__clkbuf_8 output366 (.A(net366),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[6]));
 sky130_fd_sc_hd__clkbuf_8 output367 (.A(net367),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat1_b[7]));
 sky130_fd_sc_hd__clkbuf_8 output368 (.A(net368),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[0]));
 sky130_fd_sc_hd__clkbuf_8 output369 (.A(net369),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[1]));
 sky130_fd_sc_hd__clkbuf_8 output370 (.A(net370),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[2]));
 sky130_fd_sc_hd__clkbuf_8 output371 (.A(net371),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[3]));
 sky130_fd_sc_hd__clkbuf_8 output372 (.A(net372),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[4]));
 sky130_fd_sc_hd__clkbuf_8 output373 (.A(net373),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[5]));
 sky130_fd_sc_hd__clkbuf_8 output374 (.A(net374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[6]));
 sky130_fd_sc_hd__clkbuf_8 output375 (.A(net375),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_rheostat2_b[7]));
 sky130_fd_sc_hd__clkbuf_8 output376 (.A(net376),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(left_vref_to_user));
 sky130_fd_sc_hd__clkbuf_8 output377 (.A(net377),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(overvoltage_ena));
 sky130_fd_sc_hd__clkbuf_8 output378 (.A(net378),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(overvoltage_trim[0]));
 sky130_fd_sc_hd__clkbuf_8 output379 (.A(net379),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(overvoltage_trim[1]));
 sky130_fd_sc_hd__clkbuf_8 output380 (.A(net380),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(overvoltage_trim[2]));
 sky130_fd_sc_hd__clkbuf_8 output381 (.A(net381),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(overvoltage_trim[3]));
 sky130_fd_sc_hd__clkbuf_8 output382 (.A(net382),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_ena));
 sky130_fd_sc_hd__clkbuf_8 output383 (.A(net383),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[0]));
 sky130_fd_sc_hd__clkbuf_8 output384 (.A(net384),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[10]));
 sky130_fd_sc_hd__clkbuf_8 output385 (.A(net385),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[11]));
 sky130_fd_sc_hd__clkbuf_8 output386 (.A(net386),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[1]));
 sky130_fd_sc_hd__clkbuf_8 output387 (.A(net387),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[2]));
 sky130_fd_sc_hd__clkbuf_8 output388 (.A(net388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[3]));
 sky130_fd_sc_hd__clkbuf_8 output389 (.A(net389),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[4]));
 sky130_fd_sc_hd__clkbuf_8 output390 (.A(net390),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[5]));
 sky130_fd_sc_hd__clkbuf_8 output391 (.A(net391),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[6]));
 sky130_fd_sc_hd__clkbuf_8 output392 (.A(net392),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[7]));
 sky130_fd_sc_hd__clkbuf_8 output393 (.A(net393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[8]));
 sky130_fd_sc_hd__clkbuf_8 output394 (.A(net394),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac0_value[9]));
 sky130_fd_sc_hd__clkbuf_8 output395 (.A(net395),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_ena));
 sky130_fd_sc_hd__clkbuf_8 output396 (.A(net396),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[0]));
 sky130_fd_sc_hd__clkbuf_8 output397 (.A(net397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[10]));
 sky130_fd_sc_hd__clkbuf_8 output398 (.A(net398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[11]));
 sky130_fd_sc_hd__clkbuf_8 output399 (.A(net399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[1]));
 sky130_fd_sc_hd__clkbuf_8 output400 (.A(net400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[2]));
 sky130_fd_sc_hd__clkbuf_8 output401 (.A(net401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[3]));
 sky130_fd_sc_hd__clkbuf_8 output402 (.A(net402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[4]));
 sky130_fd_sc_hd__clkbuf_8 output403 (.A(net403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[5]));
 sky130_fd_sc_hd__clkbuf_8 output404 (.A(net404),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[6]));
 sky130_fd_sc_hd__clkbuf_8 output405 (.A(net405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[7]));
 sky130_fd_sc_hd__clkbuf_8 output406 (.A(net406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[8]));
 sky130_fd_sc_hd__clkbuf_8 output407 (.A(net407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(rdac1_value[9]));
 sky130_fd_sc_hd__clkbuf_8 output408 (.A(net408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_ena));
 sky130_fd_sc_hd__clkbuf_8 output409 (.A(net409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_amuxbusB));
 sky130_fd_sc_hd__clkbuf_8 output410 (.A(net410),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output411 (.A(net411),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_dac1));
 sky130_fd_sc_hd__clkbuf_8 output412 (.A(net412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_gpio2_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output413 (.A(net413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_gpio2_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output414 (.A(net414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_gpio5_1[0]));
 sky130_fd_sc_hd__clkbuf_8 output415 (.A(net415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_gpio5_1[1]));
 sky130_fd_sc_hd__clkbuf_8 output416 (.A(net416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output417 (.A(net417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_rheostat_tap));
 sky130_fd_sc_hd__clkbuf_8 output418 (.A(net418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output419 (.A(net419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output420 (.A(net420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_vbgsc));
 sky130_fd_sc_hd__clkbuf_8 output421 (.A(net421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output422 (.A(net422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_amuxbusA));
 sky130_fd_sc_hd__clkbuf_8 output423 (.A(net423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output424 (.A(net424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_dac0));
 sky130_fd_sc_hd__clkbuf_8 output425 (.A(net425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_gpio2_3[0]));
 sky130_fd_sc_hd__clkbuf_8 output426 (.A(net426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_gpio2_3[1]));
 sky130_fd_sc_hd__clkbuf_8 output427 (.A(net427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_gpio5_0[0]));
 sky130_fd_sc_hd__clkbuf_8 output428 (.A(net428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_gpio5_0[1]));
 sky130_fd_sc_hd__clkbuf_8 output429 (.A(net429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output430 (.A(net430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output431 (.A(net431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output432 (.A(net432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output433 (.A(net433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_adc1[0]));
 sky130_fd_sc_hd__clkbuf_8 output434 (.A(net434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_adc1[1]));
 sky130_fd_sc_hd__clkbuf_8 output435 (.A(net435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_amuxbusA[0]));
 sky130_fd_sc_hd__clkbuf_8 output436 (.A(net436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_amuxbusA[1]));
 sky130_fd_sc_hd__clkbuf_8 output437 (.A(net437),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_analog0[0]));
 sky130_fd_sc_hd__clkbuf_8 output438 (.A(net438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_analog0[1]));
 sky130_fd_sc_hd__clkbuf_8 output439 (.A(net439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_comp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output440 (.A(net440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_comp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output441 (.A(net441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio3_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output442 (.A(net442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio3_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output443 (.A(net443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio3_6[0]));
 sky130_fd_sc_hd__clkbuf_8 output444 (.A(net444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio3_6[1]));
 sky130_fd_sc_hd__clkbuf_8 output445 (.A(net445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio4_2[0]));
 sky130_fd_sc_hd__clkbuf_8 output446 (.A(net446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio4_2[1]));
 sky130_fd_sc_hd__clkbuf_8 output447 (.A(net447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio4_6[0]));
 sky130_fd_sc_hd__clkbuf_8 output448 (.A(net448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_gpio4_6[1]));
 sky130_fd_sc_hd__clkbuf_8 output449 (.A(net449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_ulpcomp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output450 (.A(net450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_hgbw_opamp_to_ulpcomp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output451 (.A(net451),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G1[0]));
 sky130_fd_sc_hd__clkbuf_8 output452 (.A(net452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G1[1]));
 sky130_fd_sc_hd__clkbuf_8 output453 (.A(net453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G1[2]));
 sky130_fd_sc_hd__clkbuf_8 output454 (.A(net454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G1[3]));
 sky130_fd_sc_hd__clkbuf_8 output455 (.A(net455),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G1[4]));
 sky130_fd_sc_hd__clkbuf_8 output456 (.A(net456),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G2[0]));
 sky130_fd_sc_hd__clkbuf_8 output457 (.A(net457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G2[1]));
 sky130_fd_sc_hd__clkbuf_8 output458 (.A(net458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G2[2]));
 sky130_fd_sc_hd__clkbuf_8 output459 (.A(net459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G2[3]));
 sky130_fd_sc_hd__clkbuf_8 output460 (.A(net460),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_G2[4]));
 sky130_fd_sc_hd__clkbuf_8 output461 (.A(net461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_ena));
 sky130_fd_sc_hd__clkbuf_8 output462 (.A(net462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_n_to_amuxbusB));
 sky130_fd_sc_hd__clkbuf_8 output463 (.A(net463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_n_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output464 (.A(net464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_n_to_gpio2_6[0]));
 sky130_fd_sc_hd__clkbuf_8 output465 (.A(net465),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_n_to_gpio2_6[1]));
 sky130_fd_sc_hd__clkbuf_8 output466 (.A(net466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output467 (.A(net467),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output468 (.A(net468),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output469 (.A(net469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_amuxbusA));
 sky130_fd_sc_hd__clkbuf_8 output470 (.A(net470),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output471 (.A(net471),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_gpio2_7[0]));
 sky130_fd_sc_hd__clkbuf_8 output472 (.A(net472),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_gpio2_7[1]));
 sky130_fd_sc_hd__clkbuf_8 output473 (.A(net473),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output474 (.A(net474),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output475 (.A(net475),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_tempsense));
 sky130_fd_sc_hd__clkbuf_8 output476 (.A(net476),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output477 (.A(net477),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_adc1[0]));
 sky130_fd_sc_hd__clkbuf_8 output478 (.A(net478),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_adc1[1]));
 sky130_fd_sc_hd__clkbuf_8 output479 (.A(net479),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_amuxbusA[0]));
 sky130_fd_sc_hd__clkbuf_8 output480 (.A(net480),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_amuxbusA[1]));
 sky130_fd_sc_hd__clkbuf_8 output481 (.A(net481),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_analog0[0]));
 sky130_fd_sc_hd__clkbuf_8 output482 (.A(net482),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_analog0[1]));
 sky130_fd_sc_hd__clkbuf_8 output483 (.A(net483),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_comp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output484 (.A(net484),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_comp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output485 (.A(net485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_gpio3_0[0]));
 sky130_fd_sc_hd__clkbuf_8 output486 (.A(net486),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_gpio3_0[1]));
 sky130_fd_sc_hd__clkbuf_8 output487 (.A(net487),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_ulpcomp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output488 (.A(net488),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_instramp_to_ulpcomp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output489 (.A(net489),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_ena));
 sky130_fd_sc_hd__clkbuf_8 output490 (.A(net490),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_amuxbusB));
 sky130_fd_sc_hd__clkbuf_8 output491 (.A(net491),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output492 (.A(net492),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_dac1));
 sky130_fd_sc_hd__clkbuf_8 output493 (.A(net493),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_gpio2_4[0]));
 sky130_fd_sc_hd__clkbuf_8 output494 (.A(net494),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_gpio2_4[1]));
 sky130_fd_sc_hd__clkbuf_8 output495 (.A(net495),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output496 (.A(net496),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_rheostat_tap));
 sky130_fd_sc_hd__clkbuf_8 output497 (.A(net497),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output498 (.A(net498),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output499 (.A(net499),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_vbgtc));
 sky130_fd_sc_hd__clkbuf_8 output500 (.A(net500),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output501 (.A(net501),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_amuxbusA));
 sky130_fd_sc_hd__clkbuf_8 output502 (.A(net502),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output503 (.A(net503),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_dac0));
 sky130_fd_sc_hd__clkbuf_8 output504 (.A(net504),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_gpio2_5[0]));
 sky130_fd_sc_hd__clkbuf_8 output505 (.A(net505),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_gpio2_5[1]));
 sky130_fd_sc_hd__clkbuf_8 output506 (.A(net506),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output507 (.A(net507),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_rheostat_out));
 sky130_fd_sc_hd__clkbuf_8 output508 (.A(net508),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output509 (.A(net509),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_tempsense));
 sky130_fd_sc_hd__clkbuf_8 output510 (.A(net510),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output511 (.A(net511),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_adc0[0]));
 sky130_fd_sc_hd__clkbuf_8 output512 (.A(net512),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_adc0[1]));
 sky130_fd_sc_hd__clkbuf_8 output513 (.A(net513),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_amuxbusB[0]));
 sky130_fd_sc_hd__clkbuf_8 output514 (.A(net514),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_amuxbusB[1]));
 sky130_fd_sc_hd__clkbuf_8 output515 (.A(net515),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_analog1[0]));
 sky130_fd_sc_hd__clkbuf_8 output516 (.A(net516),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_analog1[1]));
 sky130_fd_sc_hd__clkbuf_8 output517 (.A(net517),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_comp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output518 (.A(net518),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_comp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output519 (.A(net519),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio3_3[0]));
 sky130_fd_sc_hd__clkbuf_8 output520 (.A(net520),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio3_3[1]));
 sky130_fd_sc_hd__clkbuf_8 output521 (.A(net521),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio3_7[0]));
 sky130_fd_sc_hd__clkbuf_8 output522 (.A(net522),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio3_7[1]));
 sky130_fd_sc_hd__clkbuf_8 output523 (.A(net523),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio4_3[0]));
 sky130_fd_sc_hd__clkbuf_8 output524 (.A(net524),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio4_3[1]));
 sky130_fd_sc_hd__clkbuf_8 output525 (.A(net525),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio4_7[0]));
 sky130_fd_sc_hd__clkbuf_8 output526 (.A(net526),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_gpio4_7[1]));
 sky130_fd_sc_hd__clkbuf_8 output527 (.A(net527),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_ulpcomp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output528 (.A(net528),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_lp_opamp_to_ulpcomp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output529 (.A(net529),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[0]));
 sky130_fd_sc_hd__clkbuf_8 output530 (.A(net530),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[1]));
 sky130_fd_sc_hd__clkbuf_8 output531 (.A(net531),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[2]));
 sky130_fd_sc_hd__clkbuf_8 output532 (.A(net532),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[3]));
 sky130_fd_sc_hd__clkbuf_8 output533 (.A(net533),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[4]));
 sky130_fd_sc_hd__clkbuf_8 output534 (.A(net534),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[5]));
 sky130_fd_sc_hd__clkbuf_8 output535 (.A(net535),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[6]));
 sky130_fd_sc_hd__clkbuf_8 output536 (.A(net536),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat1_b[7]));
 sky130_fd_sc_hd__clkbuf_8 output537 (.A(net537),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[0]));
 sky130_fd_sc_hd__clkbuf_8 output538 (.A(net538),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[1]));
 sky130_fd_sc_hd__clkbuf_8 output539 (.A(net539),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[2]));
 sky130_fd_sc_hd__clkbuf_8 output540 (.A(net540),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[3]));
 sky130_fd_sc_hd__clkbuf_8 output541 (.A(net541),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[4]));
 sky130_fd_sc_hd__clkbuf_8 output542 (.A(net542),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[5]));
 sky130_fd_sc_hd__clkbuf_8 output543 (.A(net543),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[6]));
 sky130_fd_sc_hd__clkbuf_8 output544 (.A(net544),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_rheostat2_b[7]));
 sky130_fd_sc_hd__clkbuf_8 output545 (.A(net545),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(right_vref_to_user));
 sky130_fd_sc_hd__clkbuf_8 output546 (.A(net546),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(sio0_connect[0]));
 sky130_fd_sc_hd__clkbuf_8 output547 (.A(net547),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(sio0_connect[1]));
 sky130_fd_sc_hd__clkbuf_8 output548 (.A(net548),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(sio1_connect[0]));
 sky130_fd_sc_hd__clkbuf_8 output549 (.A(net549),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(sio1_connect[1]));
 sky130_fd_sc_hd__clkbuf_8 output550 (.A(net550),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(tempsense_ena));
 sky130_fd_sc_hd__clkbuf_8 output551 (.A(net551),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(tempsense_sel));
 sky130_fd_sc_hd__clkbuf_8 output552 (.A(net552),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(tempsense_to_user));
 sky130_fd_sc_hd__clkbuf_8 output553 (.A(net553),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_clk));
 sky130_fd_sc_hd__clkbuf_8 output554 (.A(net554),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_ena));
 sky130_fd_sc_hd__clkbuf_8 output555 (.A(net555),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_analog0));
 sky130_fd_sc_hd__clkbuf_8 output556 (.A(net556),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_dac1));
 sky130_fd_sc_hd__clkbuf_8 output557 (.A(net557),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_gpio1_6[0]));
 sky130_fd_sc_hd__clkbuf_8 output558 (.A(net558),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_gpio1_6[1]));
 sky130_fd_sc_hd__clkbuf_8 output559 (.A(net559),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_gpio6_1[0]));
 sky130_fd_sc_hd__clkbuf_8 output560 (.A(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_gpio6_1[1]));
 sky130_fd_sc_hd__clkbuf_8 output561 (.A(net561),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_right_vref));
 sky130_fd_sc_hd__clkbuf_8 output562 (.A(net562),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_sio1));
 sky130_fd_sc_hd__clkbuf_8 output563 (.A(net563),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_vbgsc));
 sky130_fd_sc_hd__clkbuf_8 output564 (.A(net564),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_n_to_vinref));
 sky130_fd_sc_hd__clkbuf_8 output565 (.A(net565),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_analog1));
 sky130_fd_sc_hd__clkbuf_8 output566 (.A(net566),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_dac0));
 sky130_fd_sc_hd__clkbuf_8 output567 (.A(net567),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_gpio1_7[0]));
 sky130_fd_sc_hd__clkbuf_8 output568 (.A(net568),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_gpio1_7[1]));
 sky130_fd_sc_hd__clkbuf_8 output569 (.A(net569),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_gpio6_0[0]));
 sky130_fd_sc_hd__clkbuf_8 output570 (.A(net570),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_gpio6_0[1]));
 sky130_fd_sc_hd__clkbuf_8 output571 (.A(net571),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_left_vref));
 sky130_fd_sc_hd__clkbuf_8 output572 (.A(net572),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_sio0));
 sky130_fd_sc_hd__clkbuf_8 output573 (.A(net573),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_tempsense));
 sky130_fd_sc_hd__clkbuf_8 output574 (.A(net574),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_vbgtc));
 sky130_fd_sc_hd__clkbuf_8 output575 (.A(net575),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(ulpcomp_p_to_voutref));
 sky130_fd_sc_hd__clkbuf_8 output576 (.A(net576),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_adc0[0]));
 sky130_fd_sc_hd__clkbuf_8 output577 (.A(net577),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_adc0[1]));
 sky130_fd_sc_hd__clkbuf_8 output578 (.A(net578),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_adc1[0]));
 sky130_fd_sc_hd__clkbuf_8 output579 (.A(net579),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_adc1[1]));
 sky130_fd_sc_hd__clkbuf_8 output580 (.A(net580),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_comp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output581 (.A(net581),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_comp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output582 (.A(net582),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_comp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output583 (.A(net583),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_comp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output584 (.A(net584),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_ulpcomp_n[0]));
 sky130_fd_sc_hd__clkbuf_8 output585 (.A(net585),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_ulpcomp_n[1]));
 sky130_fd_sc_hd__clkbuf_8 output586 (.A(net586),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_ulpcomp_p[0]));
 sky130_fd_sc_hd__clkbuf_8 output587 (.A(net587),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(user_to_ulpcomp_p[1]));
 sky130_fd_sc_hd__clkbuf_8 output588 (.A(net588),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(vbg_test_to_gpio1_1[0]));
 sky130_fd_sc_hd__clkbuf_8 output589 (.A(net589),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(vbg_test_to_gpio1_1[1]));
 sky130_fd_sc_hd__clkbuf_8 output590 (.A(net590),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(vbgsc_to_user));
 sky130_fd_sc_hd__clkbuf_8 output591 (.A(net591),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(vbgtc_to_user));
 sky130_fd_sc_hd__clkbuf_8 output592 (.A(net592),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(vinref_to_user));
 sky130_fd_sc_hd__clkbuf_8 output593 (.A(net593),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(voutref_to_user));
 sky130_fd_sc_hd__buf_12 fanout594 (.A(n1457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net594));
 sky130_fd_sc_hd__buf_12 fanout595 (.A(n1456),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net595));
 sky130_fd_sc_hd__buf_12 fanout596 (.A(n1454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_8 fanout597 (.A(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net597));
 sky130_fd_sc_hd__clkbuf_8 fanout598 (.A(n1404),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_8 fanout599 (.A(n1400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net599));
 sky130_fd_sc_hd__clkbuf_8 fanout600 (.A(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net600));
 sky130_fd_sc_hd__buf_6 fanout601 (.A(n1396),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net601));
 sky130_fd_sc_hd__clkbuf_8 fanout602 (.A(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net602));
 sky130_fd_sc_hd__buf_8 fanout603 (.A(n1395),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net603));
 sky130_fd_sc_hd__clkbuf_8 fanout604 (.A(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net604));
 sky130_fd_sc_hd__buf_4 fanout605 (.A(n1389),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net605));
 sky130_fd_sc_hd__buf_8 fanout606 (.A(n1466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net606));
 sky130_fd_sc_hd__buf_12 fanout607 (.A(n1022),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_16 fanout608 (.A(n1455),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net608));
 sky130_fd_sc_hd__buf_8 fanout609 (.A(n1403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net609));
 sky130_fd_sc_hd__buf_12 fanout610 (.A(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net610));
 sky130_fd_sc_hd__buf_6 fanout611 (.A(n1399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net611));
 sky130_fd_sc_hd__buf_8 fanout612 (.A(n1012),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net612));
 sky130_fd_sc_hd__buf_8 fanout613 (.A(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net613));
 sky130_fd_sc_hd__buf_6 fanout614 (.A(n1001),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net614));
 sky130_fd_sc_hd__buf_8 fanout615 (.A(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net615));
 sky130_fd_sc_hd__buf_6 fanout616 (.A(n1000),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_16 max_cap617 (.A(n1230),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net617));
 sky130_fd_sc_hd__buf_12 max_cap618 (.A(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net618));
 sky130_fd_sc_hd__buf_12 fanout619 (.A(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net619));
 sky130_fd_sc_hd__buf_12 fanout620 (.A(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net620));
 sky130_fd_sc_hd__buf_12 fanout621 (.A(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net621));
 sky130_fd_sc_hd__buf_12 fanout622 (.A(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net622));
 sky130_fd_sc_hd__buf_6 fanout623 (.A(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net623));
 sky130_fd_sc_hd__clkbuf_16 fanout624 (.A(net49),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net624));
 sky130_fd_sc_hd__buf_6 fanout625 (.A(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net625));
 sky130_fd_sc_hd__buf_6 fanout626 (.A(net48),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net626));
 sky130_fd_sc_hd__buf_12 wire627 (.A(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net627));
 sky130_fd_sc_hd__buf_8 fanout628 (.A(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net628));
 sky130_fd_sc_hd__buf_6 fanout629 (.A(net631),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net629));
 sky130_fd_sc_hd__clkbuf_16 wire630 (.A(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net630));
 sky130_fd_sc_hd__buf_12 wire631 (.A(net47),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net631));
 sky130_fd_sc_hd__buf_8 fanout632 (.A(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net632));
 sky130_fd_sc_hd__buf_8 fanout633 (.A(net46),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net633));
 sky130_fd_sc_hd__buf_8 wire634 (.A(net46),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net634));
 sky130_fd_sc_hd__buf_8 fanout635 (.A(net45),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net635));
 sky130_fd_sc_hd__buf_8 fanout636 (.A(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net636));
 sky130_fd_sc_hd__buf_12 wire637 (.A(net45),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net637));
 sky130_fd_sc_hd__buf_6 fanout638 (.A(net44),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net638));
 sky130_fd_sc_hd__buf_8 fanout639 (.A(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net639));
 sky130_fd_sc_hd__buf_12 wire640 (.A(net44),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net640));
 sky130_fd_sc_hd__buf_8 fanout641 (.A(net643),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net641));
 sky130_fd_sc_hd__buf_6 fanout642 (.A(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net642));
 sky130_fd_sc_hd__buf_6 fanout643 (.A(net43),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net643));
 sky130_fd_sc_hd__buf_12 wire644 (.A(net643),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net644));
 sky130_fd_sc_hd__buf_6 fanout645 (.A(net647),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net645));
 sky130_fd_sc_hd__buf_6 fanout646 (.A(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net646));
 sky130_fd_sc_hd__buf_6 fanout647 (.A(net42),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net647));
 sky130_fd_sc_hd__clkbuf_16 wire648 (.A(net647),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net648));
 sky130_fd_sc_hd__clkbuf_8 fanout649 (.A(net31),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net649));
 sky130_fd_sc_hd__buf_4 fanout650 (.A(net652),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net650));
 sky130_fd_sc_hd__buf_8 fanout651 (.A(net652),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net651));
 sky130_fd_sc_hd__buf_12 wire652 (.A(net31),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net652));
 sky130_fd_sc_hd__buf_8 wire653 (.A(net28),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net653));
 sky130_fd_sc_hd__buf_12 wire654 (.A(net27),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net654));
 sky130_fd_sc_hd__buf_8 wire655 (.A(net26),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net655));
 sky130_fd_sc_hd__buf_12 wire656 (.A(net25),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net656));
 sky130_fd_sc_hd__clkbuf_16 wire657 (.A(net22),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net657));
 sky130_fd_sc_hd__buf_12 fanout658 (.A(net21),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net658));
 sky130_fd_sc_hd__clkbuf_4 fanout659 (.A(net21),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net659));
 sky130_fd_sc_hd__clkbuf_8 fanout660 (.A(net20),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net660));
 sky130_fd_sc_hd__buf_4 fanout661 (.A(net663),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net661));
 sky130_fd_sc_hd__buf_6 fanout662 (.A(net663),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net662));
 sky130_fd_sc_hd__buf_8 wire663 (.A(net20),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net663));
 sky130_fd_sc_hd__clkbuf_8 fanout664 (.A(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net664));
 sky130_fd_sc_hd__clkbuf_8 fanout665 (.A(net666),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_8 fanout666 (.A(net667),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_4 fanout667 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net667));
 sky130_fd_sc_hd__clkbuf_8 fanout668 (.A(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_8 fanout669 (.A(net670),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net669));
 sky130_fd_sc_hd__clkbuf_4 fanout670 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net670));
 sky130_fd_sc_hd__clkbuf_8 fanout671 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net671));
 sky130_fd_sc_hd__clkbuf_4 fanout672 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_8 fanout673 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net673));
 sky130_fd_sc_hd__clkbuf_8 fanout674 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net674));
 sky130_fd_sc_hd__buf_4 fanout675 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_8 fanout676 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_4 fanout677 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_8 fanout678 (.A(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_8 fanout679 (.A(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net679));
 sky130_fd_sc_hd__clkbuf_4 fanout680 (.A(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net680));
 sky130_fd_sc_hd__buf_4 fanout681 (.A(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net681));
 sky130_fd_sc_hd__buf_8 fanout682 (.A(net18),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net682));
 sky130_fd_sc_hd__clkbuf_8 fanout683 (.A(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net683));
 sky130_fd_sc_hd__buf_4 fanout684 (.A(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_8 fanout685 (.A(net686),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_4 fanout686 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_8 fanout687 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net687));
 sky130_fd_sc_hd__buf_4 fanout688 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net688));
 sky130_fd_sc_hd__clkbuf_8 fanout689 (.A(net690),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_8 fanout690 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_8 fanout691 (.A(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net691));
 sky130_fd_sc_hd__clkbuf_8 fanout692 (.A(net693),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net692));
 sky130_fd_sc_hd__buf_4 fanout693 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net693));
 sky130_fd_sc_hd__clkbuf_8 fanout694 (.A(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_8 fanout695 (.A(net696),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net695));
 sky130_fd_sc_hd__buf_4 fanout696 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net696));
 sky130_fd_sc_hd__clkbuf_8 fanout697 (.A(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net697));
 sky130_fd_sc_hd__clkbuf_8 fanout698 (.A(net699),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net698));
 sky130_fd_sc_hd__buf_4 fanout699 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_8 fanout700 (.A(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_8 fanout701 (.A(net702),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_4 fanout702 (.A(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net702));
 sky130_fd_sc_hd__buf_8 fanout703 (.A(net18),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net703));
 sky130_fd_sc_hd__conb_1 U1060_704 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .LO(net704));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_1_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_2_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_3_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_4_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_5_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_6_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_7_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_8_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_9_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_10_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_10_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_11_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_11_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_12_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_12_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_13_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_13_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_14_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_14_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_15_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_15_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_16_PCLK (.A(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_16_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_17_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_17_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_18_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_18_PCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_19_PCLK (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_leaf_19_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_PCLK (.A(PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_0_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_PCLK (.A(clknet_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_1_0__leaf_PCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_PCLK (.A(clknet_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(clknet_1_1__leaf_PCLK));
 sky130_fd_sc_hd__clkinvlp_4 clkload0 (.A(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload3 (.A(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload5 (.A(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload6 (.A(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload7 (.A(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload8 (.A(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload9 (.A(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload10 (.A(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload11 (.A(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload12 (.A(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload13 (.A(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload14 (.A(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload15 (.A(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload16 (.A(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload17 (.A(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__clkbuf_4 clkload18 (.A(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__buf_4 rebuffer1 (.A(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net705));
 sky130_fd_sc_hd__nor2_4 clone2 (.A(net722),
    .B(net709),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(net706));
 sky130_fd_sc_hd__buf_12 rebuffer3 (.A(n1101),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net707));
 sky130_fd_sc_hd__dlymetal6s2s_1 rebuffer4 (.A(net707),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer5 (.A(net707),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net709));
 sky130_fd_sc_hd__buf_4 rebuffer6 (.A(n1122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net710));
 sky130_fd_sc_hd__clkbuf_4 rebuffer7 (.A(n1122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net711));
 sky130_fd_sc_hd__buf_6 rebuffer8 (.A(n1214),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer9 (.A(net712),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net713));
 sky130_fd_sc_hd__buf_2 rebuffer10 (.A(n1416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net714));
 sky130_fd_sc_hd__buf_8 rebuffer11 (.A(n1013),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net715));
 sky130_fd_sc_hd__nor2_4 clone12 (.A(net617),
    .B(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(net716));
 sky130_fd_sc_hd__nor2_4 clone13 (.A(net719),
    .B(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(net717));
 sky130_fd_sc_hd__clkbuf_16 clone14 (.A(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net718));
 sky130_fd_sc_hd__nand2_4 clone15 (.A(n1033),
    .B(n1018),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(net719));
 sky130_fd_sc_hd__nor2_4 clone16 (.A(net722),
    .B(n1127),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(net720));
 sky130_fd_sc_hd__nor2_4 clone17 (.A(net722),
    .B(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .Y(net721));
 sky130_fd_sc_hd__clkbuf_16 clone18 (.A(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0),
    .X(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(PADDR[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(PADDR[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(PADDR[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(PADDR[12]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(PADDR[13]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(PADDR[14]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(PADDR[15]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(PADDR[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(PADDR[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(PADDR[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(PADDR[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(PADDR[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(PADDR[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(PADDR[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(PADDR[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(PADDR[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_PCLK_A (.DIODE(PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(PENABLE),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output62_X (.DIODE(PRDATA[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_X (.DIODE(PRDATA[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_X (.DIODE(PRDATA[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_X (.DIODE(PRDATA[12]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output66_X (.DIODE(PRDATA[13]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_X (.DIODE(PRDATA[14]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_X (.DIODE(PRDATA[15]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_X (.DIODE(PRDATA[16]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_X (.DIODE(PRDATA[17]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_X (.DIODE(PRDATA[18]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_X (.DIODE(PRDATA[19]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_X (.DIODE(PRDATA[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_X (.DIODE(PRDATA[20]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_X (.DIODE(PRDATA[21]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_X (.DIODE(PRDATA[22]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_X (.DIODE(PRDATA[23]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_X (.DIODE(PRDATA[24]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_X (.DIODE(PRDATA[25]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_X (.DIODE(PRDATA[26]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_X (.DIODE(PRDATA[27]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_X (.DIODE(PRDATA[28]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_X (.DIODE(PRDATA[29]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_X (.DIODE(PRDATA[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_X (.DIODE(PRDATA[30]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_X (.DIODE(PRDATA[31]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_X (.DIODE(PRDATA[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_X (.DIODE(PRDATA[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_X (.DIODE(PRDATA[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_X (.DIODE(PRDATA[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_X (.DIODE(PRDATA[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_X (.DIODE(PRDATA[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_X (.DIODE(PRDATA[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1060_Y (.DIODE(PREADY),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(PRESETn),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(PSEL),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(PWDATA[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(PWDATA[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(PWDATA[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(PWDATA[12]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(PWDATA[13]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(PWDATA[14]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(PWDATA[15]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(PWDATA[16]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(PWDATA[17]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(PWDATA[18]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(PWDATA[19]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(PWDATA[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(PWDATA[20]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(PWDATA[21]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(PWDATA[22]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(PWDATA[23]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(PWDATA[24]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(PWDATA[25]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(PWDATA[26]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(PWDATA[27]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(PWDATA[28]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(PWDATA[29]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(PWDATA[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(PWDATA[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(PWDATA[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(PWDATA[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(PWDATA[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(PWDATA[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(PWDATA[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(PWDATA[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(PWRITE),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_X (.DIODE(adc0_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_X (.DIODE(adc0_to_dac0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_X (.DIODE(adc0_to_gpio1_3[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_X (.DIODE(adc0_to_gpio1_3[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_X (.DIODE(adc0_to_gpio6_4[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_X (.DIODE(adc0_to_gpio6_4[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_X (.DIODE(adc0_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_X (.DIODE(adc0_to_tempsense),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_X (.DIODE(adc0_to_vbgtc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_X (.DIODE(adc0_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_X (.DIODE(adc1_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_X (.DIODE(adc1_to_dac1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_X (.DIODE(adc1_to_gpio1_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_X (.DIODE(adc1_to_gpio1_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_X (.DIODE(adc1_to_gpio6_5[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_X (.DIODE(adc1_to_gpio6_5[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_X (.DIODE(adc1_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_X (.DIODE(adc1_to_vbgsc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_X (.DIODE(adc1_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_X (.DIODE(adc_refh_to_gpio6_6[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_X (.DIODE(adc_refh_to_gpio6_6[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_X (.DIODE(adc_refl_to_gpio6_7[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_X (.DIODE(adc_refl_to_gpio6_7[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_X (.DIODE(analog0_connect[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output118_X (.DIODE(analog0_connect[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_X (.DIODE(analog1_connect[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_X (.DIODE(analog1_connect[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_X (.DIODE(audiodac_out_to_analog1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_X (.DIODE(audiodac_out_to_analog1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output123_X (.DIODE(audiodac_outb_to_analog0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_X (.DIODE(audiodac_outb_to_analog0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output125_X (.DIODE(bandgap_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output126_X (.DIODE(bandgap_sel),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output127_X (.DIODE(bandgap_trim[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output128_X (.DIODE(bandgap_trim[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output129_X (.DIODE(bandgap_trim[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output130_X (.DIODE(bandgap_trim[12]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output131_X (.DIODE(bandgap_trim[13]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_X (.DIODE(bandgap_trim[14]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_X (.DIODE(bandgap_trim[15]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output134_X (.DIODE(bandgap_trim[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_X (.DIODE(bandgap_trim[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_X (.DIODE(bandgap_trim[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_X (.DIODE(bandgap_trim[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_X (.DIODE(bandgap_trim[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output139_X (.DIODE(bandgap_trim[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_X (.DIODE(bandgap_trim[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_X (.DIODE(bandgap_trim[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output142_X (.DIODE(bandgap_trim[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output143_X (.DIODE(brownout_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(brownout_filt),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_X (.DIODE(brownout_isrc_sel),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_X (.DIODE(brownout_oneshot),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output146_X (.DIODE(brownout_otrip[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output147_X (.DIODE(brownout_otrip[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_X (.DIODE(brownout_otrip[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_X (.DIODE(brownout_rc_dis),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output150_X (.DIODE(brownout_rc_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(brownout_timeout),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(brownout_unfilt),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output151_X (.DIODE(brownout_vtrip[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output152_X (.DIODE(brownout_vtrip[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output153_X (.DIODE(brownout_vtrip[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(brownout_vunder),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output154_X (.DIODE(comp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_X (.DIODE(comp_hyst[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_X (.DIODE(comp_hyst[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_X (.DIODE(comp_n_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_X (.DIODE(comp_n_to_dac1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_X (.DIODE(comp_n_to_gpio1_4[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_X (.DIODE(comp_n_to_gpio1_4[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_X (.DIODE(comp_n_to_gpio6_3[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_X (.DIODE(comp_n_to_gpio6_3[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_X (.DIODE(comp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_X (.DIODE(comp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_X (.DIODE(comp_n_to_vbgsc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_X (.DIODE(comp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(comp_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output167_X (.DIODE(comp_p_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_X (.DIODE(comp_p_to_dac0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_X (.DIODE(comp_p_to_gpio1_5[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_X (.DIODE(comp_p_to_gpio1_5[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_X (.DIODE(comp_p_to_gpio6_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_X (.DIODE(comp_p_to_gpio6_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output173_X (.DIODE(comp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_X (.DIODE(comp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output175_X (.DIODE(comp_p_to_tempsense),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_X (.DIODE(comp_p_to_vbgtc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_X (.DIODE(comp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_X (.DIODE(comp_trim[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_X (.DIODE(comp_trim[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_X (.DIODE(comp_trim[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_X (.DIODE(comp_trim[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_X (.DIODE(comp_trim[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_X (.DIODE(comp_trim[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_X (.DIODE(dac0_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_X (.DIODE(dac0_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_X (.DIODE(dac1_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_X (.DIODE(dac1_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_X (.DIODE(dac_refh_to_gpio1_1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_X (.DIODE(dac_refh_to_gpio1_1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_X (.DIODE(dac_refl_to_gpio1_0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_X (.DIODE(dac_refl_to_gpio1_0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_X (.DIODE(ibias_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_X (.DIODE(ibias_ref_select),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_X (.DIODE(ibias_snk_ena[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_X (.DIODE(ibias_snk_ena[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_X (.DIODE(ibias_snk_ena[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_X (.DIODE(ibias_snk_ena[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_X (.DIODE(ibias_src_ena[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_X (.DIODE(ibias_src_ena[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output200_X (.DIODE(ibias_src_ena[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_X (.DIODE(ibias_src_ena[12]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output202_X (.DIODE(ibias_src_ena[13]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_X (.DIODE(ibias_src_ena[14]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_X (.DIODE(ibias_src_ena[15]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_X (.DIODE(ibias_src_ena[16]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output206_X (.DIODE(ibias_src_ena[17]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_X (.DIODE(ibias_src_ena[18]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output208_X (.DIODE(ibias_src_ena[19]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output209_X (.DIODE(ibias_src_ena[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_X (.DIODE(ibias_src_ena[20]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output211_X (.DIODE(ibias_src_ena[21]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output212_X (.DIODE(ibias_src_ena[22]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output213_X (.DIODE(ibias_src_ena[23]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output214_X (.DIODE(ibias_src_ena[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output215_X (.DIODE(ibias_src_ena[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output216_X (.DIODE(ibias_src_ena[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output217_X (.DIODE(ibias_src_ena[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output218_X (.DIODE(ibias_src_ena[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output219_X (.DIODE(ibias_src_ena[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output220_X (.DIODE(ibias_src_ena[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output221_X (.DIODE(ibias_src_ena[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output222_X (.DIODE(ibias_test_to_gpio1_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output223_X (.DIODE(ibias_test_to_gpio1_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output224_X (.DIODE(idac_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output225_X (.DIODE(idac_to_gpio1_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output226_X (.DIODE(idac_to_gpio1_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output227_X (.DIODE(idac_to_gpio1_3[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output228_X (.DIODE(idac_to_gpio1_3[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output229_X (.DIODE(idac_value[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output230_X (.DIODE(idac_value[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output231_X (.DIODE(idac_value[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output232_X (.DIODE(idac_value[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output233_X (.DIODE(idac_value[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output234_X (.DIODE(idac_value[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output235_X (.DIODE(idac_value[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output236_X (.DIODE(idac_value[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output237_X (.DIODE(idac_value[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output238_X (.DIODE(idac_value[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output239_X (.DIODE(idac_value[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output240_X (.DIODE(idac_value[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output241_X (.DIODE(ldo_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output242_X (.DIODE(ldo_ref_sel),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output243_X (.DIODE(left_hgbw_opamp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output244_X (.DIODE(left_hgbw_opamp_n_to_amuxbusB),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output245_X (.DIODE(left_hgbw_opamp_n_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output246_X (.DIODE(left_hgbw_opamp_n_to_dac1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output247_X (.DIODE(left_hgbw_opamp_n_to_gpio2_0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output248_X (.DIODE(left_hgbw_opamp_n_to_gpio2_0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output249_X (.DIODE(left_hgbw_opamp_n_to_gpio5_3[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output250_X (.DIODE(left_hgbw_opamp_n_to_gpio5_3[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output251_X (.DIODE(left_hgbw_opamp_n_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output252_X (.DIODE(left_hgbw_opamp_n_to_rheostat_tap),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output253_X (.DIODE(left_hgbw_opamp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output254_X (.DIODE(left_hgbw_opamp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output255_X (.DIODE(left_hgbw_opamp_n_to_vbgtc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output256_X (.DIODE(left_hgbw_opamp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output257_X (.DIODE(left_hgbw_opamp_p_to_amuxbusA),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_X (.DIODE(left_hgbw_opamp_p_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output259_X (.DIODE(left_hgbw_opamp_p_to_dac0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_X (.DIODE(left_hgbw_opamp_p_to_gpio2_1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output261_X (.DIODE(left_hgbw_opamp_p_to_gpio2_1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output262_X (.DIODE(left_hgbw_opamp_p_to_gpio5_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_X (.DIODE(left_hgbw_opamp_p_to_gpio5_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output264_X (.DIODE(left_hgbw_opamp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output265_X (.DIODE(left_hgbw_opamp_p_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output266_X (.DIODE(left_hgbw_opamp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output267_X (.DIODE(left_hgbw_opamp_p_to_tempsense),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output268_X (.DIODE(left_hgbw_opamp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output269_X (.DIODE(left_hgbw_opamp_to_adc0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output270_X (.DIODE(left_hgbw_opamp_to_adc0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output271_X (.DIODE(left_hgbw_opamp_to_amuxbusB[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output272_X (.DIODE(left_hgbw_opamp_to_amuxbusB[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output273_X (.DIODE(left_hgbw_opamp_to_analog1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output274_X (.DIODE(left_hgbw_opamp_to_analog1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_X (.DIODE(left_hgbw_opamp_to_comp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output276_X (.DIODE(left_hgbw_opamp_to_comp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output277_X (.DIODE(left_hgbw_opamp_to_gpio3_1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output278_X (.DIODE(left_hgbw_opamp_to_gpio3_1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output279_X (.DIODE(left_hgbw_opamp_to_gpio3_5[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output280_X (.DIODE(left_hgbw_opamp_to_gpio3_5[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output281_X (.DIODE(left_hgbw_opamp_to_gpio4_1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_X (.DIODE(left_hgbw_opamp_to_gpio4_1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output283_X (.DIODE(left_hgbw_opamp_to_gpio4_5[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output284_X (.DIODE(left_hgbw_opamp_to_gpio4_5[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output285_X (.DIODE(left_hgbw_opamp_to_ulpcomp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output286_X (.DIODE(left_hgbw_opamp_to_ulpcomp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output287_X (.DIODE(left_instramp_G1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output288_X (.DIODE(left_instramp_G1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output289_X (.DIODE(left_instramp_G1[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output290_X (.DIODE(left_instramp_G1[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output291_X (.DIODE(left_instramp_G1[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_X (.DIODE(left_instramp_G2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output293_X (.DIODE(left_instramp_G2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_X (.DIODE(left_instramp_G2[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_X (.DIODE(left_instramp_G2[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_X (.DIODE(left_instramp_G2[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_X (.DIODE(left_instramp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_X (.DIODE(left_instramp_n_to_amuxbusB),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_X (.DIODE(left_instramp_n_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output300_X (.DIODE(left_instramp_n_to_gpio5_7[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output301_X (.DIODE(left_instramp_n_to_gpio5_7[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output302_X (.DIODE(left_instramp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output303_X (.DIODE(left_instramp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output304_X (.DIODE(left_instramp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_X (.DIODE(left_instramp_p_to_amuxbusA),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output306_X (.DIODE(left_instramp_p_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_X (.DIODE(left_instramp_p_to_gpio5_6[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_X (.DIODE(left_instramp_p_to_gpio5_6[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output309_X (.DIODE(left_instramp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output310_X (.DIODE(left_instramp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output311_X (.DIODE(left_instramp_p_to_tempsense),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output312_X (.DIODE(left_instramp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output313_X (.DIODE(left_instramp_to_adc0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output314_X (.DIODE(left_instramp_to_adc0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output315_X (.DIODE(left_instramp_to_amuxbusB[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output316_X (.DIODE(left_instramp_to_amuxbusB[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output317_X (.DIODE(left_instramp_to_analog1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output318_X (.DIODE(left_instramp_to_analog1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output319_X (.DIODE(left_instramp_to_comp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output320_X (.DIODE(left_instramp_to_comp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output321_X (.DIODE(left_instramp_to_gpio4_4[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output322_X (.DIODE(left_instramp_to_gpio4_4[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output323_X (.DIODE(left_instramp_to_ulpcomp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output324_X (.DIODE(left_instramp_to_ulpcomp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output325_X (.DIODE(left_lp_opamp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output326_X (.DIODE(left_lp_opamp_n_to_amuxbusB),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output327_X (.DIODE(left_lp_opamp_n_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output328_X (.DIODE(left_lp_opamp_n_to_dac1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output329_X (.DIODE(left_lp_opamp_n_to_gpio5_5[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output330_X (.DIODE(left_lp_opamp_n_to_gpio5_5[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output331_X (.DIODE(left_lp_opamp_n_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output332_X (.DIODE(left_lp_opamp_n_to_rheostat_tap),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output333_X (.DIODE(left_lp_opamp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output334_X (.DIODE(left_lp_opamp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output335_X (.DIODE(left_lp_opamp_n_to_vbgsc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output336_X (.DIODE(left_lp_opamp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output337_X (.DIODE(left_lp_opamp_p_to_amuxbusA),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output338_X (.DIODE(left_lp_opamp_p_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output339_X (.DIODE(left_lp_opamp_p_to_dac0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output340_X (.DIODE(left_lp_opamp_p_to_gpio5_4[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output341_X (.DIODE(left_lp_opamp_p_to_gpio5_4[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output342_X (.DIODE(left_lp_opamp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output343_X (.DIODE(left_lp_opamp_p_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output344_X (.DIODE(left_lp_opamp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output345_X (.DIODE(left_lp_opamp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output346_X (.DIODE(left_lp_opamp_to_adc1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output347_X (.DIODE(left_lp_opamp_to_adc1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output348_X (.DIODE(left_lp_opamp_to_amuxbusA[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output349_X (.DIODE(left_lp_opamp_to_amuxbusA[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output350_X (.DIODE(left_lp_opamp_to_analog0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output351_X (.DIODE(left_lp_opamp_to_analog0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output352_X (.DIODE(left_lp_opamp_to_comp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output353_X (.DIODE(left_lp_opamp_to_comp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output354_X (.DIODE(left_lp_opamp_to_gpio3_4[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output355_X (.DIODE(left_lp_opamp_to_gpio3_4[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output356_X (.DIODE(left_lp_opamp_to_gpio4_0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output357_X (.DIODE(left_lp_opamp_to_gpio4_0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output358_X (.DIODE(left_lp_opamp_to_ulpcomp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output359_X (.DIODE(left_lp_opamp_to_ulpcomp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output360_X (.DIODE(left_rheostat1_b[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output361_X (.DIODE(left_rheostat1_b[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output362_X (.DIODE(left_rheostat1_b[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output363_X (.DIODE(left_rheostat1_b[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output364_X (.DIODE(left_rheostat1_b[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output365_X (.DIODE(left_rheostat1_b[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output366_X (.DIODE(left_rheostat1_b[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output367_X (.DIODE(left_rheostat1_b[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output368_X (.DIODE(left_rheostat2_b[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output369_X (.DIODE(left_rheostat2_b[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output370_X (.DIODE(left_rheostat2_b[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output371_X (.DIODE(left_rheostat2_b[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output372_X (.DIODE(left_rheostat2_b[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output373_X (.DIODE(left_rheostat2_b[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output374_X (.DIODE(left_rheostat2_b[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output375_X (.DIODE(left_rheostat2_b[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output376_X (.DIODE(left_vref_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output377_X (.DIODE(overvoltage_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(overvoltage_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output378_X (.DIODE(overvoltage_trim[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output379_X (.DIODE(overvoltage_trim[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output380_X (.DIODE(overvoltage_trim[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output381_X (.DIODE(overvoltage_trim[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output382_X (.DIODE(rdac0_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output383_X (.DIODE(rdac0_value[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output384_X (.DIODE(rdac0_value[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output385_X (.DIODE(rdac0_value[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output386_X (.DIODE(rdac0_value[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output387_X (.DIODE(rdac0_value[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output388_X (.DIODE(rdac0_value[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output389_X (.DIODE(rdac0_value[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output390_X (.DIODE(rdac0_value[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output391_X (.DIODE(rdac0_value[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output392_X (.DIODE(rdac0_value[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output393_X (.DIODE(rdac0_value[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output394_X (.DIODE(rdac0_value[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output395_X (.DIODE(rdac1_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output396_X (.DIODE(rdac1_value[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output397_X (.DIODE(rdac1_value[10]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output398_X (.DIODE(rdac1_value[11]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output399_X (.DIODE(rdac1_value[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output400_X (.DIODE(rdac1_value[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output401_X (.DIODE(rdac1_value[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output402_X (.DIODE(rdac1_value[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output403_X (.DIODE(rdac1_value[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output404_X (.DIODE(rdac1_value[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output405_X (.DIODE(rdac1_value[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output406_X (.DIODE(rdac1_value[8]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output407_X (.DIODE(rdac1_value[9]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output408_X (.DIODE(right_hgbw_opamp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output409_X (.DIODE(right_hgbw_opamp_n_to_amuxbusB),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output410_X (.DIODE(right_hgbw_opamp_n_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output411_X (.DIODE(right_hgbw_opamp_n_to_dac1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output412_X (.DIODE(right_hgbw_opamp_n_to_gpio2_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output413_X (.DIODE(right_hgbw_opamp_n_to_gpio2_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output414_X (.DIODE(right_hgbw_opamp_n_to_gpio5_1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output415_X (.DIODE(right_hgbw_opamp_n_to_gpio5_1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output416_X (.DIODE(right_hgbw_opamp_n_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output417_X (.DIODE(right_hgbw_opamp_n_to_rheostat_tap),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output418_X (.DIODE(right_hgbw_opamp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output419_X (.DIODE(right_hgbw_opamp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output420_X (.DIODE(right_hgbw_opamp_n_to_vbgsc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output421_X (.DIODE(right_hgbw_opamp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output422_X (.DIODE(right_hgbw_opamp_p_to_amuxbusA),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output423_X (.DIODE(right_hgbw_opamp_p_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output424_X (.DIODE(right_hgbw_opamp_p_to_dac0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output425_X (.DIODE(right_hgbw_opamp_p_to_gpio2_3[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output426_X (.DIODE(right_hgbw_opamp_p_to_gpio2_3[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output427_X (.DIODE(right_hgbw_opamp_p_to_gpio5_0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output428_X (.DIODE(right_hgbw_opamp_p_to_gpio5_0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output429_X (.DIODE(right_hgbw_opamp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output430_X (.DIODE(right_hgbw_opamp_p_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output431_X (.DIODE(right_hgbw_opamp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output432_X (.DIODE(right_hgbw_opamp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output433_X (.DIODE(right_hgbw_opamp_to_adc1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output434_X (.DIODE(right_hgbw_opamp_to_adc1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output435_X (.DIODE(right_hgbw_opamp_to_amuxbusA[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output436_X (.DIODE(right_hgbw_opamp_to_amuxbusA[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output437_X (.DIODE(right_hgbw_opamp_to_analog0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output438_X (.DIODE(right_hgbw_opamp_to_analog0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output439_X (.DIODE(right_hgbw_opamp_to_comp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output440_X (.DIODE(right_hgbw_opamp_to_comp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output441_X (.DIODE(right_hgbw_opamp_to_gpio3_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output442_X (.DIODE(right_hgbw_opamp_to_gpio3_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output443_X (.DIODE(right_hgbw_opamp_to_gpio3_6[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output444_X (.DIODE(right_hgbw_opamp_to_gpio3_6[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output445_X (.DIODE(right_hgbw_opamp_to_gpio4_2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output446_X (.DIODE(right_hgbw_opamp_to_gpio4_2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output447_X (.DIODE(right_hgbw_opamp_to_gpio4_6[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output448_X (.DIODE(right_hgbw_opamp_to_gpio4_6[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output449_X (.DIODE(right_hgbw_opamp_to_ulpcomp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output450_X (.DIODE(right_hgbw_opamp_to_ulpcomp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output451_X (.DIODE(right_instramp_G1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output452_X (.DIODE(right_instramp_G1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output453_X (.DIODE(right_instramp_G1[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output454_X (.DIODE(right_instramp_G1[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output455_X (.DIODE(right_instramp_G1[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output456_X (.DIODE(right_instramp_G2[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output457_X (.DIODE(right_instramp_G2[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output458_X (.DIODE(right_instramp_G2[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output459_X (.DIODE(right_instramp_G2[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output460_X (.DIODE(right_instramp_G2[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output461_X (.DIODE(right_instramp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output462_X (.DIODE(right_instramp_n_to_amuxbusB),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output463_X (.DIODE(right_instramp_n_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output464_X (.DIODE(right_instramp_n_to_gpio2_6[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output465_X (.DIODE(right_instramp_n_to_gpio2_6[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output466_X (.DIODE(right_instramp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output467_X (.DIODE(right_instramp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output468_X (.DIODE(right_instramp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output469_X (.DIODE(right_instramp_p_to_amuxbusA),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output470_X (.DIODE(right_instramp_p_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output471_X (.DIODE(right_instramp_p_to_gpio2_7[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output472_X (.DIODE(right_instramp_p_to_gpio2_7[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output473_X (.DIODE(right_instramp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output474_X (.DIODE(right_instramp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output475_X (.DIODE(right_instramp_p_to_tempsense),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output476_X (.DIODE(right_instramp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output477_X (.DIODE(right_instramp_to_adc1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output478_X (.DIODE(right_instramp_to_adc1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output479_X (.DIODE(right_instramp_to_amuxbusA[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output480_X (.DIODE(right_instramp_to_amuxbusA[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output481_X (.DIODE(right_instramp_to_analog0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output482_X (.DIODE(right_instramp_to_analog0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output483_X (.DIODE(right_instramp_to_comp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output484_X (.DIODE(right_instramp_to_comp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output485_X (.DIODE(right_instramp_to_gpio3_0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output486_X (.DIODE(right_instramp_to_gpio3_0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output487_X (.DIODE(right_instramp_to_ulpcomp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output488_X (.DIODE(right_instramp_to_ulpcomp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output489_X (.DIODE(right_lp_opamp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output490_X (.DIODE(right_lp_opamp_n_to_amuxbusB),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output491_X (.DIODE(right_lp_opamp_n_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output492_X (.DIODE(right_lp_opamp_n_to_dac1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output493_X (.DIODE(right_lp_opamp_n_to_gpio2_4[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output494_X (.DIODE(right_lp_opamp_n_to_gpio2_4[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output495_X (.DIODE(right_lp_opamp_n_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output496_X (.DIODE(right_lp_opamp_n_to_rheostat_tap),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output497_X (.DIODE(right_lp_opamp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output498_X (.DIODE(right_lp_opamp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output499_X (.DIODE(right_lp_opamp_n_to_vbgtc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output500_X (.DIODE(right_lp_opamp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output501_X (.DIODE(right_lp_opamp_p_to_amuxbusA),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output502_X (.DIODE(right_lp_opamp_p_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output503_X (.DIODE(right_lp_opamp_p_to_dac0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output504_X (.DIODE(right_lp_opamp_p_to_gpio2_5[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output505_X (.DIODE(right_lp_opamp_p_to_gpio2_5[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output506_X (.DIODE(right_lp_opamp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output507_X (.DIODE(right_lp_opamp_p_to_rheostat_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output508_X (.DIODE(right_lp_opamp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output509_X (.DIODE(right_lp_opamp_p_to_tempsense),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output510_X (.DIODE(right_lp_opamp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output511_X (.DIODE(right_lp_opamp_to_adc0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output512_X (.DIODE(right_lp_opamp_to_adc0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output513_X (.DIODE(right_lp_opamp_to_amuxbusB[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output514_X (.DIODE(right_lp_opamp_to_amuxbusB[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output515_X (.DIODE(right_lp_opamp_to_analog1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output516_X (.DIODE(right_lp_opamp_to_analog1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output517_X (.DIODE(right_lp_opamp_to_comp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output518_X (.DIODE(right_lp_opamp_to_comp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output519_X (.DIODE(right_lp_opamp_to_gpio3_3[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output520_X (.DIODE(right_lp_opamp_to_gpio3_3[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output521_X (.DIODE(right_lp_opamp_to_gpio3_7[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output522_X (.DIODE(right_lp_opamp_to_gpio3_7[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output523_X (.DIODE(right_lp_opamp_to_gpio4_3[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output524_X (.DIODE(right_lp_opamp_to_gpio4_3[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output525_X (.DIODE(right_lp_opamp_to_gpio4_7[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output526_X (.DIODE(right_lp_opamp_to_gpio4_7[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output527_X (.DIODE(right_lp_opamp_to_ulpcomp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output528_X (.DIODE(right_lp_opamp_to_ulpcomp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output529_X (.DIODE(right_rheostat1_b[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output530_X (.DIODE(right_rheostat1_b[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output531_X (.DIODE(right_rheostat1_b[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output532_X (.DIODE(right_rheostat1_b[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output533_X (.DIODE(right_rheostat1_b[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output534_X (.DIODE(right_rheostat1_b[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output535_X (.DIODE(right_rheostat1_b[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output536_X (.DIODE(right_rheostat1_b[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output537_X (.DIODE(right_rheostat2_b[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output538_X (.DIODE(right_rheostat2_b[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output539_X (.DIODE(right_rheostat2_b[2]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output540_X (.DIODE(right_rheostat2_b[3]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output541_X (.DIODE(right_rheostat2_b[4]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output542_X (.DIODE(right_rheostat2_b[5]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output543_X (.DIODE(right_rheostat2_b[6]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output544_X (.DIODE(right_rheostat2_b[7]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output545_X (.DIODE(right_vref_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output546_X (.DIODE(sio0_connect[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output547_X (.DIODE(sio0_connect[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output548_X (.DIODE(sio1_connect[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output549_X (.DIODE(sio1_connect[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output550_X (.DIODE(tempsense_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output551_X (.DIODE(tempsense_sel),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output552_X (.DIODE(tempsense_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output553_X (.DIODE(ulpcomp_clk),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output554_X (.DIODE(ulpcomp_ena),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output555_X (.DIODE(ulpcomp_n_to_analog0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output556_X (.DIODE(ulpcomp_n_to_dac1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output557_X (.DIODE(ulpcomp_n_to_gpio1_6[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output558_X (.DIODE(ulpcomp_n_to_gpio1_6[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output559_X (.DIODE(ulpcomp_n_to_gpio6_1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output560_X (.DIODE(ulpcomp_n_to_gpio6_1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output561_X (.DIODE(ulpcomp_n_to_right_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output562_X (.DIODE(ulpcomp_n_to_sio1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output563_X (.DIODE(ulpcomp_n_to_vbgsc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output564_X (.DIODE(ulpcomp_n_to_vinref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(ulpcomp_out),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output565_X (.DIODE(ulpcomp_p_to_analog1),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output566_X (.DIODE(ulpcomp_p_to_dac0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output567_X (.DIODE(ulpcomp_p_to_gpio1_7[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output568_X (.DIODE(ulpcomp_p_to_gpio1_7[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output569_X (.DIODE(ulpcomp_p_to_gpio6_0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output570_X (.DIODE(ulpcomp_p_to_gpio6_0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output571_X (.DIODE(ulpcomp_p_to_left_vref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output572_X (.DIODE(ulpcomp_p_to_sio0),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output573_X (.DIODE(ulpcomp_p_to_tempsense),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output574_X (.DIODE(ulpcomp_p_to_vbgtc),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output575_X (.DIODE(ulpcomp_p_to_voutref),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output576_X (.DIODE(user_to_adc0[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output577_X (.DIODE(user_to_adc0[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output578_X (.DIODE(user_to_adc1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output579_X (.DIODE(user_to_adc1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output580_X (.DIODE(user_to_comp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output581_X (.DIODE(user_to_comp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output582_X (.DIODE(user_to_comp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output583_X (.DIODE(user_to_comp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output584_X (.DIODE(user_to_ulpcomp_n[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output585_X (.DIODE(user_to_ulpcomp_n[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output586_X (.DIODE(user_to_ulpcomp_p[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output587_X (.DIODE(user_to_ulpcomp_p[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output588_X (.DIODE(vbg_test_to_gpio1_1[0]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output589_X (.DIODE(vbg_test_to_gpio1_1[1]),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output590_X (.DIODE(vbgsc_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output591_X (.DIODE(vbgtc_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(vccd1_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(vccd2_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(vdda1_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(vdda2_pwr_good),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output592_X (.DIODE(vinref_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output593_X (.DIODE(voutref_to_user),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1090_A (.DIODE(n1010),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1085_A (.DIODE(n1010),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1079_Y (.DIODE(n1010),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(n1012),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1161_B1 (.DIODE(n1012),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1155_B1 (.DIODE(n1012),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1146_B1 (.DIODE(n1012),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1094_Y (.DIODE(n1012),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1860_A (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1465_A1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1439_A1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1411_A1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1403_A2 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1348_A1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1320_B1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1281_A1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1263_B1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1257_B1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1213_B2 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1193_A1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1133_A1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1109_B1 (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1108_Y (.DIODE(n1019),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(n1022),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1369_A1 (.DIODE(n1022),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1224_B1 (.DIODE(n1022),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1292_A1 (.DIODE(n1022),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1123_Y (.DIODE(n1022),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1126_D (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1125_X (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1132_Y (.DIODE(n1035),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1055_C (.DIODE(n1035),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1130_X (.DIODE(n1037),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1055_A_N (.DIODE(n1037),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1142_A (.DIODE(n1044),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1055_Y (.DIODE(n1044),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1145_A (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1143_X (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1153_C (.DIODE(n1051),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1097_X (.DIODE(n1051),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1153_A (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1146_X (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1159_B (.DIODE(n1057),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1155_X (.DIODE(n1057),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1165_B (.DIODE(n1062),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1161_X (.DIODE(n1062),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1172_B (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1168_X (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1178_B (.DIODE(n1072),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1174_X (.DIODE(n1072),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1486_A (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1456_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1430_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1390_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1368_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1335_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1315_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1294_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1278_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1246_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1226_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1181_A1 (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1180_Y (.DIODE(n1074),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1913_A (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1466_A1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1440_A1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1434_A2 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1412_A1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1348_B1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1322_A1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1282_A1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1264_B1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1259_A1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1214_A1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1193_B1 (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1192_Y (.DIODE(n1078),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1203_A (.DIODE(n1084),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1199_X (.DIODE(n1084),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1205_D (.DIODE(n1089),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1204_X (.DIODE(n1089),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1205_B (.DIODE(n1091),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1181_X (.DIODE(n1091),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1214_Y (.DIODE(n1094),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1058_D (.DIODE(n1094),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1222_B (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1218_X (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1227_D (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1226_X (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1227_A (.DIODE(n1109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1223_X (.DIODE(n1109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1241_B (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1238_X (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1057_C (.DIODE(n1135),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1045_X (.DIODE(n1135),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1260_A (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1234_X (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1374_B1 (.DIODE(n1142),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1268_X (.DIODE(n1142),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1275_A (.DIODE(n1153),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1271_X (.DIODE(n1153),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1289_C (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1287_X (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1289_B (.DIODE(n1167),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1286_X (.DIODE(n1167),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1301_C (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1295_X (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1312_C (.DIODE(n1189),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1310_X (.DIODE(n1189),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1315_X (.DIODE(n1193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1043_C (.DIODE(n1193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1320_X (.DIODE(n1201),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1066_A (.DIODE(n1201),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1324_A (.DIODE(n1205),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1043_X (.DIODE(n1205),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1325_A (.DIODE(n1208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1307_X (.DIODE(n1208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1329_X (.DIODE(n1209),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1067_D (.DIODE(n1209),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1327_X (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1067_B (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1447_B1 (.DIODE(n1224),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1345_X (.DIODE(n1224),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone18_A (.DIODE(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer1_A (.DIODE(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap618_A (.DIODE(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1244_B (.DIODE(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1113_Y (.DIODE(n1231),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1353_X (.DIODE(n1232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1053_D (.DIODE(n1232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1356_X (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1064_C (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1362_X (.DIODE(n1247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1068_C (.DIODE(n1247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1364_X (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1035_A (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1372_C1 (.DIODE(n1254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1371_X (.DIODE(n1254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1380_A (.DIODE(n1263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1378_X (.DIODE(n1263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1384_X (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1037_B (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_B (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1198_B (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_B (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1112_B (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_B (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1211_B (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1340_A (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1267_A (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1220_A (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1121_A (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1111_Y (.DIODE(n1287),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1420_D (.DIODE(n1312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1417_X (.DIODE(n1312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1421_C (.DIODE(n1316),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1052_X (.DIODE(n1316),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1426_X (.DIODE(n1323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1032_D (.DIODE(n1323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1423_X (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1032_A (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1438_B1 (.DIODE(n1332),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1436_X (.DIODE(n1332),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1431_X (.DIODE(n1337),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1395_A (.DIODE(n1337),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1444_X (.DIODE(n1344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1041_B (.DIODE(n1344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1347_B (.DIODE(n1347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1042_X (.DIODE(n1347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1452_X (.DIODE(n1352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1033_D (.DIODE(n1352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1449_X (.DIODE(n1355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1033_A (.DIODE(n1355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1462_X (.DIODE(n1362),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1437_B1 (.DIODE(n1362),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1457_X (.DIODE(n1367),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1394_A (.DIODE(n1367),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1470_X (.DIODE(n1374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1065_B (.DIODE(n1374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1346_B (.DIODE(n1377),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1054_X (.DIODE(n1377),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1497_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1496_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1495_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1494_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1493_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1492_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1491_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1490_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1489_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1488_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1487_S (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1486_Y (.DIODE(n1388),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1528_A (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1456_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1430_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1391_A1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1369_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1336_A1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1315_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1293_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1277_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1247_A1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1225_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1179_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1140_A1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1122_B1 (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1121_Y (.DIODE(n1393),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1599_A (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1469_B1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1443_B1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1417_A1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1361_A1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1355_A1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1304_A1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1283_B1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1268_A1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1228_B1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1217_A1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1191_A1 (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1190_Y (.DIODE(n1397),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(n1399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1164_A2 (.DIODE(n1399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1158_A2 (.DIODE(n1399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1436_A1 (.DIODE(n1399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1103_Y (.DIODE(n1399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1630_A (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1451_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1425_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1385_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1365_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1327_B1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1309_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1288_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1272_B1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1239_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1219_B1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1202_A1 (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1200_Y (.DIODE(n1401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_A (.DIODE(n1403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1377_B2 (.DIODE(n1403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1154_B1 (.DIODE(n1403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1160_B1 (.DIODE(n1403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1116_Y (.DIODE(n1403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1366_B1 (.DIODE(n1405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1328_A1 (.DIODE(n1405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1310_A1 (.DIODE(n1405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1290_A1 (.DIODE(n1405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1273_B1 (.DIODE(n1405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1202_B1 (.DIODE(n1405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1201_Y (.DIODE(n1405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1461_B1 (.DIODE(n1407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1435_B1 (.DIODE(n1407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1344_B1 (.DIODE(n1407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1254_A1 (.DIODE(n1407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1253_Y (.DIODE(n1407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1049_B (.DIODE(n1407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone14_A (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1442_B1 (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1468_B1 (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1115_B1 (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1131_B1 (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1157_B1 (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1163_B1 (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1114_Y (.DIODE(n1408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout597_A (.DIODE(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1700_S (.DIODE(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1696_S (.DIODE(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1682_S (.DIODE(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1681_S (.DIODE(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1680_S (.DIODE(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1679_Y (.DIODE(n1409),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1701_A (.DIODE(n1410),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1466_B1 (.DIODE(n1410),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1440_B1 (.DIODE(n1410),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1414_A1 (.DIODE(n1410),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1351_B1 (.DIODE(n1410),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1350_Y (.DIODE(n1410),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1706_A (.DIODE(n1412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1467_B1 (.DIODE(n1412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1441_B1 (.DIODE(n1412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1416_B1 (.DIODE(n1412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1353_B1 (.DIODE(n1412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1352_Y (.DIODE(n1412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1711_A (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1449_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1423_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1383_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1365_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1357_A1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1308_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1287_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1271_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1236_B1 (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1235_Y (.DIODE(n1414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1720_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1719_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1718_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1717_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1716_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1715_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1714_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1713_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1712_S (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1711_Y (.DIODE(n1415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1731_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1730_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1729_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1728_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1727_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1726_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1725_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1724_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1723_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1722_S (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1721_Y (.DIODE(n1417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1732_A (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1459_A1 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1433_A1 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1408_A1_N (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1402_A2 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1342_A1 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1319_A2 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1298_B1 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1261_A1 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1254_B1 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1209_A2 (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1207_Y (.DIODE(n1418),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1742_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1741_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1740_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1739_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1738_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1737_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1736_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1735_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1734_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1733_S (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1732_Y (.DIODE(n1419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1471_B1 (.DIODE(n1420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1445_B1 (.DIODE(n1420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1418_B1 (.DIODE(n1420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1356_B1 (.DIODE(n1420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1268_B1 (.DIODE(n1420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1199_B1 (.DIODE(n1420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1198_Y (.DIODE(n1420),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1754_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1753_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1752_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1751_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1750_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1749_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1748_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1747_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1746_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1745_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1744_S (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1743_Y (.DIODE(n1421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1468_A1 (.DIODE(n1422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1413_B1 (.DIODE(n1422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1376_B1 (.DIODE(n1422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1375_A2 (.DIODE(n1422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1351_A1 (.DIODE(n1422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1323_A1 (.DIODE(n1422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1211_Y (.DIODE(n1422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1765_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1764_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1763_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1762_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1761_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1760_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1759_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1758_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1757_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1756_S (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1755_Y (.DIODE(n1423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1766_A (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1462_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1436_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1411_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1400_A2 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1345_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1299_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1266_B2 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1261_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1256_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1208_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1184_B1 (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1183_Y (.DIODE(n1424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1777_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1776_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1775_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1774_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1773_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1772_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1771_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1770_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1769_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1768_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1767_S (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1766_Y (.DIODE(n1425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1778_A (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1450_A1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1424_A1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1384_B1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1366_A1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1326_B1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1309_B1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1288_B1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1238_B1 (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1237_Y (.DIODE(n1426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1419_B1 (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1787_A (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1472_B1 (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1446_B1 (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1364_B1 (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1357_B1 (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1306_B1 (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1233_B1 (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1232_Y (.DIODE(n1428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1795_A (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1471_A1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1445_A1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1418_A1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1362_B1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1355_B1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1305_A1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1284_B1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1230_B1 (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1229_Y (.DIODE(n1430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1803_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1802_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1801_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1800_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1799_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1798_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1797_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1796_S (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1795_Y (.DIODE(n1431),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1804_A (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1453_B1 (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1427_B1 (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1387_A1 (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1378_A1 (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1329_B1 (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1311_B1 (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1245_B1 (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1244_Y (.DIODE(n1432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1811_S (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1810_S (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1809_S (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1808_S (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1807_S (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1806_S (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1805_S (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1804_Y (.DIODE(n1433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1812_A (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1452_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1426_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1387_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1378_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1330_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1313_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1292_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1274_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1240_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1223_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1187_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1130_B1 (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1129_Y (.DIODE(n1434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1824_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1823_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1822_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1821_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1820_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1819_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1818_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1817_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1816_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1815_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1814_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1813_S (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1812_Y (.DIODE(n1435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1825_A (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1454_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1428_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1388_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1379_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1330_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1314_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1291_B1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1277_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1242_B1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1225_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1187_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1138_A1 (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1137_Y (.DIODE(n1436),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1838_A (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1452_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1426_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1386_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1367_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1329_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1311_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1291_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1276_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1242_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1224_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1189_A1 (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1188_Y (.DIODE(n1438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1849_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1848_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1847_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1846_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1845_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1844_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1843_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1842_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1841_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1840_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1839_S (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1838_Y (.DIODE(n1439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1850_A (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1458_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1432_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1391_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1368_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1336_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1316_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1294_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1278_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1249_B1 (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1248_Y (.DIODE(n1440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1859_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1858_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1857_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1856_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1855_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1854_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1853_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1852_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1851_S (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1850_Y (.DIODE(n1441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1873_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1872_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1871_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1870_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1869_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1868_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1867_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1866_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1865_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1864_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1863_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1862_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1861_S (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1860_Y (.DIODE(n1442),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1874_A (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1450_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1424_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1386_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1367_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1328_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1310_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1290_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1274_A1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1239_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1223_A1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1189_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1135_B1 (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1134_Y (.DIODE(n1443),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1886_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1885_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1884_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1883_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1882_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1881_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1880_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1879_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1878_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1877_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1876_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1875_S (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1874_Y (.DIODE(n1444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1887_A (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1470_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1444_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1419_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1362_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1356_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1304_B1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1285_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1271_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1231_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1218_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1191_B1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1130_A1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1119_B1 (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1118_Y (.DIODE(n1445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1900_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1899_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1898_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1897_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1896_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1895_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1894_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1893_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1892_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1891_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1890_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1889_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1888_S (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1887_Y (.DIODE(n1446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1901_A (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1465_B1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1439_B1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1434_B2 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1412_B1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1377_A2 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1349_A1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1321_B1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1299_A1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1258_A1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1214_B1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1196_A1 (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1195_Y (.DIODE(n1447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1912_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1911_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1910_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1909_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1908_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1907_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1906_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1905_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1904_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1903_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1902_S (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1901_Y (.DIODE(n1448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1925_A (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1449_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1423_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1384_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1364_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1327_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1308_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1287_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1273_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1238_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1221_A1 (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1220_Y (.DIODE(n1450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1467_A1 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1441_A1 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1413_A1 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1376_A1 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1375_B2 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1349_B1 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1322_B1 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1258_B1 (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1112_Y (.DIODE(n1452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1950_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1949_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1948_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1947_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1946_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1945_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1944_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1943_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1942_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1941_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1940_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1939_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1938_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1937_S (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1936_Y (.DIODE(n1453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(n1455),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1306_A1 (.DIODE(n1455),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1970_A (.DIODE(n1455),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1272_A1 (.DIODE(n1455),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1120_Y (.DIODE(n1455),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(n1457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1990_S (.DIODE(n1457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1991_S (.DIODE(n1457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1989_Y (.DIODE(n1457),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2008_A (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1453_A1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1427_A1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1389_A1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1379_B1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1332_B1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1313_A1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1293_A1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1245_A1 (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1243_Y (.DIODE(n1458),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2016_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2015_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2014_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2013_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2012_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2011_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2010_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2009_S (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2008_Y (.DIODE(n1459),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2021_S (.DIODE(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2020_S (.DIODE(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2019_S (.DIODE(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2018_S (.DIODE(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2017_Y (.DIODE(n1461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_A (.DIODE(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_A (.DIODE(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1525_A (.DIODE(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1701_B (.DIODE(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1485_X (.DIODE(n1462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2022_A (.DIODE(n1463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1455_A1 (.DIODE(n1463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1429_A1 (.DIODE(n1463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1388_B1 (.DIODE(n1463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1332_A1 (.DIODE(n1463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1331_Y (.DIODE(n1463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_A (.DIODE(n1466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1458_A1 (.DIODE(n1466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1069_X (.DIODE(n1466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2035_A1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2034_A1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2033_A1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1542_A (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1206_B1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1175_B1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1169_B1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1166_A (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1162_B1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1156_B1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1148_B2 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1144_B1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1101_B1 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1100_Y (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1096_B2 (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1069_A (.DIODE(n1469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1434_X (.DIODE(n1485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1400_B1 (.DIODE(n1485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload1_A (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_3__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_1__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_0__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_1__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_15__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_17__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_0__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_11__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_PCLK_X (.DIODE(clknet_leaf_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_X (.DIODE(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1404_A1 (.DIODE(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1152_B (.DIODE(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1113_C (.DIODE(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1106_A (.DIODE(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1099_B (.DIODE(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1091_A (.DIODE(net9),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1080_B (.DIODE(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_X (.DIODE(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1136_B (.DIODE(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1117_B (.DIODE(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1111_B (.DIODE(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1104_A (.DIODE(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1089_C (.DIODE(net10),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_X (.DIODE(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1111_C (.DIODE(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1095_B (.DIODE(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1081_A (.DIODE(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1050_B (.DIODE(net11),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1080_A (.DIODE(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_X (.DIODE(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1124_C (.DIODE(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1117_C (.DIODE(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1088_A (.DIODE(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1050_A (.DIODE(net12),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_X (.DIODE(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1252_A_N (.DIODE(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1128_B (.DIODE(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1113_B (.DIODE(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1106_B (.DIODE(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1092_A (.DIODE(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1083_A (.DIODE(net13),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1063_B (.DIODE(net14),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_X (.DIODE(net14),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1252_B (.DIODE(net14),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1083_B (.DIODE(net14),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout703_A (.DIODE(net18),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout682_A (.DIODE(net18),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_X (.DIODE(net18),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire663_A (.DIODE(net20),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout660_A (.DIODE(net20),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net20),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout659_A (.DIODE(net21),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout658_A (.DIODE(net21),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_X (.DIODE(net21),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_X (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1994_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1975_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1956_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1937_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1889_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1862_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1687_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1645_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1614_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1593_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1559_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1529_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1523_A0 (.DIODE(net23),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_X (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1995_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1976_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1957_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1938_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1688_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1646_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1615_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1594_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1560_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1511_A0 (.DIODE(net24),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire656_A (.DIODE(net25),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_X (.DIODE(net25),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire655_A (.DIODE(net26),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net26),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire654_A (.DIODE(net27),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net27),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire653_A (.DIODE(net28),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_X (.DIODE(net28),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_X (.DIODE(net29),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1682_A0 (.DIODE(net29),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1580_A0 (.DIODE(net29),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1565_A0 (.DIODE(net29),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1503_A0 (.DIODE(net29),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_X (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1681_A0 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1579_A0 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1566_A0 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1504_A0 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire652_A (.DIODE(net31),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout649_A (.DIODE(net31),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_X (.DIODE(net31),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_X (.DIODE(net32),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1680_A0 (.DIODE(net32),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1575_A0 (.DIODE(net32),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1567_A0 (.DIODE(net32),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1505_A0 (.DIODE(net32),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_X (.DIODE(net33),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1576_A0 (.DIODE(net33),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1568_A0 (.DIODE(net33),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1506_A0 (.DIODE(net33),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_X (.DIODE(net34),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1577_A0 (.DIODE(net34),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1569_A0 (.DIODE(net34),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1507_A0 (.DIODE(net34),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_X (.DIODE(net35),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1578_A0 (.DIODE(net35),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1570_A0 (.DIODE(net35),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1508_A0 (.DIODE(net35),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_X (.DIODE(net36),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1574_A0 (.DIODE(net36),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1571_A0 (.DIODE(net36),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1509_A0 (.DIODE(net36),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout647_A (.DIODE(net42),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_X (.DIODE(net42),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout643_A (.DIODE(net43),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_X (.DIODE(net43),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire640_A (.DIODE(net44),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout638_A (.DIODE(net44),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_X (.DIODE(net44),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire637_A (.DIODE(net45),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout635_A (.DIODE(net45),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_X (.DIODE(net45),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire634_A (.DIODE(net46),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout633_A (.DIODE(net46),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_X (.DIODE(net46),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_X (.DIODE(net50),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1485_B (.DIODE(net50),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output63_A (.DIODE(net63),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1205_X (.DIODE(net63),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output64_A (.DIODE(net64),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1142_X (.DIODE(net64),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output65_A (.DIODE(net65),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1127_X (.DIODE(net65),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output67_A (.DIODE(net67),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1178_X (.DIODE(net67),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output68_A (.DIODE(net68),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1165_X (.DIODE(net68),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output69_A (.DIODE(net69),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1159_X (.DIODE(net69),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output70_A (.DIODE(net70),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1172_X (.DIODE(net70),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output71_A (.DIODE(net71),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1477_X (.DIODE(net71),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1480_X (.DIODE(net72),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1359_X (.DIODE(net73),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1474_X (.DIODE(net84),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout619_A (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1478_B1 (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1475_B1 (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1459_B1 (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1433_B1 (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1370_B1 (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1319_B1 (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1071_Y (.DIODE(net85),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1448_X (.DIODE(net87),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1260_X (.DIODE(net88),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1325_X (.DIODE(net89),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1382_X (.DIODE(net90),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1302_X (.DIODE(net91),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1070_X (.DIODE(net92),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1056_X (.DIODE(net93),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1417_B1 (.DIODE(net95),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_0__Q (.DIODE(net95),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1731_A1 (.DIODE(net95),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_8__Q (.DIODE(net96),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1722_A1 (.DIODE(net96),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1374_A1 (.DIODE(net96),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_9__Q (.DIODE(net97),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1723_A1 (.DIODE(net97),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1217_B2 (.DIODE(net97),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_6__Q (.DIODE(net98),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1724_A1 (.DIODE(net98),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1361_B2 (.DIODE(net98),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_7__Q (.DIODE(net99),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1725_A1 (.DIODE(net99),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1285_B2 (.DIODE(net99),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_1__Q (.DIODE(net104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1719_A1 (.DIODE(net104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1357_A2 (.DIODE(net104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_7__Q (.DIODE(net106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1712_A1 (.DIODE(net106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1287_B2 (.DIODE(net106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output107_A (.DIODE(net107),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_8__Q (.DIODE(net107),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1713_A1 (.DIODE(net107),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1271_B2 (.DIODE(net107),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output108_A (.DIODE(net108),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_5__Q (.DIODE(net108),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1714_A1 (.DIODE(net108),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1308_B2 (.DIODE(net108),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_6__Q (.DIODE(net109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1715_A1 (.DIODE(net109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1365_B2 (.DIODE(net109),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_4__Q (.DIODE(net112),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1716_A1 (.DIODE(net112),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1236_B2 (.DIODE(net112),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_0__Q (.DIODE(net113),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2015_A1 (.DIODE(net113),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1389_A2 (.DIODE(net113),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_1__Q (.DIODE(net114),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2016_A1 (.DIODE(net114),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1332_B2 (.DIODE(net114),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_4__Q (.DIODE(net115),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2011_A1 (.DIODE(net115),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1245_A2 (.DIODE(net115),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output116_A (.DIODE(net116),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_5__Q (.DIODE(net116),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2012_A1 (.DIODE(net116),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1313_A2 (.DIODE(net116),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output117_A (.DIODE(net117),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_ana_REG_reg_0__Q (.DIODE(net117),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1704_A1 (.DIODE(net117),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1414_A2 (.DIODE(net117),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output119_A (.DIODE(net119),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_ana_REG_reg_2__Q (.DIODE(net119),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1702_A1 (.DIODE(net119),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1466_B2 (.DIODE(net119),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_ana_REG_reg_3__Q (.DIODE(net120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1703_A1 (.DIODE(net120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1440_B2 (.DIODE(net120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_2__Q (.DIODE(net121),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1675_A1 (.DIODE(net121),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1461_B2 (.DIODE(net121),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output122_A (.DIODE(net122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_3__Q (.DIODE(net122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1676_A1 (.DIODE(net122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1435_B2 (.DIODE(net122),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output124_A (.DIODE(net124),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_5__Q (.DIODE(net124),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1674_A1 (.DIODE(net124),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1266_A1 (.DIODE(net124),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output132_A (.DIODE(net132),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_15__Q (.DIODE(net132),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1596_A1 (.DIODE(net132),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1163_A2 (.DIODE(net132),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output133_A (.DIODE(net133),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_16__Q (.DIODE(net133),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1597_A1 (.DIODE(net133),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1157_A2 (.DIODE(net133),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_4__Q (.DIODE(net136),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1585_A1 (.DIODE(net136),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1256_A2 (.DIODE(net136),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output140_A (.DIODE(net140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_8__Q (.DIODE(net140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1589_A1 (.DIODE(net140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1263_A2 (.DIODE(net140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output141_A (.DIODE(net141),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_9__Q (.DIODE(net141),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1590_A1 (.DIODE(net141),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1208_A2 (.DIODE(net141),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output144_A (.DIODE(net144),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_7__Q (.DIODE(net144),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1490_A1 (.DIODE(net144),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1294_A2 (.DIODE(net144),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output145_A (.DIODE(net145),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_8__Q (.DIODE(net145),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1489_A1 (.DIODE(net145),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1278_A2 (.DIODE(net145),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output148_A (.DIODE(net148),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_6__Q (.DIODE(net148),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1493_A1 (.DIODE(net148),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1368_A2 (.DIODE(net148),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output149_A (.DIODE(net149),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_10__Q (.DIODE(net149),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1487_A1 (.DIODE(net149),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1181_A2 (.DIODE(net149),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_1__Q (.DIODE(net157),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1741_A1 (.DIODE(net157),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1342_A2 (.DIODE(net157),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output158_A (.DIODE(net158),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_0__Q (.DIODE(net158),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1742_A1 (.DIODE(net158),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1408_A2_N (.DIODE(net158),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output159_A (.DIODE(net159),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_8__Q (.DIODE(net159),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1733_A1 (.DIODE(net159),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1261_A2 (.DIODE(net159),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output160_A (.DIODE(net160),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_9__Q (.DIODE(net160),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1734_A1 (.DIODE(net160),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1209_A1 (.DIODE(net160),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_6__Q (.DIODE(net161),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1735_A1 (.DIODE(net161),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1402_A1 (.DIODE(net161),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output162_A (.DIODE(net162),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_7__Q (.DIODE(net162),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1736_A1 (.DIODE(net162),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1298_B2 (.DIODE(net162),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output163_A (.DIODE(net163),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_4__Q (.DIODE(net163),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1738_A1 (.DIODE(net163),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1254_B2 (.DIODE(net163),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output164_A (.DIODE(net164),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_2__Q (.DIODE(net164),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1740_A1 (.DIODE(net164),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1459_A2 (.DIODE(net164),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output165_A (.DIODE(net165),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_3__Q (.DIODE(net165),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1739_A1 (.DIODE(net165),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1433_A2 (.DIODE(net165),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output166_A (.DIODE(net166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_5__Q (.DIODE(net166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1737_A1 (.DIODE(net166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1319_A1 (.DIODE(net166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_9__Q (.DIODE(net169),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1744_A1 (.DIODE(net169),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1218_B2 (.DIODE(net169),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output170_A (.DIODE(net170),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_10__Q (.DIODE(net170),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1745_A1 (.DIODE(net170),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1199_B2 (.DIODE(net170),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output171_A (.DIODE(net171),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_7__Q (.DIODE(net171),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1746_A1 (.DIODE(net171),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1286_B2 (.DIODE(net171),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output172_A (.DIODE(net172),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_8__Q (.DIODE(net172),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1747_A1 (.DIODE(net172),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1268_B2 (.DIODE(net172),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output174_A (.DIODE(net174),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_2__Q (.DIODE(net174),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1752_A1 (.DIODE(net174),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1471_B2 (.DIODE(net174),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output176_A (.DIODE(net176),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_3__Q (.DIODE(net176),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1751_A1 (.DIODE(net176),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1445_B2 (.DIODE(net176),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_6__Q (.DIODE(net177),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1748_A1 (.DIODE(net177),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1363_B2 (.DIODE(net177),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_4__Q (.DIODE(net181),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1607_A1 (.DIODE(net181),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1228_B2 (.DIODE(net181),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_5__Q (.DIODE(net182),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1608_A1 (.DIODE(net182),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1304_A2 (.DIODE(net182),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_14__Q (.DIODE(net185),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1686_A1 (.DIODE(net185),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1173_B2 (.DIODE(net185),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_1__Q (.DIODE(net186),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1677_A1 (.DIODE(net186),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1344_B2 (.DIODE(net186),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_A (.DIODE(net188),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_2__Q (.DIODE(net188),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2013_A1 (.DIODE(net188),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1453_A2 (.DIODE(net188),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_3__Q (.DIODE(net189),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2014_A1 (.DIODE(net189),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1427_A2 (.DIODE(net189),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_6__Q (.DIODE(net190),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2009_A1 (.DIODE(net190),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1379_B2 (.DIODE(net190),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_7__Q (.DIODE(net191),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2010_A1 (.DIODE(net191),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1293_A2 (.DIODE(net191),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_0__Q (.DIODE(net192),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1572_A1 (.DIODE(net192),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1406_A2 (.DIODE(net192),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_29__Q (.DIODE(net193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1543_A1 (.DIODE(net193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1166_B (.DIODE(net193),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_25__Q (.DIODE(net194),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1544_A1 (.DIODE(net194),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1096_B1 (.DIODE(net194),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output195_A (.DIODE(net195),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_26__Q (.DIODE(net195),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2033_A2 (.DIODE(net195),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1545_A1 (.DIODE(net195),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_27__Q (.DIODE(net196),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2034_A2 (.DIODE(net196),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1546_A1 (.DIODE(net196),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output197_A (.DIODE(net197),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_28__Q (.DIODE(net197),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2035_A2 (.DIODE(net197),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1547_A1 (.DIODE(net197),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output208_A (.DIODE(net208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_20__Q (.DIODE(net208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1567_A1 (.DIODE(net208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1144_B2 (.DIODE(net208),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_21__Q (.DIODE(net210),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1568_A1 (.DIODE(net210),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1481_A2 (.DIODE(net210),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output211_A (.DIODE(net211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_22__Q (.DIODE(net211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2027_A2 (.DIODE(net211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1569_A1 (.DIODE(net211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output212_A (.DIODE(net212),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_23__Q (.DIODE(net212),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1570_A1 (.DIODE(net212),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1483_A2 (.DIODE(net212),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output213_A (.DIODE(net213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_24__Q (.DIODE(net213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2029_A2 (.DIODE(net213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1571_A1 (.DIODE(net213),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output215_A (.DIODE(net215),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_4__Q (.DIODE(net215),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1551_A1 (.DIODE(net215),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1249_A2 (.DIODE(net215),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output222_A (.DIODE(net222),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_0__Q (.DIODE(net222),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2025_A1 (.DIODE(net222),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1388_B2 (.DIODE(net222),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output223_A (.DIODE(net223),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_1__Q (.DIODE(net223),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2026_A1 (.DIODE(net223),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1332_A2 (.DIODE(net223),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output225_A (.DIODE(net225),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_2__Q (.DIODE(net225),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2018_A1 (.DIODE(net225),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1454_B2 (.DIODE(net225),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output226_A (.DIODE(net226),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_3__Q (.DIODE(net226),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2019_A1 (.DIODE(net226),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1428_B2 (.DIODE(net226),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output227_A (.DIODE(net227),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_0__Q (.DIODE(net227),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2020_A1 (.DIODE(net227),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1389_B2 (.DIODE(net227),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output228_A (.DIODE(net228),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_1__Q (.DIODE(net228),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2021_A1 (.DIODE(net228),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1334_A2 (.DIODE(net228),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output229_A (.DIODE(net229),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_0__Q (.DIODE(net229),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1530_A1 (.DIODE(net229),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1391_A2 (.DIODE(net229),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output232_A (.DIODE(net232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_1__Q (.DIODE(net232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1531_A1 (.DIODE(net232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1336_A2 (.DIODE(net232),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output233_A (.DIODE(net233),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_2__Q (.DIODE(net233),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1532_A1 (.DIODE(net233),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1456_B2 (.DIODE(net233),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output234_A (.DIODE(net234),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_3__Q (.DIODE(net234),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1533_A1 (.DIODE(net234),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1430_B2 (.DIODE(net234),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output235_A (.DIODE(net235),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_4__Q (.DIODE(net235),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1534_A1 (.DIODE(net235),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1247_A2 (.DIODE(net235),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output236_A (.DIODE(net236),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_5__Q (.DIODE(net236),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1535_A1 (.DIODE(net236),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1315_B2 (.DIODE(net236),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output242_A (.DIODE(net242),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_24__Q (.DIODE(net242),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2029_B2 (.DIODE(net242),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1574_A1 (.DIODE(net242),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output243_A (.DIODE(net243),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_0__Q (.DIODE(net243),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1660_A1 (.DIODE(net243),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1416_A2 (.DIODE(net243),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output244_A (.DIODE(net244),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_4__Q (.DIODE(net244),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1869_A1 (.DIODE(net244),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1257_B2 (.DIODE(net244),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output245_A (.DIODE(net245),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_3__Q (.DIODE(net245),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1870_A1 (.DIODE(net245),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1439_A2 (.DIODE(net245),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output246_A (.DIODE(net246),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_2__Q (.DIODE(net246),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1871_A1 (.DIODE(net246),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1465_A2 (.DIODE(net246),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output247_A (.DIODE(net247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_11__Q (.DIODE(net247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1861_A1 (.DIODE(net247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1133_A2 (.DIODE(net247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output248_A (.DIODE(net248),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_12__Q (.DIODE(net248),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1862_A1 (.DIODE(net248),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1109_B2 (.DIODE(net248),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output249_A (.DIODE(net249),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_0__Q (.DIODE(net249),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1872_A1 (.DIODE(net249),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1411_A2 (.DIODE(net249),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output250_A (.DIODE(net250),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_1__Q (.DIODE(net250),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1873_A1 (.DIODE(net250),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1348_A2 (.DIODE(net250),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output251_A (.DIODE(net251),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_5__Q (.DIODE(net251),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1868_A1 (.DIODE(net251),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1320_B2 (.DIODE(net251),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output252_A (.DIODE(net252),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_6__Q (.DIODE(net252),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1867_A1 (.DIODE(net252),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1403_A1 (.DIODE(net252),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output253_A (.DIODE(net253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_9__Q (.DIODE(net253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1864_A1 (.DIODE(net253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1213_B1 (.DIODE(net253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output254_A (.DIODE(net254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_7__Q (.DIODE(net254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1866_A1 (.DIODE(net254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1281_A2 (.DIODE(net254),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output255_A (.DIODE(net255),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_8__Q (.DIODE(net255),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1865_A1 (.DIODE(net255),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1263_B2 (.DIODE(net255),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output257_A (.DIODE(net257),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_4__Q (.DIODE(net257),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1882_A1 (.DIODE(net257),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1239_B2 (.DIODE(net257),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_A (.DIODE(net258),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_3__Q (.DIODE(net258),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1883_A1 (.DIODE(net258),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1424_B2 (.DIODE(net258),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output259_A (.DIODE(net259),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_2__Q (.DIODE(net259),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1884_A1 (.DIODE(net259),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1450_B2 (.DIODE(net259),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_A (.DIODE(net260),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_10__Q (.DIODE(net260),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1875_A1 (.DIODE(net260),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1189_B2 (.DIODE(net260),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output261_A (.DIODE(net261),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_11__Q (.DIODE(net261),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1876_A1 (.DIODE(net261),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1135_B2 (.DIODE(net261),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_A (.DIODE(net263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_1__Q (.DIODE(net263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1886_A1 (.DIODE(net263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1328_B2 (.DIODE(net263),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output265_A (.DIODE(net265),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_5__Q (.DIODE(net265),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1881_A1 (.DIODE(net265),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1310_B2 (.DIODE(net265),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output266_A (.DIODE(net266),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_6__Q (.DIODE(net266),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1880_A1 (.DIODE(net266),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1367_B2 (.DIODE(net266),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output267_A (.DIODE(net267),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_7__Q (.DIODE(net267),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1879_A1 (.DIODE(net267),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1290_B2 (.DIODE(net267),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output272_A (.DIODE(net272),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_13__Q (.DIODE(net272),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1957_A1 (.DIODE(net272),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1147_A2 (.DIODE(net272),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output273_A (.DIODE(net273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_10__Q (.DIODE(net273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1958_A1 (.DIODE(net273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1179_A2 (.DIODE(net273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output274_A (.DIODE(net274),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_11__Q (.DIODE(net274),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1959_A1 (.DIODE(net274),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1135_A2 (.DIODE(net274),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_A (.DIODE(net275),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_2__Q (.DIODE(net275),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1966_A1 (.DIODE(net275),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1455_B2 (.DIODE(net275),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output276_A (.DIODE(net276),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_3__Q (.DIODE(net276),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1967_A1 (.DIODE(net276),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1429_B2 (.DIODE(net276),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output281_A (.DIODE(net281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_8__Q (.DIODE(net281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1960_A1 (.DIODE(net281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1276_B2 (.DIODE(net281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output282_A (.DIODE(net282),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_9__Q (.DIODE(net282),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1961_A1 (.DIODE(net282),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1224_B2 (.DIODE(net282),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output283_A (.DIODE(net283),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_6__Q (.DIODE(net283),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1962_A1 (.DIODE(net283),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1369_A2 (.DIODE(net283),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output284_A (.DIODE(net284),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_7__Q (.DIODE(net284),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1963_A1 (.DIODE(net284),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1292_A2 (.DIODE(net284),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_6__Q (.DIODE(net292),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1662_A1 (.DIODE(net292),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1366_B2 (.DIODE(net292),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output293_A (.DIODE(net293),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_7__Q (.DIODE(net293),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1663_A1 (.DIODE(net293),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1290_A2 (.DIODE(net293),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_A (.DIODE(net294),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_8__Q (.DIODE(net294),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1664_A1 (.DIODE(net294),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1273_B2 (.DIODE(net294),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_A (.DIODE(net295),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_9__Q (.DIODE(net295),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1665_A1 (.DIODE(net295),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1221_B2 (.DIODE(net295),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_A (.DIODE(net296),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_10__Q (.DIODE(net296),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1666_A1 (.DIODE(net296),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1202_B2 (.DIODE(net296),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net298),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_3__Q (.DIODE(net298),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1808_A1 (.DIODE(net298),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1427_B2 (.DIODE(net298),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_A (.DIODE(net299),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_2__Q (.DIODE(net299),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1809_A1 (.DIODE(net299),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1453_B2 (.DIODE(net299),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output302_A (.DIODE(net302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_5__Q (.DIODE(net302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1806_A1 (.DIODE(net302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1311_B2 (.DIODE(net302),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output303_A (.DIODE(net303),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_4__Q (.DIODE(net303),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1807_A1 (.DIODE(net303),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1245_B2 (.DIODE(net303),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_A (.DIODE(net305),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_3__Q (.DIODE(net305),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1800_A1 (.DIODE(net305),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1445_A2 (.DIODE(net305),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output306_A (.DIODE(net306),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_2__Q (.DIODE(net306),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1801_A1 (.DIODE(net306),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1471_A2 (.DIODE(net306),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_0__Q (.DIODE(net307),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1802_A1 (.DIODE(net307),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1418_A2 (.DIODE(net307),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_A (.DIODE(net308),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_1__Q (.DIODE(net308),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1803_A1 (.DIODE(net308),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1355_B2 (.DIODE(net308),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output312_A (.DIODE(net312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_7__Q (.DIODE(net312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1796_A1 (.DIODE(net312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1284_B2 (.DIODE(net312),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output315_A (.DIODE(net315),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_10__Q (.DIODE(net315),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1826_A1 (.DIODE(net315),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1187_A2 (.DIODE(net315),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output316_A (.DIODE(net316),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_11__Q (.DIODE(net316),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1827_A1 (.DIODE(net316),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1138_A2 (.DIODE(net316),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output317_A (.DIODE(net317),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_8__Q (.DIODE(net317),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1828_A1 (.DIODE(net317),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1277_A2 (.DIODE(net317),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output318_A (.DIODE(net318),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_9__Q (.DIODE(net318),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1829_A1 (.DIODE(net318),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1225_A2 (.DIODE(net318),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output319_A (.DIODE(net319),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_2__Q (.DIODE(net319),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1834_A1 (.DIODE(net319),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1454_A2 (.DIODE(net319),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output320_A (.DIODE(net320),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_3__Q (.DIODE(net320),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1835_A1 (.DIODE(net320),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1428_A2 (.DIODE(net320),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output321_A (.DIODE(net321),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_6__Q (.DIODE(net321),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1830_A1 (.DIODE(net321),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1379_A2 (.DIODE(net321),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output322_A (.DIODE(net322),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_7__Q (.DIODE(net322),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1831_A1 (.DIODE(net322),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1291_B2 (.DIODE(net322),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output323_A (.DIODE(net323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_0__Q (.DIODE(net323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1836_A1 (.DIODE(net323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1388_A2 (.DIODE(net323),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output331_A (.DIODE(net331),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_5__Q (.DIODE(net331),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1844_A1 (.DIODE(net331),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1311_A2 (.DIODE(net331),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output332_A (.DIODE(net332),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_6__Q (.DIODE(net332),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1843_A1 (.DIODE(net332),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1367_A2 (.DIODE(net332),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output333_A (.DIODE(net333),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_9__Q (.DIODE(net333),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1840_A1 (.DIODE(net333),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1224_A2 (.DIODE(net333),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output334_A (.DIODE(net334),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_7__Q (.DIODE(net334),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1842_A1 (.DIODE(net334),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1291_A2 (.DIODE(net334),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output335_A (.DIODE(net335),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_8__Q (.DIODE(net335),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1841_A1 (.DIODE(net335),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1276_A2 (.DIODE(net335),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output338_A (.DIODE(net338),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_3__Q (.DIODE(net338),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1856_A1 (.DIODE(net338),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1432_B2 (.DIODE(net338),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output339_A (.DIODE(net339),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_2__Q (.DIODE(net339),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1857_A1 (.DIODE(net339),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1458_B2 (.DIODE(net339),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output340_A (.DIODE(net340),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_0__Q (.DIODE(net340),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1858_A1 (.DIODE(net340),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1391_B2 (.DIODE(net340),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output341_A (.DIODE(net341),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_1__Q (.DIODE(net341),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1859_A1 (.DIODE(net341),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1336_B2 (.DIODE(net341),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output342_A (.DIODE(net342),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_7__Q (.DIODE(net342),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1852_A1 (.DIODE(net342),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1294_B2 (.DIODE(net342),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output344_A (.DIODE(net344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_6__Q (.DIODE(net344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1853_A1 (.DIODE(net344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1368_B2 (.DIODE(net344),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output345_A (.DIODE(net345),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_8__Q (.DIODE(net345),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1851_A1 (.DIODE(net345),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1278_B2 (.DIODE(net345),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output346_A (.DIODE(net346),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_4__Q (.DIODE(net346),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1945_A1 (.DIODE(net346),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1258_B2 (.DIODE(net346),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output347_A (.DIODE(net347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_5__Q (.DIODE(net347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1946_A1 (.DIODE(net347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1322_B2 (.DIODE(net347),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output348_A (.DIODE(net348),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_10__Q (.DIODE(net348),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1939_A1 (.DIODE(net348),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1196_B2 (.DIODE(net348),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output349_A (.DIODE(net349),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_11__Q (.DIODE(net349),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1940_A1 (.DIODE(net349),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1132_B2 (.DIODE(net349),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output350_A (.DIODE(net350),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_8__Q (.DIODE(net350),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1941_A1 (.DIODE(net350),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1375_B1 (.DIODE(net350),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output351_A (.DIODE(net351),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_9__Q (.DIODE(net351),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1942_A1 (.DIODE(net351),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1212_A2 (.DIODE(net351),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output352_A (.DIODE(net352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_2__Q (.DIODE(net352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1947_A1 (.DIODE(net352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1467_A2 (.DIODE(net352),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output353_A (.DIODE(net353),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_3__Q (.DIODE(net353),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1948_A1 (.DIODE(net353),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1441_A2 (.DIODE(net353),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output354_A (.DIODE(net354),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_12__Q (.DIODE(net354),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1937_A1 (.DIODE(net354),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1115_A2 (.DIODE(net354),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output355_A (.DIODE(net355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_13__Q (.DIODE(net355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1938_A1 (.DIODE(net355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1150_B2 (.DIODE(net355),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output356_A (.DIODE(net356),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_6__Q (.DIODE(net356),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1943_A1 (.DIODE(net356),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1376_A2 (.DIODE(net356),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output357_A (.DIODE(net357),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_7__Q (.DIODE(net357),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1944_A1 (.DIODE(net357),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1281_B2 (.DIODE(net357),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output358_A (.DIODE(net358),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_0__Q (.DIODE(net358),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1949_A1 (.DIODE(net358),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1413_A2 (.DIODE(net358),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output359_A (.DIODE(net359),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_1__Q (.DIODE(net359),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1950_A1 (.DIODE(net359),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1349_B2 (.DIODE(net359),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output362_A (.DIODE(net362),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_4__Q (.DIODE(net362),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1653_A1 (.DIODE(net362),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1230_A2 (.DIODE(net362),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output363_A (.DIODE(net363),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_5__Q (.DIODE(net363),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1654_A1 (.DIODE(net363),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1303_A2 (.DIODE(net363),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output364_A (.DIODE(net364),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_6__Q (.DIODE(net364),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1655_A1 (.DIODE(net364),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1360_A2 (.DIODE(net364),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output365_A (.DIODE(net365),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_7__Q (.DIODE(net365),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1656_A1 (.DIODE(net365),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1284_A2 (.DIODE(net365),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output366_A (.DIODE(net366),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_8__Q (.DIODE(net366),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1657_A1 (.DIODE(net366),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1377_B1 (.DIODE(net366),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output367_A (.DIODE(net367),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_9__Q (.DIODE(net367),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1658_A1 (.DIODE(net367),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1210_A2 (.DIODE(net367),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output368_A (.DIODE(net368),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_10__Q (.DIODE(net368),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1643_A1 (.DIODE(net368),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1194_A2 (.DIODE(net368),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output369_A (.DIODE(net369),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_11__Q (.DIODE(net369),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1644_A1 (.DIODE(net369),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1133_B2 (.DIODE(net369),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output370_A (.DIODE(net370),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_12__Q (.DIODE(net370),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1645_A1 (.DIODE(net370),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1119_A2 (.DIODE(net370),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output371_A (.DIODE(net371),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_13__Q (.DIODE(net371),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1646_A1 (.DIODE(net371),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1151_A2 (.DIODE(net371),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output372_A (.DIODE(net372),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_14__Q (.DIODE(net372),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1647_A1 (.DIODE(net372),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1173_A2 (.DIODE(net372),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output373_A (.DIODE(net373),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_15__Q (.DIODE(net373),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1648_A1 (.DIODE(net373),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1160_B2 (.DIODE(net373),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output374_A (.DIODE(net374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_16__Q (.DIODE(net374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1649_A1 (.DIODE(net374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1154_B2 (.DIODE(net374),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output375_A (.DIODE(net375),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_17__Q (.DIODE(net375),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1650_A1 (.DIODE(net375),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1167_A2 (.DIODE(net375),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output376_A (.DIODE(net376),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_18__Q (.DIODE(net376),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1682_A1 (.DIODE(net376),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1475_A2 (.DIODE(net376),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output379_A (.DIODE(net379),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_21__Q (.DIODE(net379),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1576_A1 (.DIODE(net379),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1481_B2 (.DIODE(net379),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output380_A (.DIODE(net380),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_22__Q (.DIODE(net380),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2027_B2 (.DIODE(net380),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1577_A1 (.DIODE(net380),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output381_A (.DIODE(net381),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_23__Q (.DIODE(net381),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1578_A1 (.DIODE(net381),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1483_B2 (.DIODE(net381),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output384_A (.DIODE(net384),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_11__Q (.DIODE(net384),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1522_A1 (.DIODE(net384),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1140_B2 (.DIODE(net384),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output386_A (.DIODE(net386),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_2__Q (.DIODE(net386),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1513_A1 (.DIODE(net386),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1457_B2 (.DIODE(net386),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output387_A (.DIODE(net387),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_3__Q (.DIODE(net387),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1514_A1 (.DIODE(net387),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1431_B2 (.DIODE(net387),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output389_A (.DIODE(net389),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_5__Q (.DIODE(net389),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1516_A1 (.DIODE(net389),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1317_A2 (.DIODE(net389),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output392_A (.DIODE(net392),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_8__Q (.DIODE(net392),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1519_A1 (.DIODE(net392),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1262_A2 (.DIODE(net392),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output396_A (.DIODE(net396),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_14__Q (.DIODE(net396),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1499_A1 (.DIODE(net396),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1177_A2 (.DIODE(net396),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output398_A (.DIODE(net398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_25__Q (.DIODE(net398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1510_A1 (.DIODE(net398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1096_A1 (.DIODE(net398),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output399_A (.DIODE(net399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_15__Q (.DIODE(net399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1500_A1 (.DIODE(net399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1162_A2 (.DIODE(net399),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output400_A (.DIODE(net400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_16__Q (.DIODE(net400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1501_A1 (.DIODE(net400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1156_A2 (.DIODE(net400),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output401_A (.DIODE(net401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_17__Q (.DIODE(net401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1502_A1 (.DIODE(net401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1171_A2 (.DIODE(net401),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output402_A (.DIODE(net402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_18__Q (.DIODE(net402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1503_A1 (.DIODE(net402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1476_A2 (.DIODE(net402),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output403_A (.DIODE(net403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_19__Q (.DIODE(net403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1504_A1 (.DIODE(net403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1479_A2 (.DIODE(net403),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output405_A (.DIODE(net405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_21__Q (.DIODE(net405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1506_A1 (.DIODE(net405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1482_A2 (.DIODE(net405),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output406_A (.DIODE(net406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_22__Q (.DIODE(net406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2028_A2 (.DIODE(net406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1507_A1 (.DIODE(net406),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output407_A (.DIODE(net407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_23__Q (.DIODE(net407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1508_A1 (.DIODE(net407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1484_A2 (.DIODE(net407),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output408_A (.DIODE(net408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_0__Q (.DIODE(net408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1629_A1 (.DIODE(net408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1409_B2 (.DIODE(net408),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output412_A (.DIODE(net412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_11__Q (.DIODE(net412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1888_A1 (.DIODE(net412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1130_A2 (.DIODE(net412),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output413_A (.DIODE(net413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_12__Q (.DIODE(net413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1889_A1 (.DIODE(net413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1119_B2 (.DIODE(net413),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output414_A (.DIODE(net414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_0__Q (.DIODE(net414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1899_A1 (.DIODE(net414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1419_A2 (.DIODE(net414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output415_A (.DIODE(net415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_1__Q (.DIODE(net415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1900_A1 (.DIODE(net415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1356_A2 (.DIODE(net415),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output416_A (.DIODE(net416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_5__Q (.DIODE(net416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1895_A1 (.DIODE(net416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1304_B2 (.DIODE(net416),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output417_A (.DIODE(net417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_6__Q (.DIODE(net417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1894_A1 (.DIODE(net417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1362_A2 (.DIODE(net417),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output419_A (.DIODE(net419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_7__Q (.DIODE(net419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1893_A1 (.DIODE(net419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1285_A2 (.DIODE(net419),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output421_A (.DIODE(net421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_10__Q (.DIODE(net421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1890_A1 (.DIODE(net421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1191_B2 (.DIODE(net421),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output422_A (.DIODE(net422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_4__Q (.DIODE(net422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1908_A1 (.DIODE(net422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1258_A2 (.DIODE(net422),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output423_A (.DIODE(net423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_3__Q (.DIODE(net423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1909_A1 (.DIODE(net423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1439_B2 (.DIODE(net423),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output424_A (.DIODE(net424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_2__Q (.DIODE(net424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1910_A1 (.DIODE(net424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1465_B2 (.DIODE(net424),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output425_A (.DIODE(net425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_9__Q (.DIODE(net425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1902_A1 (.DIODE(net425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1214_B2 (.DIODE(net425),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output426_A (.DIODE(net426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_10__Q (.DIODE(net426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1903_A1 (.DIODE(net426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1196_A2 (.DIODE(net426),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output427_A (.DIODE(net427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_0__Q (.DIODE(net427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1911_A1 (.DIODE(net427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1412_B2 (.DIODE(net427),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output428_A (.DIODE(net428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_1__Q (.DIODE(net428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1912_A1 (.DIODE(net428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1349_A2 (.DIODE(net428),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output429_A (.DIODE(net429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_7__Q (.DIODE(net429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1905_A1 (.DIODE(net429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1299_A2 (.DIODE(net429),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output430_A (.DIODE(net430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_5__Q (.DIODE(net430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1907_A1 (.DIODE(net430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1321_B2 (.DIODE(net430),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output432_A (.DIODE(net432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_8__Q (.DIODE(net432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1904_A1 (.DIODE(net432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1377_A1 (.DIODE(net432),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output433_A (.DIODE(net433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_4__Q (.DIODE(net433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1983_A1 (.DIODE(net433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1236_A2 (.DIODE(net433),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output434_A (.DIODE(net434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_5__Q (.DIODE(net434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1984_A1 (.DIODE(net434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1306_A2 (.DIODE(net434),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output435_A (.DIODE(net435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_12__Q (.DIODE(net435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1975_A1 (.DIODE(net435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1122_A2 (.DIODE(net435),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output438_A (.DIODE(net438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_11__Q (.DIODE(net438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1978_A1 (.DIODE(net438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1131_A2 (.DIODE(net438),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output439_A (.DIODE(net439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_2__Q (.DIODE(net439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1985_A1 (.DIODE(net439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1472_A2 (.DIODE(net439),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output440_A (.DIODE(net440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_3__Q (.DIODE(net440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1986_A1 (.DIODE(net440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1446_A2 (.DIODE(net440),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output441_A (.DIODE(net441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_16__Q (.DIODE(net441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1971_A1 (.DIODE(net441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1154_A2 (.DIODE(net441),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output444_A (.DIODE(net444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_15__Q (.DIODE(net444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1974_A1 (.DIODE(net444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1160_A2 (.DIODE(net444),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output445_A (.DIODE(net445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_8__Q (.DIODE(net445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1979_A1 (.DIODE(net445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1272_A2 (.DIODE(net445),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output446_A (.DIODE(net446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_9__Q (.DIODE(net446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1980_A1 (.DIODE(net446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1219_A2 (.DIODE(net446),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output447_A (.DIODE(net447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_6__Q (.DIODE(net447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1981_A1 (.DIODE(net447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1363_A2 (.DIODE(net447),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output448_A (.DIODE(net448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_7__Q (.DIODE(net448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1982_A1 (.DIODE(net448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1286_A2 (.DIODE(net448),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output449_A (.DIODE(net449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_0__Q (.DIODE(net449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1987_A1 (.DIODE(net449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1383_A2 (.DIODE(net449),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output450_A (.DIODE(net450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_1__Q (.DIODE(net450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1988_A1 (.DIODE(net450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1326_A2 (.DIODE(net450),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output452_A (.DIODE(net452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_2__Q (.DIODE(net452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1637_A1 (.DIODE(net452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1451_A2 (.DIODE(net452),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output453_A (.DIODE(net453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_3__Q (.DIODE(net453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1638_A1 (.DIODE(net453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1425_A2 (.DIODE(net453),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output454_A (.DIODE(net454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_4__Q (.DIODE(net454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1639_A1 (.DIODE(net454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1239_A2 (.DIODE(net454),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output461_A (.DIODE(net461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_0__Q (.DIODE(net461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1641_A1 (.DIODE(net461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1385_A2 (.DIODE(net461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output462_A (.DIODE(net462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_1__Q (.DIODE(net462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1793_A1 (.DIODE(net462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1357_B2 (.DIODE(net462),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1419_B2 (.DIODE(net463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output463_A (.DIODE(net463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_0__Q (.DIODE(net463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1794_A1 (.DIODE(net463),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output464_A (.DIODE(net464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_5__Q (.DIODE(net464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1788_A1 (.DIODE(net464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1306_B2 (.DIODE(net464),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output465_A (.DIODE(net465),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_6__Q (.DIODE(net465),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1789_A1 (.DIODE(net465),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1364_B2 (.DIODE(net465),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output466_A (.DIODE(net466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_3__Q (.DIODE(net466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1791_A1 (.DIODE(net466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1446_B2 (.DIODE(net466),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output467_A (.DIODE(net467),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_2__Q (.DIODE(net467),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1792_A1 (.DIODE(net467),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1472_B2 (.DIODE(net467),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output468_A (.DIODE(net468),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_4__Q (.DIODE(net468),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1790_A1 (.DIODE(net468),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1233_B2 (.DIODE(net468),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output469_A (.DIODE(net469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_1__Q (.DIODE(net469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1785_A1 (.DIODE(net469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1326_B2 (.DIODE(net469),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output471_A (.DIODE(net471),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_6__Q (.DIODE(net471),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1779_A1 (.DIODE(net471),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1366_A2 (.DIODE(net471),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output472_A (.DIODE(net472),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_7__Q (.DIODE(net472),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1780_A1 (.DIODE(net472),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1288_B2 (.DIODE(net472),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output474_A (.DIODE(net474),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_2__Q (.DIODE(net474),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1784_A1 (.DIODE(net474),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1450_A2 (.DIODE(net474),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output475_A (.DIODE(net475),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_3__Q (.DIODE(net475),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1783_A1 (.DIODE(net475),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1424_A2 (.DIODE(net475),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output476_A (.DIODE(net476),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_5__Q (.DIODE(net476),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1781_A1 (.DIODE(net476),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1309_B2 (.DIODE(net476),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output477_A (.DIODE(net477),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_4__Q (.DIODE(net477),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1819_A1 (.DIODE(net477),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1240_B2 (.DIODE(net477),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output479_A (.DIODE(net479),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_8__Q (.DIODE(net479),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1815_A1 (.DIODE(net479),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1274_B2 (.DIODE(net479),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output480_A (.DIODE(net480),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_9__Q (.DIODE(net480),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1816_A1 (.DIODE(net480),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1223_B2 (.DIODE(net480),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output481_A (.DIODE(net481),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_6__Q (.DIODE(net481),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1817_A1 (.DIODE(net481),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1378_B2 (.DIODE(net481),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output482_A (.DIODE(net482),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_7__Q (.DIODE(net482),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1818_A1 (.DIODE(net482),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1292_B2 (.DIODE(net482),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output485_A (.DIODE(net485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_10__Q (.DIODE(net485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1813_A1 (.DIODE(net485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1187_B2 (.DIODE(net485),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output490_A (.DIODE(net490),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_2__Q (.DIODE(net490),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1922_A1 (.DIODE(net490),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1466_A2 (.DIODE(net490),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output491_A (.DIODE(net491),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_1__Q (.DIODE(net491),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1923_A1 (.DIODE(net491),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1348_B2 (.DIODE(net491),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output492_A (.DIODE(net492),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_0__Q (.DIODE(net492),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1924_A1 (.DIODE(net492),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1412_A2 (.DIODE(net492),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output493_A (.DIODE(net493),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_9__Q (.DIODE(net493),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1914_A1 (.DIODE(net493),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1214_A2 (.DIODE(net493),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output494_A (.DIODE(net494),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_10__Q (.DIODE(net494),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1915_A1 (.DIODE(net494),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1193_B2 (.DIODE(net494),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output495_A (.DIODE(net495),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_3__Q (.DIODE(net495),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1921_A1 (.DIODE(net495),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1440_A2 (.DIODE(net495),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output496_A (.DIODE(net496),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_4__Q (.DIODE(net496),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1920_A1 (.DIODE(net496),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1259_A2 (.DIODE(net496),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output497_A (.DIODE(net497),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_7__Q (.DIODE(net497),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1917_A1 (.DIODE(net497),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1282_A2 (.DIODE(net497),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output498_A (.DIODE(net498),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_5__Q (.DIODE(net498),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1919_A1 (.DIODE(net498),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1322_A2 (.DIODE(net498),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output500_A (.DIODE(net500),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_8__Q (.DIODE(net500),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1916_A1 (.DIODE(net500),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1264_B2 (.DIODE(net500),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output502_A (.DIODE(net502),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_1__Q (.DIODE(net502),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1934_A1 (.DIODE(net502),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1327_A2 (.DIODE(net502),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output504_A (.DIODE(net504),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_8__Q (.DIODE(net504),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1926_A1 (.DIODE(net504),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1273_A2 (.DIODE(net504),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output505_A (.DIODE(net505),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_9__Q (.DIODE(net505),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1927_A1 (.DIODE(net505),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1221_A2 (.DIODE(net505),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output509_A (.DIODE(net509),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_5__Q (.DIODE(net509),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1930_A1 (.DIODE(net509),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1308_A2 (.DIODE(net509),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output511_A (.DIODE(net511),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_4__Q (.DIODE(net511),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2002_A1 (.DIODE(net511),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1247_B2 (.DIODE(net511),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output513_A (.DIODE(net513),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_12__Q (.DIODE(net513),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1994_A1 (.DIODE(net513),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1101_A2 (.DIODE(net513),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output515_A (.DIODE(net515),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_10__Q (.DIODE(net515),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1996_A1 (.DIODE(net515),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1182_A2 (.DIODE(net515),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output516_A (.DIODE(net516),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_11__Q (.DIODE(net516),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1997_A1 (.DIODE(net516),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1138_B2 (.DIODE(net516),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output518_A (.DIODE(net518),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_3__Q (.DIODE(net518),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2005_A1 (.DIODE(net518),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1431_A2 (.DIODE(net518),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output520_A (.DIODE(net520),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_17__Q (.DIODE(net520),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1991_A1 (.DIODE(net520),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1169_A2 (.DIODE(net520),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output521_A (.DIODE(net521),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_14__Q (.DIODE(net521),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1992_A1 (.DIODE(net521),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1175_A2 (.DIODE(net521),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output523_A (.DIODE(net523),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_8__Q (.DIODE(net523),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1998_A1 (.DIODE(net523),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1279_A2 (.DIODE(net523),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output524_A (.DIODE(net524),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_9__Q (.DIODE(net524),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1999_A1 (.DIODE(net524),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1206_A2 (.DIODE(net524),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output525_A (.DIODE(net525),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_6__Q (.DIODE(net525),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2000_A1 (.DIODE(net525),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1371_A2 (.DIODE(net525),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output526_A (.DIODE(net526),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_7__Q (.DIODE(net526),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2001_A1 (.DIODE(net526),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1295_A2 (.DIODE(net526),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output527_A (.DIODE(net527),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_0__Q (.DIODE(net527),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2006_A1 (.DIODE(net527),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1392_A2 (.DIODE(net527),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output540_A (.DIODE(net540),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_13__Q (.DIODE(net540),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1615_A1 (.DIODE(net540),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1148_A1 (.DIODE(net540),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output541_A (.DIODE(net541),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_14__Q (.DIODE(net541),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1616_A1 (.DIODE(net541),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1176_B2 (.DIODE(net541),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output544_A (.DIODE(net544),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_17__Q (.DIODE(net544),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1619_A1 (.DIODE(net544),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1170_B2 (.DIODE(net544),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output545_A (.DIODE(net545),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_17__Q (.DIODE(net545),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1683_A1 (.DIODE(net545),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1167_B2 (.DIODE(net545),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output550_A (.DIODE(net550),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_tempsense_ctrl_REG_reg_0__Q (.DIODE(net550),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1527_A0 (.DIODE(net550),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1269_A2 (.DIODE(net550),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output553_A (.DIODE(net553),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_10__Q (.DIODE(net553),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1600_A1 (.DIODE(net553),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1191_A2 (.DIODE(net553),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output554_A (.DIODE(net554),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_9__Q (.DIODE(net554),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1601_A1 (.DIODE(net554),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1217_A2 (.DIODE(net554),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output555_A (.DIODE(net555),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_1__Q (.DIODE(net555),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1764_A1 (.DIODE(net555),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1351_A2 (.DIODE(net555),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output557_A (.DIODE(net557),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_8__Q (.DIODE(net557),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1756_A1 (.DIODE(net557),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1375_A1 (.DIODE(net557),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output558_A (.DIODE(net558),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_9__Q (.DIODE(net558),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1757_A1 (.DIODE(net558),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1212_B2 (.DIODE(net558),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output559_A (.DIODE(net559),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_6__Q (.DIODE(net559),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1758_A1 (.DIODE(net559),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1376_B2 (.DIODE(net559),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output560_A (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_7__Q (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1759_A1 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1283_A2 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output567_A (.DIODE(net567),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_9__Q (.DIODE(net567),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1767_A1 (.DIODE(net567),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1208_B2 (.DIODE(net567),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output568_A (.DIODE(net568),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_10__Q (.DIODE(net568),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1768_A1 (.DIODE(net568),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1184_B2 (.DIODE(net568),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output569_A (.DIODE(net569),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_7__Q (.DIODE(net569),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1769_A1 (.DIODE(net569),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1299_B2 (.DIODE(net569),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output570_A (.DIODE(net570),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_8__Q (.DIODE(net570),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1770_A1 (.DIODE(net570),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1261_B2 (.DIODE(net570),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output571_A (.DIODE(net571),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_5__Q (.DIODE(net571),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1772_A1 (.DIODE(net571),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1266_B1 (.DIODE(net571),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output575_A (.DIODE(net575),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_6__Q (.DIODE(net575),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1771_A1 (.DIODE(net575),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1400_A1 (.DIODE(net575),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output579_A (.DIODE(net579),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_13__Q (.DIODE(net579),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1688_A1 (.DIODE(net579),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1151_B2 (.DIODE(net579),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output584_A (.DIODE(net584),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_6__Q (.DIODE(net584),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1693_A1 (.DIODE(net584),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1360_B2 (.DIODE(net584),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output588_A (.DIODE(net588),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_2__Q (.DIODE(net588),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2023_A1 (.DIODE(net588),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1455_A2 (.DIODE(net588),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output589_A (.DIODE(net589),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_3__Q (.DIODE(net589),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2024_A1 (.DIODE(net589),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1429_A2 (.DIODE(net589),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output592_A (.DIODE(net592),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_19__Q (.DIODE(net592),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1681_A1 (.DIODE(net592),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1478_A2 (.DIODE(net592),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output593_A (.DIODE(net593),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_20__Q (.DIODE(net593),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1680_A1 (.DIODE(net593),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1143_B2 (.DIODE(net593),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_X (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1992_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1993_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1994_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1995_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1997_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1996_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1998_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1999_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2000_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2001_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2002_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2003_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2004_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2005_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2006_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2007_S (.DIODE(net594),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout595_X (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1973_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1974_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1975_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1976_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1978_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1977_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1979_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1980_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1981_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1982_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1983_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1984_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1985_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1986_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1987_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1988_S (.DIODE(net595),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_X (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1955_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1954_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1956_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1957_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1958_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1959_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1960_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1961_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1962_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1963_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1964_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1965_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1966_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1967_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1968_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1969_S (.DIODE(net596),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout601_X (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1584_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1597_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1598_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1581_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout600_A (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1575_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1578_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1577_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1576_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1574_S (.DIODE(net601),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_X (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1572_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1548_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout602_A (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1549_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1567_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1543_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1544_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1545_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1546_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1547_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1571_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1570_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1569_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1568_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1551_S (.DIODE(net603),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_X (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1519_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1511_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1515_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1509_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1510_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1508_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1507_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1506_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1514_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1513_S (.DIODE(net605),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout606_X (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1432_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1372_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1297_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1182_B1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1141_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1480_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1477_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1406_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1317_B1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1279_B1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1337_B1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2029_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2027_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1483_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1481_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1249_A1 (.DIODE(net606),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_X (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1174_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1168_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1155_A1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1951_A (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1161_A1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1135_A1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1334_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1390_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1314_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1276_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1246_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1179_A1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1147_A1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1125_A1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1429_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1455_B1 (.DIODE(net607),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_X (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1199_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1174_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1146_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1131_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1168_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1154_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1160_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1219_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1363_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1446_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1472_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1122_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1383_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1326_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1286_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1236_A1 (.DIODE(net608),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_X (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1303_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1284_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1230_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1210_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1194_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1360_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1416_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1133_B1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1119_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1151_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1167_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1173_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1642_A (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1469_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1443_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1354_A1 (.DIODE(net609),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_X (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1373_A2 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1323_B1 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1194_B1 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1414_B1 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1259_B1 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1282_B1 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1210_B1 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1353_A1 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_X (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1462_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1611_A (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1345_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1321_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1264_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1109_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1184_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1213_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1298_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1257_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1139_A1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1403_B2 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1409_B1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1176_B1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1170_B1 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1148_A2 (.DIODE(net611),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_X (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1175_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1169_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1206_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1182_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1101_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1989_A (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1457_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1431_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1392_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1371_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1335_B1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1316_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1295_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1279_A1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1247_B1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1138_B1 (.DIODE(net612),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout613_X (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1110_A2 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1157_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1163_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1296_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1479_B1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1461_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1409_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1476_B1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1320_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1185_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1176_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1170_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1150_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1132_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1370_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1435_A1 (.DIODE(net613),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout614_X (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1208_A1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1256_A1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1263_A1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1143_A1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout613_A (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2029_B1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2027_B1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1573_A (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1483_B1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1481_B1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1344_A1 (.DIODE(net614),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_X (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1337_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1476_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1479_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1317_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1262_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1177_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1171_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1162_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1156_A1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1140_B1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout615_A (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1295_B1 (.DIODE(net616),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_A (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1211_A (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_cap617_X (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1229_B (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1350_B (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1251_A (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1207_B (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1237_B (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1235_B (.DIODE(net617),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout619_X (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1296_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1209_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1185_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1164_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1158_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1139_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1110_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1097_C (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2035_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2034_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2033_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1484_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1482_B1 (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1087_A (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1051_B (.DIODE(net619),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_X (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2017_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1642_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1599_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1486_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1850_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1812_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1989_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1661_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1573_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1825_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1804_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1498_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1049_A (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2008_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1542_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1838_B (.DIODE(net620),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_X (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1787_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1778_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1951_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2022_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1711_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1721_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1743_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1874_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1860_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1901_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1795_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1936_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1706_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1679_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1755_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1766_B (.DIODE(net621),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_X (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1887_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1913_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1925_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1970_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_A (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1528_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1732_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1630_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1611_B (.DIODE(net622),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_X (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1891_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1877_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1864_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1840_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1816_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1767_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1757_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1744_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1734_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1723_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1692_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1634_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1627_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1590_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1556_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1539_A0 (.DIODE(net623),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout624_X (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1902_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1914_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1927_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_A (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1999_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1980_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1961_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1942_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1829_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1665_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1658_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1601_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1520_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1488_A0 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout625_X (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1878_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1865_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1851_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1841_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1815_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1756_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1733_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1722_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1713_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1770_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1691_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1633_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1626_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1589_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1555_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1538_A0 (.DIODE(net625),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire627_A (.DIODE(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout626_X (.DIODE(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1998_A0 (.DIODE(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1979_A0 (.DIODE(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1960_A0 (.DIODE(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1828_A0 (.DIODE(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1747_A0 (.DIODE(net626),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire627_X (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1904_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1892_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1926_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1916_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout625_A (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1603_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1489_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1657_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1664_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1519_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1941_A0 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout628_X (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1879_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1866_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1852_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1842_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1818_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1796_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1780_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1712_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1769_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1736_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1694_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1632_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1625_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1588_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1554_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1537_A0 (.DIODE(net628),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire630_A (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout629_X (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2001_A0 (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1982_A0 (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1963_A0 (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1944_A0 (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1831_A0 (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1746_A0 (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1725_A0 (.DIODE(net629),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire630_X (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2010_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1928_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout628_A (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1602_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1759_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1490_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1656_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1663_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1518_A0 (.DIODE(net630),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire631_X (.DIODE(net631),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1893_A0 (.DIODE(net631),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1905_A0 (.DIODE(net631),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1917_A0 (.DIODE(net631),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout629_A (.DIODE(net631),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout632_X (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1880_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1853_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1817_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1805_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1797_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1789_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1779_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1771_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1748_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1735_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1693_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1631_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1624_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1587_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1553_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1536_A0 (.DIODE(net632),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout633_X (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout632_A (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2000_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1981_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1962_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1943_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1867_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1843_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1830_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1758_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1724_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1715_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1662_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1655_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1609_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1517_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1493_A0 (.DIODE(net633),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire634_X (.DIODE(net634),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1894_A0 (.DIODE(net634),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2009_A0 (.DIODE(net634),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1906_A0 (.DIODE(net634),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1918_A0 (.DIODE(net634),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1929_A0 (.DIODE(net634),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout635_X (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1671_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1654_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1608_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1516_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1492_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2012_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2003_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1984_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1965_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1946_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1881_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1868_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1854_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1833_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1820_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1714_A0 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout636_X (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1895_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1806_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1798_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1788_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1781_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1772_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1760_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1749_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1737_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1726_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1696_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1640_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1623_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1586_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1552_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1535_A0 (.DIODE(net636),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire637_X (.DIODE(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1907_A0 (.DIODE(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1919_A0 (.DIODE(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1930_A0 (.DIODE(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout636_A (.DIODE(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1674_A0 (.DIODE(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1844_A0 (.DIODE(net637),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout638_X (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1653_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1551_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1515_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1491_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1048_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2011_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2002_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1983_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1964_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1945_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1882_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1869_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1855_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1845_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1832_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1819_A0 (.DIODE(net638),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout639_X (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1807_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1799_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1790_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1782_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1773_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1761_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1750_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1738_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1727_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1716_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1695_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1639_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1622_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1607_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1585_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1534_A0 (.DIODE(net639),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire640_X (.DIODE(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1896_A0 (.DIODE(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1908_A0 (.DIODE(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1920_A0 (.DIODE(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1931_A0 (.DIODE(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout639_A (.DIODE(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1670_A0 (.DIODE(net640),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout641_X (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1550_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1496_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2005_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1986_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1967_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1948_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1883_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1870_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1856_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1846_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1835_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1822_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1808_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1800_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1676_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1514_A0 (.DIODE(net641),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout642_X (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1921_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1909_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1897_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1791_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1783_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1762_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1728_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1717_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1774_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1751_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1739_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1708_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1698_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1638_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1621_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1533_A0 (.DIODE(net642),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire644_X (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2019_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2014_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2024_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1932_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout642_A (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1584_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1606_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1703_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1652_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1669_A0 (.DIODE(net644),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout645_X (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1549_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1495_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2004_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1985_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1966_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1947_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1884_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1871_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1857_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1847_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1834_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1821_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1809_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1801_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1675_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1513_A0 (.DIODE(net645),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout646_X (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1922_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1910_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1898_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1792_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1784_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1763_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1729_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1718_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1775_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1752_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1740_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1707_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1697_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1637_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1620_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1532_A0 (.DIODE(net646),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire648_X (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2018_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2013_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2023_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1933_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout646_A (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1583_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1605_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1702_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1651_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1668_A0 (.DIODE(net648),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout649_X (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1494_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2016_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2007_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1988_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1969_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1950_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1886_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1873_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1859_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1849_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1837_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1824_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1811_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1803_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1730_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1719_A0 (.DIODE(net649),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout650_X (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1705_A0 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1677_A0 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1667_A0 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1659_A0 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1604_A0 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1582_A0 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1526_A1 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1512_A0 (.DIODE(net650),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout651_X (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1934_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1923_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1793_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1785_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1776_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1764_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1912_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1900_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1753_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1741_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1710_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1699_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1636_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1628_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1548_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1531_A0 (.DIODE(net651),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire652_X (.DIODE(net652),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2021_A0 (.DIODE(net652),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2026_A0 (.DIODE(net652),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout651_A (.DIODE(net652),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout650_A (.DIODE(net652),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire653_X (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1953_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1991_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1972_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1683_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1619_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1564_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1581_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1650_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1502_A0 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire654_X (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1952_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1990_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1971_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1684_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1618_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1563_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1597_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1649_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1501_A0 (.DIODE(net654),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire655_X (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1955_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1993_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1974_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1685_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1617_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1562_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1596_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1648_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1500_A0 (.DIODE(net655),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire656_X (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1954_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1973_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1992_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1686_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1616_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1561_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1595_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1647_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1499_A0 (.DIODE(net656),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire657_X (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1888_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1814_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1978_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1997_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1861_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1876_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1690_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1613_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1541_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1558_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1592_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1644_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1522_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1940_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1959_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1827_A0 (.DIODE(net657),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout658_X (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1768_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1745_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1689_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1635_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1612_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1557_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1540_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1958_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1939_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1826_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1666_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1643_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1600_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1591_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1521_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1487_A0 (.DIODE(net658),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout660_X (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1497_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2015_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2006_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1987_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1968_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1949_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1885_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1872_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1858_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1848_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1836_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1823_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1810_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1802_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1731_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1720_A0 (.DIODE(net660),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout661_X (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1704_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1678_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1672_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1660_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1610_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1598_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1572_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1527_A1 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1524_A0 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout662_X (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2020_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1935_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1924_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1794_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1786_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1777_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1765_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1742_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1911_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1899_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1754_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1709_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1700_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1641_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1629_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1530_A0 (.DIODE(net662),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire663_X (.DIODE(net663),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2025_A0 (.DIODE(net663),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout662_A (.DIODE(net663),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout661_A (.DIODE(net663),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout681_X (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout679_A (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout680_A (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_5__RESET_B (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_6__RESET_B (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_7__RESET_B (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_0__RESET_B (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_tempsense_ctrl_REG_reg_0__RESET_B (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_tempsense_ctrl_REG_reg_1__RESET_B (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout678_A (.DIODE(net681),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout682_X (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout676_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout677_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout674_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout675_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout681_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout667_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout672_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout671_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout673_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_5__RESET_B (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_4__RESET_B (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout670_A (.DIODE(net682),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout703_X (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout696_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout693_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout702_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout699_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout686_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_1__RESET_B (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_iso_REG_reg_0__RESET_B (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_0__RESET_B (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout690_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout687_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout688_A (.DIODE(net703),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload2_A (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_0__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_9__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_7__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_10__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_9__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_8__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_8__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_4__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_9__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_2__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_10__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_2__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_9__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_5__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_10__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_4__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_3__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_2__CLK (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_PCLK_X (.DIODE(clknet_leaf_1_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload3_A (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_4__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_7__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_1__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_7__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_6__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_3__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_6__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_7__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_6__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_8__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_6__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_2__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_5__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_4__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_2__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_6__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_5__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_8__CLK (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_PCLK_X (.DIODE(clknet_leaf_2_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload4_A (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_5__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_3__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_1__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_0__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_8__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_4__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_0__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_5__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_0__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_1__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_5__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_0__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_5__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_7__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_1__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_1__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_7__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_6__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_5__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_0__CLK (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_PCLK_X (.DIODE(clknet_leaf_3_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload5_A (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_2__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_dac_out_REG_reg_4__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_1__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_4__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_1__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_3__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_PCLK_X (.DIODE(clknet_leaf_4_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_15__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_instramp_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_7__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_brownout_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_PCLK_X (.DIODE(clknet_leaf_5_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_8__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_7__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_PCLK_X (.DIODE(clknet_leaf_6_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload9_A (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_8__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_8__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_7__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_2__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_8__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_4__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_7__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_9__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_5__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_4__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_0__CLK (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_PCLK_X (.DIODE(clknet_leaf_7_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload10_A (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_2__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_2__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_7__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_7__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_0__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_3__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_3__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_ref_REG_reg_6__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_idac_REG_reg_1__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_6__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_3__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_8__CLK (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_PCLK_X (.DIODE(clknet_leaf_8_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload11_A (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_2__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_0__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_3__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_test_REG_reg_1__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_9__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_10__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_8__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_9__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_10__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_9__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_9__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_9__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_8__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_PCLK_X (.DIODE(clknet_leaf_9_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload12_A (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_1__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc0_in_REG_reg_5__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_9__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_10__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp1_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_8__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_3__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_10__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_7__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inn_REG_reg_10__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_2__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_15__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_9__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_3__CLK (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_PCLK_X (.DIODE(clknet_leaf_10_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload13_A (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_2__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_9__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_12__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_10__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_1__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_10__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_iso_REG_reg_2__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_iso_REG_reg_1__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_8__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_7__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_3__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_0__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_iso_REG_reg_0__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_9__CLK (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_PCLK_X (.DIODE(clknet_leaf_11_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload14_A (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_9__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_8__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_11__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inn_REG_reg_11__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_8__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_9__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_4__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_10__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_14__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_16__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_17__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_10__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_11__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_17__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_17__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_15__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_8__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp1_out_REG_reg_10__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_7__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_adc1_in_REG_reg_4__CLK (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_PCLK_X (.DIODE(clknet_leaf_12_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload15_A (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_12__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_10__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_12__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_13__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_11__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_9__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_11__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_10__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_9__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_14__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_8__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_inn_REG_reg_7__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_16__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_16__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_15__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_14__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_8__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_PCLK_X (.DIODE(clknet_leaf_13_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload16_A (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_6__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_16__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_11__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_12__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_14__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_17__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_2__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_13__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_13__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_iso_REG_reg_3__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_12__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_7__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_out_REG_reg_13__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_11__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_13__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_12__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_comp0_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_4__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_8__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_6__CLK (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_PCLK_X (.DIODE(clknet_leaf_14_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload17_A (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_15__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_15__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_18__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_14__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_18__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_19__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_19__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_19__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_16__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_20__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_uproj_REG_reg_20__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_11__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_10__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_16__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_14__CLK (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_PCLK_X (.DIODE(clknet_leaf_15_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload18_A (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_ana_REG_reg_1__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_tempsense_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_5__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_12__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_11__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_15__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_17__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_15__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_11__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_9__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_13__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_12__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_12__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_11__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_idac_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_8__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_instramp_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_17__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_right_opamp_ctrl_REG_reg_12__CLK (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_PCLK_X (.DIODE(clknet_leaf_16_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload6_A (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_12__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_16__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_19__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_11__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_12__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_16__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_13__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_ana_REG_reg_3__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_ana_REG_reg_2__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_sio_ana_REG_reg_0__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_0__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_13__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_18__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_16__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_17__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_comparator_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_tempsense_ctrl_REG_reg_1__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_14__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_17__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_14__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_11__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_6__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_left_opamp_ctrl_REG_reg_14__CLK (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_PCLK_X (.DIODE(clknet_leaf_17_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload7_A (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_29__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_26__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_27__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_25__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_25__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_3__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_23__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_23__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_23__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_21__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_21__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_24__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_24__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_21__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_2__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_5__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_22__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_24__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_bandgap_ctrl_REG_reg_22__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_4__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_13__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_7__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_20__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_rdac_ctrl_REG_reg_18__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_20__CLK (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_PCLK_X (.DIODE(clknet_leaf_18_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload8_A (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_11__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_5__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp0_inn_REG_reg_6__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_5__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_0__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_2__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_6__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_out_REG_reg_11__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_8__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_0__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_9__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp3_out_REG_reg_3__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_inp_REG_reg_1__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_3__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_3__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_preamp0_inp_REG_reg_2__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_13__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_22__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp1_out_REG_reg_12__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_1__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_0__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ana_amp2_out_REG_reg_4__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_reg_ibias_ctrl_REG_reg_28__CLK (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_PCLK_X (.DIODE(clknet_leaf_19_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_PCLK_A (.DIODE(clknet_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_PCLK_A (.DIODE(clknet_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_PCLK_X (.DIODE(clknet_0_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload0_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_PCLK_A (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_PCLK_X (.DIODE(clknet_1_0__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_PCLK_A (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_PCLK_X (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1285_B1 (.DIODE(net706),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1217_B1 (.DIODE(net706),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1231_B1 (.DIODE(net706),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1303_B1 (.DIODE(net706),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1721_A (.DIODE(net706),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_Y (.DIODE(net706),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_B (.DIODE(net709),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer5_X (.DIODE(net709),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1470_B1 (.DIODE(net714),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1444_B1 (.DIODE(net714),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1374_A2 (.DIODE(net714),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_rebuffer10_X (.DIODE(net714),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1442_A1 (.DIODE(net716),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1212_B1 (.DIODE(net716),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1283_A1 (.DIODE(net716),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1228_A1 (.DIODE(net716),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1755_A (.DIODE(net716),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone12_Y (.DIODE(net716),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1196_B1 (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1212_A1 (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1115_A1 (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1150_B1 (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1281_B1 (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1132_B1 (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1936_A (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_Y (.DIODE(net717),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1360_B1 (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1151_B1 (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1173_B1 (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1167_B1 (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1143_B1 (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1478_A1 (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1475_A1 (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1679_A (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone14_X (.DIODE(net718),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1118_B (.DIODE(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1120_B (.DIODE(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone13_A (.DIODE(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1331_B (.DIODE(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone15_Y (.DIODE(net719),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1425_B1 (.DIODE(net720),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1385_B1 (.DIODE(net720),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1451_B1 (.DIODE(net720),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1221_B1 (.DIODE(net720),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1240_A1 (.DIODE(net720),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1661_A (.DIODE(net720),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_Y (.DIODE(net720),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1218_B1 (.DIODE(net721),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1286_B1 (.DIODE(net721),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1305_B1 (.DIODE(net721),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1233_A1 (.DIODE(net721),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1363_B1 (.DIODE(net721),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1743_A (.DIODE(net721),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_Y (.DIODE(net721),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_U1198_A (.DIODE(net722),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone17_A (.DIODE(net722),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone2_A (.DIODE(net722),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone16_A (.DIODE(net722),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_clone18_X (.DIODE(net722),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(n1025),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_37 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_38 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_39 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_40 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_41 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_42 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_43 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_44 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_45 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_46 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_47 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_48 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_49 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_50 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_51 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_52 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_53 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_54 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_55 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_56 (.DIODE(n1053),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_57 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_58 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_59 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_60 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_61 (.DIODE(n1072),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_62 (.DIODE(n1072),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_63 (.DIODE(n1072),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_64 (.DIODE(n1072),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_65 (.DIODE(n1087),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_66 (.DIODE(n1098),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_67 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_68 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_69 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_70 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_71 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_72 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_73 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_74 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_75 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_76 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_77 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_78 (.DIODE(n1104),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_79 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_80 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_81 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_82 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_83 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_84 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_85 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_86 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_87 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_88 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_89 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_90 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_91 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_92 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_93 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_94 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_95 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_96 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_97 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_98 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_99 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_100 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_101 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_102 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_103 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_104 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_105 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_106 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_107 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_108 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_109 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_110 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_111 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_112 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_113 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_114 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_115 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_116 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_117 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_118 (.DIODE(n1120),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_119 (.DIODE(n1153),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_120 (.DIODE(n1153),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_121 (.DIODE(n1153),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_122 (.DIODE(n1153),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_123 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_124 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_125 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_126 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_127 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_128 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_129 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_130 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_131 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_132 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_133 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_134 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_135 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_136 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_137 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_138 (.DIODE(n1178),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_139 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_140 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_141 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_142 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_143 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_144 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_145 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_146 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_147 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_148 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_149 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_150 (.DIODE(n1237),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_151 (.DIODE(n1247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_152 (.DIODE(n1247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_153 (.DIODE(n1247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_154 (.DIODE(n1247),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_155 (.DIODE(n1271),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_156 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_157 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_158 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_159 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_160 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_161 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_162 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_163 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_164 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_165 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_166 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_167 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_168 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_169 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_170 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_171 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_172 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_173 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_174 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_175 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_176 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_177 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_178 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_179 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_180 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_181 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_182 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_183 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_184 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_185 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_186 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_187 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_188 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_189 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_190 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_191 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_192 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_193 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_194 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_195 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_196 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_197 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_198 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_199 (.DIODE(n1273),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_200 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_201 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_202 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_203 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_204 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_205 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_206 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_207 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_208 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_209 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_210 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_211 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_212 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_213 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_214 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_215 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_216 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_217 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_218 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_219 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_220 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_221 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_222 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_223 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_224 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_225 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_226 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_227 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_228 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_229 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_230 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_231 (.DIODE(n1326),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_232 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_233 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_234 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_235 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_236 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_237 (.DIODE(net30),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_238 (.DIODE(net198),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_239 (.DIODE(net227),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_240 (.DIODE(net250),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_241 (.DIODE(net262),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_242 (.DIODE(net281),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_243 (.DIODE(net285),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_244 (.DIODE(net301),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_245 (.DIODE(net313),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_246 (.DIODE(net319),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_247 (.DIODE(net461),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_248 (.DIODE(net495),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_249 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_250 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_251 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_252 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_253 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_254 (.DIODE(net560),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_255 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_256 (.DIODE(net627),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_257 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_258 (.DIODE(net653),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_259 (.DIODE(net659),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_260 (.DIODE(net659),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_261 (.DIODE(net661),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_262 (.DIODE(clknet_1_1__leaf_PCLK),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_263 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_264 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_265 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_266 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_267 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_268 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_269 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_270 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_271 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_272 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_273 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_274 (.DIODE(n1046),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_275 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_276 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_277 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_278 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_279 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_280 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_281 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_282 (.DIODE(n1067),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_283 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_284 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_285 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_286 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_287 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_288 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_289 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_290 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_291 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_292 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_293 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_294 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_295 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_296 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_297 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_298 (.DIODE(n1106),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_299 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_300 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_301 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_302 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_303 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_304 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_305 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_306 (.DIODE(n1140),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_307 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_308 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_309 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_310 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_311 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_312 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_313 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_314 (.DIODE(n1166),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_315 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_316 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_317 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_318 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_319 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_320 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_321 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_322 (.DIODE(n1253),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_323 (.DIODE(n1261),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_324 (.DIODE(net164),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_325 (.DIODE(net414),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_326 (.DIODE(net524),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_327 (.DIODE(net610),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_328 (.DIODE(net624),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_329 (.DIODE(net635),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_330 (.DIODE(net716),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_331 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_332 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_333 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_334 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_335 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_336 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_337 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_338 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_339 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_340 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_341 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_342 (.DIODE(n1211),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_343 (.DIODE(net164),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__diode_2 ANTENNA_344 (.DIODE(net319),
    .VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_125 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_141 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_148 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_341 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_377 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_665 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_0_678 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_686 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_709 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_761 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_817 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_873 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_899 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_929 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_0_947 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1201 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1341 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1369 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1425 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1553 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1565 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1621 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1721 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1733 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1761 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1805 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1817 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1833 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1861 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1873 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1917 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1929 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1961 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1973 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1985 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2001 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2013 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2097 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2125 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2181 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2209 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2237 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2265 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2293 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2321 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2377 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2517 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2573 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2685 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2825 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2909 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2937 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_2993 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3021 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3049 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3077 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_3441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_0_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_0_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_137 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_144 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_148 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_162 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_171 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_180 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_186 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_202 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_215 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_227 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_230 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_238 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_283 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_294 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_302 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_316 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_327 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_337 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_343 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_348 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_356 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_360 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_372 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_384 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_410 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_422 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_434 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_451 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_486 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_498 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_544 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_1_556 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_585 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_609 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_782 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_1_883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_887 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_895 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_941 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_949 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1001 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1007 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1169 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1175 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1225 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1287 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1337 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1343 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1399 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1481 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1537 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1649 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1705 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1735 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1761 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1805 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1817 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1861 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1873 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1917 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1929 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_1953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1961 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1973 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1985 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_1997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2041 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2097 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2183 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2295 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2345 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2351 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2401 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2407 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2501 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2519 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2569 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2669 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2681 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2725 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2737 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2849 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2893 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_2961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_1_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_1_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_1_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_1_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_255 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_263 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_268 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_276 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_282 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_294 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_306 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_450 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_462 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_465 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_473 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_495 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_507 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_519 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_552 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_571 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_583 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_634 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_642 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_669 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_748 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_768 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_782 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_794 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_798 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_806 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_826 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_838 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_850 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_854 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_866 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_872 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_876 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_879 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_891 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_904 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_908 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_917 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_969 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_976 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1039 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1042 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1050 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1062 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1074 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1086 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1145 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_1251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1315 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1453 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1477 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1522 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1534 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1553 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1565 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1621 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1679 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1691 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1703 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1707 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_1709 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1715 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1727 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1739 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1751 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1789 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_1813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1827 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1839 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1851 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1863 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_2_1889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1915 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1927 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1957 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_1981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2001 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2026 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2038 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2053 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2078 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2090 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_2_2098 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2149 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2267 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2585 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2648 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_2_2697 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2710 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2751 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_2_2763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2771 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2921 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_2_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_2_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_417 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_428 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_440 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_473 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_480 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_644 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_683 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_691 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_756 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_787 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_795 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_800 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_835 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_908 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_928 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_935 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_947 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_985 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_997 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1005 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1048 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1077 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1092 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1104 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1150 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1162 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1174 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1204 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1216 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1228 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1260 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1272 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1284 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1291 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1296 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1308 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1320 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1345 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1350 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1362 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1368 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1396 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1401 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1407 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1564 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1590 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1598 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1622 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_1657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1683 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_1695 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1739 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1779 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_1793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1917 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1929 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_1953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_1961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_1998 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2010 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2041 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2053 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2061 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2098 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2110 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2122 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2158 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2170 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2178 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2182 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2208 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_3_2216 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2243 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2276 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2288 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2321 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2326 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2338 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2348 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2376 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2388 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2400 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2435 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2447 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2459 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2492 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2504 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2516 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2533 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2540 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2550 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2579 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2591 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2606 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2618 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2628 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2680 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2715 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2727 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2739 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_2745 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2750 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_2762 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2770 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2796 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2803 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2815 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2827 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2839 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_3_2851 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2893 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_2961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_3_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_3_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_3_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_3_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_533 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_576 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_660 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_672 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_684 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_692 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_716 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_733 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_808 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_866 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_907 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_910 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_929 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_975 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1002 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1014 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1026 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1095 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1115 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1141 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1181 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1237 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1252 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1305 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1338 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1343 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1348 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1360 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1423 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1474 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1482 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1502 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1556 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1568 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1609 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1635 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1647 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1661 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1683 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1695 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1734 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1746 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1758 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_1797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1812 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1834 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1842 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_1870 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1904 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1916 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_1928 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_4_1965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_1979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2001 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2030 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2042 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2070 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2097 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2122 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2136 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2144 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2267 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_4_2281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_4_2289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2363 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2375 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2418 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2424 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2488 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2538 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2576 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2588 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2592 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2641 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2683 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2695 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2761 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2767 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2800 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2812 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_4_2824 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2921 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_4_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_4_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_558 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_565 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_605 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_714 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_726 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_772 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_829 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_837 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_909 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_939 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_977 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1005 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1030 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1047 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1060 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1076 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1095 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1116 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1130 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1142 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1148 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1221 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1308 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1320 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1356 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1368 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1382 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1394 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1563 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1578 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1590 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1602 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1641 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_1673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1681 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1691 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1703 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1715 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1727 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1735 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1761 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1795 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1823 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1840 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1860 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_1872 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1880 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_1900 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_1930 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_1934 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1963 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1975 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_1987 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_1999 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2013 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2026 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2038 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2050 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2062 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2084 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2096 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2125 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2141 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2183 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2265 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2374 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_2386 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2424 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2436 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2448 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2456 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2476 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2488 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2500 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2504 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2518 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_2521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2552 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2579 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2606 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2618 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2630 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2674 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2686 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2689 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2739 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2761 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2827 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2839 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_5_2851 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_2902 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2910 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_5_2913 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2919 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2931 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2943 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2955 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_5_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_5_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_5_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_5_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_501 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_633 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_641 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_681 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_694 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_774 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_780 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_815 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_823 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_880 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_909 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_943 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_983 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1003 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1018 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1030 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1046 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1058 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1070 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1082 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1115 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1134 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1146 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1149 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1184 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1267 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1306 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1314 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1346 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1358 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1370 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1403 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1472 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1509 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1533 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1549 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1575 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1609 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1675 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1703 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1707 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1774 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1784 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1796 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_1808 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1830 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1842 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1854 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1866 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_1874 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1915 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_1927 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_1933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1941 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_1981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2001 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2013 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_2021 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2054 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2066 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2078 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2090 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2094 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2110 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2122 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2134 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2146 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2154 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2175 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2187 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2199 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_2265 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2287 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2321 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2346 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2358 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2370 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2378 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2418 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2430 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_2489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_6_2505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2535 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_2541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2549 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2555 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2567 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2579 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2591 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2616 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2628 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2640 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2652 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_6_2661 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_6_2677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2685 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2719 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2733 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2796 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2831 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2843 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2855 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2867 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2894 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2943 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2955 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2967 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2979 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_6_2991 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_6_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_6_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_644 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_656 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_668 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_705 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_717 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_777 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_783 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_809 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_843 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_855 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_867 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_879 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_887 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_899 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_947 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_975 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_987 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_999 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1007 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1053 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1056 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1117 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1126 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1143 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1277 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1287 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1291 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1303 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1315 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1327 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1339 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1343 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1399 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1481 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1537 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1616 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1641 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1655 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_1670 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1678 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1708 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_1720 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_7_1734 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1761 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1775 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1787 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1805 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1817 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_1841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1892 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1918 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1930 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_1942 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_1946 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1972 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1984 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_1996 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2008 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2029 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2061 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2096 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2111 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2123 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2183 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2193 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2207 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2219 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2295 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2302 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2314 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2326 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2338 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2344 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2347 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2351 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2361 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2563 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2577 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2595 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2607 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2619 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_2645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2676 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2771 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2783 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2795 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2814 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2826 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2838 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2850 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2893 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_2905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_2925 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2951 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_7_2963 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_7_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_7_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_7_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_7_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_501 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_609 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_730 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_742 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_754 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_811 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_843 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_880 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_892 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_904 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_922 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_938 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_950 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_962 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_974 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1029 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1091 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1179 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_1257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1296 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1308 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1420 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1453 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1477 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1509 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1533 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1553 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1565 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1621 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_1645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1664 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1676 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1688 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_1700 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1721 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1733 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1789 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1833 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1845 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1901 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_1925 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_1945 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1962 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1974 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_1998 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2010 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2022 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2034 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2042 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2088 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2149 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2165 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2201 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_2209 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_2213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2238 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2246 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2271 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2283 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2295 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2307 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2319 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2476 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_8_2488 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_8_2601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2670 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2682 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2694 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2704 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2765 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2771 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2868 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2880 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2896 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2908 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_8_2916 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_8_2931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_8_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_8_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_573 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_602 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_614 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_627 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_639 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_651 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_663 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_777 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_783 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_836 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_895 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_904 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_920 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_932 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_944 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_970 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_982 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1014 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1018 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1030 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1042 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1054 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_1062 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1117 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1140 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1152 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1164 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1300 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1312 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1324 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1336 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1369 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1377 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1399 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1481 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1537 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1642 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1654 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1666 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1696 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1708 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1720 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1732 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1776 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_1788 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1811 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1823 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1835 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_1858 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1866 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1880 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1892 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1917 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1929 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_1961 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_1973 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_1979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2002 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2014 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2035 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2047 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2059 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2097 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2209 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2295 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2345 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2351 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2364 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2390 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2402 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2438 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2446 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2462 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2477 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2517 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2569 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2642 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2654 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2666 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_2678 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2686 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2689 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2705 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_2741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2837 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2868 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2899 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_9_2907 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_2937 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2954 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_9_2966 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_9_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_9_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_9_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_9_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_501 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_680 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_692 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_726 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_734 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_748 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_811 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_871 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_883 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_895 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_907 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_919 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_949 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_993 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1007 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1019 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1042 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1054 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1066 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1070 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1087 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1091 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1132 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1144 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1183 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1228 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1236 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1266 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1278 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1308 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1356 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1368 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1400 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1412 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1424 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1453 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1467 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1479 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1530 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1538 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1572 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1584 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1611 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1619 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1622 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_1657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1662 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1670 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1675 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1682 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1694 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_1706 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1726 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1738 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1750 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_1785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1802 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1814 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1833 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1848 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1901 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_1924 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1957 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_1981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2001 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2013 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2097 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2109 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2145 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2237 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2260 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2420 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2432 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2502 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2514 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2526 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2538 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2546 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2592 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2670 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2682 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2694 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_10_2706 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2714 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2765 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2771 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2773 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2789 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_10_2825 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2864 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2868 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_10_2923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2927 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_10_2941 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2966 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2978 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_2990 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_10_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_10_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_302 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_314 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_326 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_334 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_563 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_596 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_608 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_652 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_658 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_670 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_697 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_777 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_783 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_895 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_921 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_945 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_973 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_977 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_980 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_992 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1004 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1089 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1107 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1145 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1199 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1235 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1337 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1341 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1354 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1366 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1378 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1390 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1398 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1451 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1580 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1638 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1641 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1690 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1702 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1710 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1735 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1768 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1780 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1805 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1817 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_1841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_1893 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_1911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1934 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1946 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1958 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_1961 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_1973 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_1998 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2004 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2075 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2087 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2183 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2208 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2220 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2232 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2284 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2292 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2322 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2334 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2346 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_2361 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2366 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2378 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2390 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2402 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2440 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2452 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2465 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2495 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2507 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2519 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2533 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2562 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2570 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2586 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2598 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2610 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2624 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2669 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2681 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2725 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2737 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_11_2740 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2751 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_11_2801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2807 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2819 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2831 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2843 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_2857 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_2865 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2906 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_2961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_11_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_11_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_11_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_11_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_504 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_516 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_528 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_533 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_577 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_585 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_616 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_620 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_697 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_728 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_740 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_752 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_784 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_796 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_808 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_844 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_856 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_884 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_896 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_904 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_925 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_930 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_942 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_954 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1001 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1013 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1085 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1089 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1118 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1130 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1142 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1149 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1243 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1255 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1306 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1314 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1394 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1398 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1406 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1418 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1426 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1436 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1518 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1530 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1538 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_1583 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1591 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1606 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1612 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_1709 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1740 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1752 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_1765 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1771 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1783 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1795 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1807 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1834 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1846 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1858 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1870 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1914 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1926 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_1957 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_1969 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1982 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_1998 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2004 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2027 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2039 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2049 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2076 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2088 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2096 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2108 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2127 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_2139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2181 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2187 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2199 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2207 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2224 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2236 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2244 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2293 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2312 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2333 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2417 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2462 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_2470 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2486 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2517 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2540 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_12_2573 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_2601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_12_2651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2677 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_12_2713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2717 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2739 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2775 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2831 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2843 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2855 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2867 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_12_2879 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2892 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2904 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2916 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2928 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_12_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_12_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_473 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_543 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_580 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_652 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_658 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_686 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_698 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_706 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_724 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_747 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_787 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_799 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_811 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_823 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_865 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_890 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_921 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_949 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_977 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_985 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1018 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1030 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1042 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1046 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1060 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1115 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1175 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1193 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1201 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1206 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1235 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1271 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1283 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1287 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1293 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1333 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1341 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1345 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1366 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1378 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1390 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1396 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1401 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1408 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1416 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1452 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1486 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1498 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_1510 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1537 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1549 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1555 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1562 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1636 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1648 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1660 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1672 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1780 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1811 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1819 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1831 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1843 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1861 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1873 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_1885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_1905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_1926 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1944 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1956 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_1961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_1965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_1998 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2010 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2029 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2055 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2097 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2137 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2162 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2174 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2182 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2263 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2271 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2290 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2355 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2367 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2379 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2391 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2403 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2407 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2438 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2450 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2462 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2559 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2571 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2654 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2664 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2683 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2689 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_13_2717 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2745 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_2849 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_13_2893 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2909 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2913 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2921 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_2933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_2959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_13_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_13_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_13_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_13_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_458 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_470 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_477 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_491 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_503 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_515 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_527 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_544 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_556 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_582 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_631 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_669 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_675 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_687 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_748 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_789 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_809 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_825 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_893 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_917 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_925 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_946 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_958 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_970 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_978 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1026 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1034 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1067 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1079 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1091 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1122 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1134 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1146 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1151 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1159 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1180 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1192 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1222 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1243 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1255 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1305 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1384 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1396 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1408 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1420 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1453 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1465 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1536 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1609 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1640 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1682 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1694 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1706 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1721 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1733 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_1745 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1751 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1765 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1791 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_1803 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1832 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1844 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1856 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1868 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_1889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1910 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_1922 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_1930 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1960 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1972 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_1984 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_1991 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2003 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2040 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2056 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2068 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2080 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2092 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2145 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2188 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2200 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2208 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2237 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2258 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2266 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2294 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2355 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2367 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2389 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2419 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2431 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2478 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2490 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2536 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2585 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_14_2629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2652 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_14_2709 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_14_2734 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2748 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2760 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_2885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2921 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_14_2933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2937 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_2950 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2972 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2984 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_14_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_14_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_460 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_468 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_486 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_498 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_585 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_609 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_615 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_642 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_654 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_666 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_777 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_796 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_808 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_820 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_832 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_899 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_911 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_929 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_945 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1001 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1005 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1019 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1031 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1043 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1055 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1170 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1218 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1287 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1307 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1319 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1327 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1343 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1375 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1387 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1399 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1401 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1553 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1565 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1654 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1666 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1690 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1702 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1714 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1726 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_1734 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1761 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_1805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1809 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1837 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1861 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1873 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_1885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_1923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_1929 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_1957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1961 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1973 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1985 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_1997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2059 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2097 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2141 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2183 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2299 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2311 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2323 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2344 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2377 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2383 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2406 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2462 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2514 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2633 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2643 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2655 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2682 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2702 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2714 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2726 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2738 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2840 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2852 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_2905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2913 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_2921 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_15_2947 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2951 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_15_2963 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_15_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_15_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_15_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_15_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_450 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_462 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_474 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_501 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_620 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_634 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_642 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_669 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_693 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_709 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_796 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_808 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_908 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_920 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_952 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_964 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_976 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1024 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1085 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1091 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1141 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1167 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1179 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1191 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1223 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1235 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1247 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1267 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1286 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1298 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1310 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1342 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1354 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1366 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1436 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1444 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1509 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1543 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1555 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1567 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1579 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1591 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1621 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1665 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_1701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1718 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1730 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1742 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_1754 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1762 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1789 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_1813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1839 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1851 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1863 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1907 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1919 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_1933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1948 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1960 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1972 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_1984 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2001 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2015 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2027 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_2039 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2069 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2149 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2165 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2170 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2182 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2194 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2225 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2235 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2247 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2267 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2401 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2422 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_2485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2511 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2523 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2535 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2549 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2557 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_2573 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2629 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2641 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_2661 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2685 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2698 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2710 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2717 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2734 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2746 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2758 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_2770 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_2785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2814 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_16_2826 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2829 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2835 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2863 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_2885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2891 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2915 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_16_2927 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_16_2935 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2941 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2967 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2979 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_16_2991 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_16_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_16_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_417 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_573 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_577 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_598 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_610 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_627 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_639 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_651 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_663 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_669 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_694 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_731 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_743 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_755 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_767 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_779 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_783 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_837 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_866 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_878 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_895 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_921 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_945 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_987 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_999 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1020 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1032 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1044 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1056 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1090 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1102 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1112 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1170 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1227 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1274 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1286 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1323 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1343 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1367 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1376 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1388 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1406 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1452 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1481 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_1513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1547 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1565 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1571 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1583 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1595 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1607 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1619 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1649 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1694 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1721 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_1733 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1761 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1820 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_1846 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1861 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1873 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1917 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1929 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_1953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1972 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_1984 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_1996 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2000 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2026 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2038 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2050 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2062 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2070 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2085 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2118 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2126 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2183 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2193 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2235 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2250 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2262 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2274 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2286 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2294 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2305 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2308 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2320 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2332 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2344 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2355 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2389 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2493 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2517 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2569 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2577 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2615 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2627 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2633 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2639 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2662 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2674 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2682 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2686 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2716 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2728 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_17_2740 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2790 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2798 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2815 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_2853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2857 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_2865 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_2904 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2934 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2946 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_2958 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_17_2966 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_17_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_17_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_17_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_17_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_456 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_468 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_471 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_509 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_574 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_586 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_656 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_671 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_750 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_832 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_840 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_856 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_902 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_914 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_994 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1006 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1047 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1083 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1091 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1130 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1162 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1174 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1186 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1198 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1221 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1227 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1255 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1305 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1404 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1431 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1436 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1447 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1459 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1471 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1507 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1519 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1535 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1621 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1646 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1665 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_1680 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1721 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1733 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1774 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1786 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1798 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1810 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1818 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1851 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_1867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1901 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1913 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_1930 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_1968 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_1980 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_1998 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2002 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2034 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_2042 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2069 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2081 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2128 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2140 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2152 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2167 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_2179 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2194 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2206 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2225 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2256 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_2281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2306 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2320 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_2393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2423 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_2469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2484 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2493 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_2545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2585 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2616 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2628 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2640 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_2657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2661 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2665 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2670 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2696 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_2708 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2717 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2738 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_18_2746 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_18_2762 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_2770 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2829 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2868 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2880 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_18_2897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2914 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2926 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_18_2938 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_18_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_18_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_333 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_337 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_354 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_366 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_383 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_420 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_424 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_511 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_523 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_550 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_579 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_591 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_619 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_635 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_767 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_779 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_783 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_835 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_895 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_927 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_939 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_966 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1021 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1033 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1059 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1086 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1094 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1151 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1164 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1210 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1222 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1230 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_1285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1324 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1336 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1388 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1410 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1422 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1434 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1451 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1481 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1547 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1607 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1619 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1649 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1705 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1735 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1737 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1761 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_1785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1805 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1817 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1829 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1860 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1872 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1884 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1896 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1939 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_1961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_1965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_1975 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_1995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_2012 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2033 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2052 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2097 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2117 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_2125 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_2141 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2178 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_19_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2227 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_2235 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2295 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2345 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2351 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_2365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2392 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_2404 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2465 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_2517 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2544 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2556 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2568 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_2625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2698 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_2710 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2718 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2747 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_2797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2849 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2893 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_2905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_19_2961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_2965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_2994 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3006 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3018 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_19_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_19_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_19_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_19_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_332 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_392 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_396 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_477 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_482 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_566 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_578 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_586 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_619 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_631 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_686 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_698 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_740 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_750 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_761 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_824 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_863 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_880 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_892 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_904 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_910 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_937 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_960 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_972 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_988 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_992 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1018 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1024 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1032 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1050 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1058 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1063 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1089 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1112 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1120 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1138 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1146 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1200 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1258 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1266 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1279 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1291 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1299 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1312 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1328 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1340 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1352 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1364 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1406 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1418 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1426 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1438 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1442 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1482 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1493 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1507 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1519 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1552 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1555 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1567 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1579 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1591 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_1621 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1646 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1677 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1707 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1721 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1733 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1789 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1833 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1845 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_1869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1910 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1922 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1930 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1935 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_1957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_1975 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_1999 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2019 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_2022 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2026 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_2042 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_2057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2070 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_2149 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2166 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2178 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2190 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2202 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_2210 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2225 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2260 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2302 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2314 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_2322 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_2353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_2389 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2406 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2418 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2430 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_2517 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_2581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2585 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2609 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_20_2617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2675 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2703 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_2765 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2771 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2782 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_20_2794 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2798 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_20_2826 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2921 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_2933 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2941 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2949 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2963 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2975 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_20_2987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_20_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_20_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_305 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_339 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_356 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_368 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_473 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_524 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_558 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_594 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_615 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_635 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_658 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_705 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_717 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_774 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_782 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_810 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_822 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_834 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_857 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_880 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_892 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_921 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_945 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_966 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_978 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_990 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1002 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1027 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1039 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1051 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1103 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1213 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1225 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1284 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1306 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1314 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1330 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1342 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1348 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1389 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1404 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1416 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1422 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1430 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1459 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1471 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1483 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1495 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1507 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1528 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1544 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1564 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_1617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1638 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1650 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1662 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1670 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1693 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1712 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1724 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1749 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1761 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1773 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1795 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1807 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1819 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1831 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_1843 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1861 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_1893 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1917 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_1953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_1968 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_2041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_2049 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2082 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2094 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2106 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2118 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2140 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2152 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2164 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_2176 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_2253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2280 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_2292 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_2349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_2365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_2405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_2409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2434 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2446 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2458 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_2465 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_21_2473 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2499 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2519 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2548 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2560 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_2572 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2577 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2633 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_2674 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_2679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2691 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2703 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2732 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_2757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_2786 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2794 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2812 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_2824 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2830 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2859 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2871 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2883 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2895 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_2907 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_21_2937 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_2981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_3021 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_21_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_21_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_21_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_21_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_336 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_348 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_360 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_392 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_404 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_416 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_462 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_479 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_491 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_503 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_515 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_527 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_548 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_560 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_572 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_656 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_678 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_690 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_726 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_742 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_784 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_788 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_818 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_830 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_834 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_850 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_862 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_917 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_971 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1029 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1035 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1110 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1126 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1162 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1174 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1221 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1255 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1306 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1314 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1370 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1467 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1479 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1509 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1533 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1553 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1565 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1605 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1630 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1642 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1650 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1674 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1686 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1698 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1706 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1721 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1733 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1756 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1774 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1786 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_1794 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1833 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1845 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_1869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1873 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1886 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1898 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1910 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_1922 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1935 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1947 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_1979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2001 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_2009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2013 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_2069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2075 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2087 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_2147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2186 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_2198 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2206 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2224 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2236 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2248 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2260 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2280 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2292 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2298 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2327 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2339 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2351 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2363 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_2375 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2418 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2430 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2459 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2471 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_2483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_2505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2522 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2534 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_2572 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2611 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_22_2632 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2640 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_2729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2758 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_2770 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_22_2797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2803 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2815 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_2877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_22_2885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2916 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2943 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2955 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_2967 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_22_2979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3022 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3034 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3046 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_22_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_22_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_333 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_400 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_412 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_424 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_436 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_444 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_462 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_474 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_486 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_498 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_585 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_590 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_598 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_614 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_629 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_641 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_658 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_670 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_697 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_717 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_753 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_762 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_773 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_781 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_853 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_865 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_899 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_911 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_923 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_935 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_947 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_979 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_991 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1006 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1109 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1112 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1169 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1175 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1196 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1208 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1220 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1244 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1256 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1268 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1280 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1334 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1342 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1399 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1455 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1481 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1537 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1605 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1621 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1681 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1686 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1698 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1710 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1739 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1751 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1763 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1775 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1787 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_1837 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_1849 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1862 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1874 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1886 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1898 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1905 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1917 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1929 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_1953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1961 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1973 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1985 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_1997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2041 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2097 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_2181 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_2197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2230 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_2264 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2290 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_2309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2342 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2348 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2351 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2364 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2376 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2388 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2400 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2501 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2519 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_2559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2577 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2622 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_2630 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_2633 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2670 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2682 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2702 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2714 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2722 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2736 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2766 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2778 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_2786 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2839 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_2851 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2857 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_2881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2915 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2927 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2939 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_2951 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_23_2963 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_2969 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_23_2977 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_2990 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3016 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_23_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_23_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_23_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_23_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_411 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_501 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_589 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_601 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_637 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_811 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_837 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_859 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_906 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_918 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_949 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1029 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1035 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1051 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1085 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1089 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1104 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1130 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1142 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1175 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1187 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1199 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1248 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1315 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1341 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1351 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1371 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1463 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1497 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1528 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1621 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1633 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1661 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1677 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1707 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1709 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1732 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1744 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1756 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1795 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_1800 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1815 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1869 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_1909 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1927 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_1957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1963 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_1979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2015 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2027 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2039 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2069 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2125 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2130 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2135 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2169 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2209 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2232 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2238 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2250 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2262 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2320 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2428 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2487 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2493 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2514 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2526 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2538 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2542 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2629 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2641 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_2685 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_24_2714 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2753 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2771 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2817 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2825 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_2885 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2891 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2914 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2935 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_2966 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_2974 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2988 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_24_2997 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3001 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_24_3041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_24_3049 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_24_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_24_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_237 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_273 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_335 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_339 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_351 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_363 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_375 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_393 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_405 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_473 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_585 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_611 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_644 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_664 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_697 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_777 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_783 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_863 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_875 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_887 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_895 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_897 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_909 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_921 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_949 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_970 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_999 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1005 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1027 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1106 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1130 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1142 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1154 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1179 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1191 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1203 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1215 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1227 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1294 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1302 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1326 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1338 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1369 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_1421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1436 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1487 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1499 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1511 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1513 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1525 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1529 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1538 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1550 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1583 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1595 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1618 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1668 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1704 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1716 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1728 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1771 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1783 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_1793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_1801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1819 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1831 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_1843 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1861 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1873 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_1905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1936 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1948 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_1961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1982 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_1994 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2006 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_2014 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2039 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2051 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_2079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2096 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2108 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2120 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2129 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_2169 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2176 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2187 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_2190 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_2209 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2243 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2255 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2267 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2279 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2295 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2306 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2318 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2330 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2342 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_2350 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2374 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2386 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2398 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2432 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_2444 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2448 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2525 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2537 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2549 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_2572 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2577 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2600 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2612 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2624 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_2633 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2649 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_2685 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2725 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2737 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2745 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_25_2777 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2794 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2849 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2857 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2871 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2883 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_25_2895 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_2903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_2981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3000 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3012 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_25_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_25_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_25_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_25_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_265 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_305 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_322 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_348 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_360 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_389 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_426 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_440 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_452 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_464 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_516 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_528 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_542 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_573 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_585 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_619 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_631 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_707 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_730 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_742 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_754 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_769 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_781 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_811 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_825 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_837 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_849 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_866 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_893 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_908 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_920 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_952 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_964 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_974 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1027 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1082 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1090 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1096 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1108 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1120 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1132 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1144 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1185 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1226 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1238 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1250 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1258 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1283 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1295 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1315 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1347 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1367 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1400 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1412 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1424 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1461 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1473 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1522 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1532 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1560 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1564 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1578 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1590 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1627 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1639 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1653 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1677 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1718 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1730 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1742 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1754 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_1762 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1765 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1777 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1789 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1813 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_1828 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1844 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1856 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1868 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1889 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1909 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1915 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_1927 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1933 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1945 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1957 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_1981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2001 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_2013 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_2021 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_2035 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2069 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2134 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_2146 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_2154 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2169 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_2203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_2213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2228 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2240 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2252 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_2264 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2325 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2349 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2381 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_2393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2429 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_26_2482 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_26_2490 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2493 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2505 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2517 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2549 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2555 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2576 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2588 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_2600 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2617 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_2629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2673 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2685 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2697 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2709 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_26_2769 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2868 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_2880 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2885 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_26_2897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2928 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2965 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2977 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_2997 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3009 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3021 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_26_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_26_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_225 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_237 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_264 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_276 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_337 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_342 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_354 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_366 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_378 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_390 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_431 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_470 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_482 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_490 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_557 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_576 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_588 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_600 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_612 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_640 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_652 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_665 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_671 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_681 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_697 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_737 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_753 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_761 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_778 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_815 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_827 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_839 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_893 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_928 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_940 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_970 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_982 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_995 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1007 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1022 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1027 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1033 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1101 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1119 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1157 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1169 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1175 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1201 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1207 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1230 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1245 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1287 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1295 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1315 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1327 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1339 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1354 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1366 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1378 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1425 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1457 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1469 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1507 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_1541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1553 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1565 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1581 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1593 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1625 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1637 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1649 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1661 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1681 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1693 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1726 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1734 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1767 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1779 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1793 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1805 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1823 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1835 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1849 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1861 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1873 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_1881 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_1897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_1909 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1917 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1929 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1941 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_1953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1972 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1984 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_1996 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2008 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2017 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2029 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_2041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_2045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2053 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2073 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2085 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2097 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2110 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_2122 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_2137 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2152 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2164 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_2176 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_2233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2271 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2283 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2295 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2297 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2321 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_2345 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2351 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2353 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_2387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_2453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_2459 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_2515 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2519 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2521 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2533 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2545 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2557 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_2569 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_27_2577 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2585 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2597 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2609 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2621 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2633 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2668 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2680 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2701 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2713 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2725 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_2737 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_2756 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_2797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2801 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2813 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2825 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_27_2833 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2848 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_2857 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2863 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2877 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_2903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2913 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2925 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2937 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2949 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_2961 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2981 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_2993 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3005 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3017 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3025 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3049 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3061 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_27_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_27_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_27_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_27_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_209 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_221 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_229 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_267 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_276 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_288 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_307 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_348 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_360 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_365 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_377 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_401 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_405 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_417 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_474 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_477 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_521 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_527 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_544 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_556 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_584 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_603 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_615 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_627 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_669 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_696 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_712 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_750 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_784 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_807 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_811 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_815 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_831 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_843 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_855 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_869 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_881 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_918 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_936 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_948 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_956 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_966 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_978 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1004 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1012 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1020 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1052 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1064 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1070 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1084 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1117 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1137 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1141 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1181 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1203 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1257 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1278 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1290 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1298 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1352 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1364 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1394 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1406 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1414 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1438 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1454 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1466 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1474 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1479 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1485 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1492 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1504 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1516 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1528 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1541 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1568 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1580 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1592 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1597 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1621 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1629 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1635 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1640 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1665 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1683 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_1697 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_1705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_1713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1717 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1729 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1741 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1778 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1790 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1802 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1814 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1821 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1833 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_1864 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1877 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1921 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1942 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1946 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_1969 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1972 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_1984 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_1989 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2001 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2013 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2030 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2038 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2052 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2082 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_2094 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2137 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2163 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2175 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2187 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2199 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2253 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2265 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2269 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2281 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2327 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2339 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2351 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2377 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2406 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2433 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2437 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2449 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_28_2461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2465 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2477 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2489 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2493 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2501 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2529 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2584 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2596 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2605 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2645 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2674 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2682 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2689 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2750 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2756 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2773 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2785 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2797 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2809 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2829 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2887 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2899 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2911 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_2923 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_28_2935 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2941 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_2979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2985 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_28_2988 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_2997 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3032 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_28_3044 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3189 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3201 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_28_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_28_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_217 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_225 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_312 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_324 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_362 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_366 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_399 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_411 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_474 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_482 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_494 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_502 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_514 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_544 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_556 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_660 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_673 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_691 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_740 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_808 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_852 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_868 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_908 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_912 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_940 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_953 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1003 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1007 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1013 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1025 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1055 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1150 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1162 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1174 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1208 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1220 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1248 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1260 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1272 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1298 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1310 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1315 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1339 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1354 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1358 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1372 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1401 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1414 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1422 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1432 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1438 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1466 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1495 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1507 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1513 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1534 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1546 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1552 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1564 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1569 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1581 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1602 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1614 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1622 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1636 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1679 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1681 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1728 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_1785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1831 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_1897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_1914 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_1922 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_1948 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2001 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_2004 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_2012 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2037 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_2049 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2073 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2089 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2095 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2131 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2137 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2178 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_2204 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2208 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2222 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2234 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2241 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_2280 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2324 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2347 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_2350 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2380 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_2392 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_2400 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2407 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_2441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2490 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2496 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_2512 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2523 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_2535 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2543 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2566 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2579 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2585 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2613 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_2625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_2642 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2648 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_2756 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2786 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_2798 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_2801 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_2806 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2841 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2895 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_2907 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_29_2913 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_2919 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2925 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_29_2964 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_2969 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_2981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3010 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_3018 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3033 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3045 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3057 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_3077 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3081 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3093 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3105 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3117 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3161 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3173 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3193 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3205 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3217 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3229 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3241 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3249 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3261 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3273 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3285 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_29_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_29_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_29_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_29_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_197 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_209 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_213 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_293 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_305 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_309 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_351 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_363 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_407 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_447 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_471 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_500 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_506 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_516 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_544 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_556 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_562 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_591 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_603 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_615 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_643 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_647 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_683 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_695 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_725 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_730 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_733 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_747 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_751 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_784 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_871 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_883 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_936 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_948 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_996 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1008 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1012 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1039 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1051 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1143 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1149 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1178 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1254 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1261 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1265 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1337 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1375 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1480 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1485 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1497 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1535 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1539 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1541 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1549 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1574 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1586 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_1617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1642 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1650 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1657 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1680 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1692 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1704 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1709 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1737 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1790 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1798 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1832 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1840 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_1871 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_1890 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1896 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1919 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_1927 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_1935 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_1947 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1955 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1964 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_1978 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_2041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_2045 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2053 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_2096 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2123 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_2154 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2179 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_2191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_2235 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_2243 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2284 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_2398 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_2437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_2483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_2493 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2551 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2576 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2588 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_2600 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_2605 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_30_2613 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2654 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_2661 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2688 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2728 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2735 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2760 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_2773 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2844 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_2887 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_30_2899 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_2977 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_2997 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3050 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3053 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3065 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3077 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3089 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3101 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3133 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3145 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3195 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3198 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_30_3210 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_30_3218 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3221 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3233 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3245 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3257 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3277 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3289 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3301 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3313 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_30_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_30_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_181 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_193 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_202 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_279 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_301 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_337 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_355 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_377 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_395 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_475 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_509 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_514 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_546 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_553 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_579 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_591 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_615 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_623 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_646 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_661 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_667 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_688 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_693 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_701 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_721 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_837 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_853 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_859 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_867 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_889 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_893 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_917 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_930 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_938 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_945 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_951 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_957 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_986 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_998 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1006 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1009 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1016 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1035 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1057 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1063 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1065 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1085 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1095 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1113 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1165 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1173 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1179 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1201 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1231 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1255 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1259 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1262 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1274 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1281 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1309 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1333 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1339 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1343 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1347 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1354 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1360 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1373 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1395 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1399 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1409 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1421 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1464 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_1476 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1503 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1507 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1536 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1567 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1571 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1587 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1600 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1612 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1618 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1621 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1627 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1648 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1683 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1688 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1696 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1699 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1707 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1749 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1753 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1778 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1784 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1789 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1797 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1800 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1806 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_1815 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1834 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1840 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1845 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1887 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1890 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1898 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_1905 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1912 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1918 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1923 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_1938 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_1946 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1954 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1963 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_1968 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_1999 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2008 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2021 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_2052 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2058 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2077 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2110 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2114 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2122 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2125 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_2129 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2136 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2144 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2147 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2170 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2178 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2181 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2185 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_2205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2230 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2283 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2293 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2297 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2342 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2369 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2398 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2407 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_2416 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2420 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_2444 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2450 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2462 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2465 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2472 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2478 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2483 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_2494 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2519 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2523 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2552 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2568 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2579 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2584 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2592 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2595 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2610 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2618 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2626 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2635 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2641 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2651 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2664 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2685 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2693 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2724 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_2730 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2738 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_2745 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2752 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2758 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_2765 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2771 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2793 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2803 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2810 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2859 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2893 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2900 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2906 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2915 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_31_2948 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2956 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2962 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2971 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_2976 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2982 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2989 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_2999 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3011 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3029 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3041 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3061 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3068 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3072 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3083 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3090 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3094 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3114 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3122 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3128 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3144 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3150 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3170 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3178 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3184 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3193 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_31_3226 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3234 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3240 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3251 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3256 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3262 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3267 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3279 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3291 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3303 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3329 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3341 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3353 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3359 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3385 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3397 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_31_3409 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_31_3415 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3441 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_31_3453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_31_3461 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_189 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_249 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_269 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_285 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_311 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_317 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_383 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_397 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_425 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_453 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_551 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_563 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_593 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_605 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_647 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_719 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_733 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_821 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_873 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_887 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_901 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_929 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_941 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_953 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_965 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_976 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_979 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_981 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1055 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1095 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1109 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1123 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1157 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1209 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1223 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1237 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1265 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1277 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1293 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1319 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1375 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1391 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1403 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1419 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1425 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_1433 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1445 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_8 FILLER_0_32_1473 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1481 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_1487 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1493 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_32_1545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1559 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1573 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_32_1711 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1727 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1739 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1751 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_1763 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3283 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3295 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3307 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3319 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3331 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3357 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3369 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_3381 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3387 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3413 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3425 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_3437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_32_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_32_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_27 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_29 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_41 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_53 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_81 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_85 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_97 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_109 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_137 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_141 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_153 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_165 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_181 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_197 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_225 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_253 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_283 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_313 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_337 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_365 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_393 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_421 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_449 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_477 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_505 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_537 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_561 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_589 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_617 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_649 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_677 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_705 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_729 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_757 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_785 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_815 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_841 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_873 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_897 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_925 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_977 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_985 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1011 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1037 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1069 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1093 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1121 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1153 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1177 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1205 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1233 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1265 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1289 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1321 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1349 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1377 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1427 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1437 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_1443 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1469 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1517 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1545 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1573 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1601 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1625 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1653 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1685 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1713 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_1741 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1745 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_1759 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1791 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1819 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1847 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1875 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1903 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1931 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1959 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_1987 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2015 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2043 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2071 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2099 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2127 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2155 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2183 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2211 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2239 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2267 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2295 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2323 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__decap_4 FILLER_0_33_2325 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2351 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2379 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2407 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2435 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2491 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2519 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2547 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2575 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2603 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2631 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2659 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2687 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2715 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2743 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2771 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2799 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2827 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2855 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2883 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2911 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2939 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2967 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_2995 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3023 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3051 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3079 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3107 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3135 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3163 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3191 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3219 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3247 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3275 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3290 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__fill_2 FILLER_0_33_3302 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3305 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3317 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3329 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3333 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3345 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3357 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3361 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3373 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3385 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3389 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3401 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3413 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3417 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3429 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_3 FILLER_0_33_3441 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3445 (.VPWR(vccd0),
    .VGND(vssd0),
    .VPB(vccd0),
    .VNB(vssd0));
 sky130_fd_sc_hd__decap_6 FILLER_0_33_3457 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
 sky130_fd_sc_hd__fill_1 FILLER_0_33_3463 (.VGND(vssd0),
    .VNB(vssd0),
    .VPB(vccd0),
    .VPWR(vccd0));
endmodule
