module analog_routes ();
endmodule