module usb_cdc_wrapper_ahbl (HCLK,
    HREADY,
    HREADYOUT,
    HRESETn,
    HSEL,
    HWRITE,
    dn_rx_i,
    dn_tx_o,
    dp_pu_o,
    dp_rx_i,
    dp_tx_o,
    irq,
    tx_en_o,
    usb_cdc_clk_48MHz,
    VPWR,
    VGND,
    HADDR,
    HRDATA,
    HSIZE,
    HTRANS,
    HWDATA);
 input HCLK;
 input HREADY;
 output HREADYOUT;
 input HRESETn;
 input HSEL;
 input HWRITE;
 input dn_rx_i;
 output dn_tx_o;
 output dp_pu_o;
 input dp_rx_i;
 output dp_tx_o;
 output irq;
 output tx_en_o;
 input usb_cdc_clk_48MHz;
 inout VPWR;
 inout VGND;
 input [31:0] HADDR;
 output [31:0] HRDATA;
 input [2:0] HSIZE;
 input [1:0] HTRANS;
 input [31:0] HWDATA;

 wire CG_REG_0_;
 wire CONTROL_REG_0_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire \ICR_REG[0] ;
 wire \ICR_REG[1] ;
 wire \ICR_REG[2] ;
 wire \ICR_REG[3] ;
 wire \ICR_REG[4] ;
 wire \ICR_REG[5] ;
 wire \IM_REG[0] ;
 wire \IM_REG[1] ;
 wire \IM_REG[2] ;
 wire \IM_REG[3] ;
 wire \IM_REG[4] ;
 wire \IM_REG[5] ;
 wire N26;
 wire N27;
 wire N28;
 wire N29;
 wire N30;
 wire N31;
 wire \RIS_REG[0] ;
 wire \RIS_REG[1] ;
 wire \RIS_REG[2] ;
 wire \RIS_REG[3] ;
 wire \RIS_REG[4] ;
 wire \RIS_REG[5] ;
 wire \RXFIFOLEVEL_REG[0] ;
 wire \RXFIFOLEVEL_REG[1] ;
 wire \RXFIFOLEVEL_REG[2] ;
 wire \RXFIFOLEVEL_REG[3] ;
 wire \TXFIFOLEVEL_REG[0] ;
 wire \TXFIFOLEVEL_REG[1] ;
 wire \TXFIFOLEVEL_REG[2] ;
 wire \TXFIFOLEVEL_REG[3] ;
 wire net56;
 wire net57;
 wire net58;
 wire eco_net;
 wire eco_net_0;
 wire eco_net_10_0;
 wire eco_net_11_0;
 wire eco_net_12_0;
 wire eco_net_13_0;
 wire eco_net_14_0;
 wire eco_net_15_0;
 wire eco_net_16_0;
 wire eco_net_17_0;
 wire eco_net_18_0;
 wire eco_net_19_0;
 wire eco_net_1_0;
 wire eco_net_20_0;
 wire eco_net_21_0;
 wire eco_net_22_0;
 wire eco_net_23_0;
 wire eco_net_24_0;
 wire eco_net_25_0;
 wire eco_net_26_0;
 wire eco_net_27_0;
 wire eco_net_28_0;
 wire eco_net_29_0;
 wire eco_net_2_0;
 wire eco_net_30_0;
 wire eco_net_3_0;
 wire eco_net_4_0;
 wire eco_net_5_0;
 wire eco_net_6_0;
 wire eco_net_7_0;
 wire eco_net_8_0;
 wire eco_net_9_0;
 wire \inst_to_wrap_out_data_o[0] ;
 wire \inst_to_wrap_out_data_o[1] ;
 wire \inst_to_wrap_out_data_o[2] ;
 wire \inst_to_wrap_out_data_o[3] ;
 wire \inst_to_wrap_out_data_o[4] ;
 wire \inst_to_wrap_out_data_o[5] ;
 wire \inst_to_wrap_out_data_o[6] ;
 wire \inst_to_wrap_out_data_o[7] ;
 wire \inst_to_wrap_rx_fifo_array_reg[0] ;
 wire \inst_to_wrap_rx_fifo_array_reg[100] ;
 wire \inst_to_wrap_rx_fifo_array_reg[101] ;
 wire \inst_to_wrap_rx_fifo_array_reg[102] ;
 wire \inst_to_wrap_rx_fifo_array_reg[103] ;
 wire \inst_to_wrap_rx_fifo_array_reg[104] ;
 wire \inst_to_wrap_rx_fifo_array_reg[105] ;
 wire \inst_to_wrap_rx_fifo_array_reg[106] ;
 wire \inst_to_wrap_rx_fifo_array_reg[107] ;
 wire \inst_to_wrap_rx_fifo_array_reg[108] ;
 wire \inst_to_wrap_rx_fifo_array_reg[109] ;
 wire \inst_to_wrap_rx_fifo_array_reg[10] ;
 wire \inst_to_wrap_rx_fifo_array_reg[110] ;
 wire \inst_to_wrap_rx_fifo_array_reg[111] ;
 wire \inst_to_wrap_rx_fifo_array_reg[112] ;
 wire \inst_to_wrap_rx_fifo_array_reg[113] ;
 wire \inst_to_wrap_rx_fifo_array_reg[114] ;
 wire \inst_to_wrap_rx_fifo_array_reg[115] ;
 wire \inst_to_wrap_rx_fifo_array_reg[116] ;
 wire \inst_to_wrap_rx_fifo_array_reg[117] ;
 wire \inst_to_wrap_rx_fifo_array_reg[118] ;
 wire \inst_to_wrap_rx_fifo_array_reg[119] ;
 wire \inst_to_wrap_rx_fifo_array_reg[11] ;
 wire \inst_to_wrap_rx_fifo_array_reg[120] ;
 wire \inst_to_wrap_rx_fifo_array_reg[121] ;
 wire \inst_to_wrap_rx_fifo_array_reg[122] ;
 wire \inst_to_wrap_rx_fifo_array_reg[123] ;
 wire \inst_to_wrap_rx_fifo_array_reg[124] ;
 wire \inst_to_wrap_rx_fifo_array_reg[125] ;
 wire \inst_to_wrap_rx_fifo_array_reg[126] ;
 wire \inst_to_wrap_rx_fifo_array_reg[127] ;
 wire \inst_to_wrap_rx_fifo_array_reg[12] ;
 wire \inst_to_wrap_rx_fifo_array_reg[13] ;
 wire \inst_to_wrap_rx_fifo_array_reg[14] ;
 wire \inst_to_wrap_rx_fifo_array_reg[15] ;
 wire \inst_to_wrap_rx_fifo_array_reg[16] ;
 wire \inst_to_wrap_rx_fifo_array_reg[17] ;
 wire \inst_to_wrap_rx_fifo_array_reg[18] ;
 wire \inst_to_wrap_rx_fifo_array_reg[19] ;
 wire \inst_to_wrap_rx_fifo_array_reg[1] ;
 wire \inst_to_wrap_rx_fifo_array_reg[20] ;
 wire \inst_to_wrap_rx_fifo_array_reg[21] ;
 wire \inst_to_wrap_rx_fifo_array_reg[22] ;
 wire \inst_to_wrap_rx_fifo_array_reg[23] ;
 wire \inst_to_wrap_rx_fifo_array_reg[24] ;
 wire \inst_to_wrap_rx_fifo_array_reg[25] ;
 wire \inst_to_wrap_rx_fifo_array_reg[26] ;
 wire \inst_to_wrap_rx_fifo_array_reg[27] ;
 wire \inst_to_wrap_rx_fifo_array_reg[28] ;
 wire \inst_to_wrap_rx_fifo_array_reg[29] ;
 wire \inst_to_wrap_rx_fifo_array_reg[2] ;
 wire \inst_to_wrap_rx_fifo_array_reg[30] ;
 wire \inst_to_wrap_rx_fifo_array_reg[31] ;
 wire \inst_to_wrap_rx_fifo_array_reg[32] ;
 wire \inst_to_wrap_rx_fifo_array_reg[33] ;
 wire \inst_to_wrap_rx_fifo_array_reg[34] ;
 wire \inst_to_wrap_rx_fifo_array_reg[35] ;
 wire \inst_to_wrap_rx_fifo_array_reg[36] ;
 wire \inst_to_wrap_rx_fifo_array_reg[37] ;
 wire \inst_to_wrap_rx_fifo_array_reg[38] ;
 wire \inst_to_wrap_rx_fifo_array_reg[39] ;
 wire \inst_to_wrap_rx_fifo_array_reg[3] ;
 wire \inst_to_wrap_rx_fifo_array_reg[40] ;
 wire \inst_to_wrap_rx_fifo_array_reg[41] ;
 wire \inst_to_wrap_rx_fifo_array_reg[42] ;
 wire \inst_to_wrap_rx_fifo_array_reg[43] ;
 wire \inst_to_wrap_rx_fifo_array_reg[44] ;
 wire \inst_to_wrap_rx_fifo_array_reg[45] ;
 wire \inst_to_wrap_rx_fifo_array_reg[46] ;
 wire \inst_to_wrap_rx_fifo_array_reg[47] ;
 wire \inst_to_wrap_rx_fifo_array_reg[48] ;
 wire \inst_to_wrap_rx_fifo_array_reg[49] ;
 wire \inst_to_wrap_rx_fifo_array_reg[4] ;
 wire \inst_to_wrap_rx_fifo_array_reg[50] ;
 wire \inst_to_wrap_rx_fifo_array_reg[51] ;
 wire \inst_to_wrap_rx_fifo_array_reg[52] ;
 wire \inst_to_wrap_rx_fifo_array_reg[53] ;
 wire \inst_to_wrap_rx_fifo_array_reg[54] ;
 wire \inst_to_wrap_rx_fifo_array_reg[55] ;
 wire \inst_to_wrap_rx_fifo_array_reg[56] ;
 wire \inst_to_wrap_rx_fifo_array_reg[57] ;
 wire \inst_to_wrap_rx_fifo_array_reg[58] ;
 wire \inst_to_wrap_rx_fifo_array_reg[59] ;
 wire \inst_to_wrap_rx_fifo_array_reg[5] ;
 wire \inst_to_wrap_rx_fifo_array_reg[60] ;
 wire \inst_to_wrap_rx_fifo_array_reg[61] ;
 wire \inst_to_wrap_rx_fifo_array_reg[62] ;
 wire \inst_to_wrap_rx_fifo_array_reg[63] ;
 wire \inst_to_wrap_rx_fifo_array_reg[64] ;
 wire \inst_to_wrap_rx_fifo_array_reg[65] ;
 wire \inst_to_wrap_rx_fifo_array_reg[66] ;
 wire \inst_to_wrap_rx_fifo_array_reg[67] ;
 wire \inst_to_wrap_rx_fifo_array_reg[68] ;
 wire \inst_to_wrap_rx_fifo_array_reg[69] ;
 wire \inst_to_wrap_rx_fifo_array_reg[6] ;
 wire \inst_to_wrap_rx_fifo_array_reg[70] ;
 wire \inst_to_wrap_rx_fifo_array_reg[71] ;
 wire \inst_to_wrap_rx_fifo_array_reg[72] ;
 wire \inst_to_wrap_rx_fifo_array_reg[73] ;
 wire \inst_to_wrap_rx_fifo_array_reg[74] ;
 wire \inst_to_wrap_rx_fifo_array_reg[75] ;
 wire \inst_to_wrap_rx_fifo_array_reg[76] ;
 wire \inst_to_wrap_rx_fifo_array_reg[77] ;
 wire \inst_to_wrap_rx_fifo_array_reg[78] ;
 wire \inst_to_wrap_rx_fifo_array_reg[79] ;
 wire \inst_to_wrap_rx_fifo_array_reg[7] ;
 wire \inst_to_wrap_rx_fifo_array_reg[80] ;
 wire \inst_to_wrap_rx_fifo_array_reg[81] ;
 wire \inst_to_wrap_rx_fifo_array_reg[82] ;
 wire \inst_to_wrap_rx_fifo_array_reg[83] ;
 wire \inst_to_wrap_rx_fifo_array_reg[84] ;
 wire \inst_to_wrap_rx_fifo_array_reg[85] ;
 wire \inst_to_wrap_rx_fifo_array_reg[86] ;
 wire \inst_to_wrap_rx_fifo_array_reg[87] ;
 wire \inst_to_wrap_rx_fifo_array_reg[88] ;
 wire \inst_to_wrap_rx_fifo_array_reg[89] ;
 wire \inst_to_wrap_rx_fifo_array_reg[8] ;
 wire \inst_to_wrap_rx_fifo_array_reg[90] ;
 wire \inst_to_wrap_rx_fifo_array_reg[91] ;
 wire \inst_to_wrap_rx_fifo_array_reg[92] ;
 wire \inst_to_wrap_rx_fifo_array_reg[93] ;
 wire \inst_to_wrap_rx_fifo_array_reg[94] ;
 wire \inst_to_wrap_rx_fifo_array_reg[95] ;
 wire \inst_to_wrap_rx_fifo_array_reg[96] ;
 wire \inst_to_wrap_rx_fifo_array_reg[97] ;
 wire \inst_to_wrap_rx_fifo_array_reg[98] ;
 wire \inst_to_wrap_rx_fifo_array_reg[99] ;
 wire \inst_to_wrap_rx_fifo_array_reg[9] ;
 wire \inst_to_wrap_rx_fifo_r_ptr_reg[0] ;
 wire \inst_to_wrap_rx_fifo_r_ptr_reg[1] ;
 wire \inst_to_wrap_rx_fifo_r_ptr_reg[2] ;
 wire \inst_to_wrap_rx_fifo_r_ptr_reg[3] ;
 wire \inst_to_wrap_rx_fifo_w_ptr_reg[0] ;
 wire \inst_to_wrap_rx_fifo_w_ptr_reg[1] ;
 wire \inst_to_wrap_rx_fifo_w_ptr_reg[2] ;
 wire \inst_to_wrap_rx_fifo_w_ptr_reg[3] ;
 wire \inst_to_wrap_tx_fifo_array_reg[0] ;
 wire \inst_to_wrap_tx_fifo_array_reg[100] ;
 wire \inst_to_wrap_tx_fifo_array_reg[101] ;
 wire \inst_to_wrap_tx_fifo_array_reg[102] ;
 wire \inst_to_wrap_tx_fifo_array_reg[103] ;
 wire \inst_to_wrap_tx_fifo_array_reg[104] ;
 wire \inst_to_wrap_tx_fifo_array_reg[105] ;
 wire \inst_to_wrap_tx_fifo_array_reg[106] ;
 wire \inst_to_wrap_tx_fifo_array_reg[107] ;
 wire \inst_to_wrap_tx_fifo_array_reg[108] ;
 wire \inst_to_wrap_tx_fifo_array_reg[109] ;
 wire \inst_to_wrap_tx_fifo_array_reg[10] ;
 wire \inst_to_wrap_tx_fifo_array_reg[110] ;
 wire \inst_to_wrap_tx_fifo_array_reg[111] ;
 wire \inst_to_wrap_tx_fifo_array_reg[112] ;
 wire \inst_to_wrap_tx_fifo_array_reg[113] ;
 wire \inst_to_wrap_tx_fifo_array_reg[114] ;
 wire \inst_to_wrap_tx_fifo_array_reg[115] ;
 wire \inst_to_wrap_tx_fifo_array_reg[116] ;
 wire \inst_to_wrap_tx_fifo_array_reg[117] ;
 wire \inst_to_wrap_tx_fifo_array_reg[118] ;
 wire \inst_to_wrap_tx_fifo_array_reg[119] ;
 wire \inst_to_wrap_tx_fifo_array_reg[11] ;
 wire \inst_to_wrap_tx_fifo_array_reg[120] ;
 wire \inst_to_wrap_tx_fifo_array_reg[121] ;
 wire \inst_to_wrap_tx_fifo_array_reg[122] ;
 wire \inst_to_wrap_tx_fifo_array_reg[123] ;
 wire \inst_to_wrap_tx_fifo_array_reg[124] ;
 wire \inst_to_wrap_tx_fifo_array_reg[125] ;
 wire \inst_to_wrap_tx_fifo_array_reg[126] ;
 wire \inst_to_wrap_tx_fifo_array_reg[127] ;
 wire \inst_to_wrap_tx_fifo_array_reg[12] ;
 wire \inst_to_wrap_tx_fifo_array_reg[13] ;
 wire \inst_to_wrap_tx_fifo_array_reg[14] ;
 wire \inst_to_wrap_tx_fifo_array_reg[15] ;
 wire \inst_to_wrap_tx_fifo_array_reg[16] ;
 wire \inst_to_wrap_tx_fifo_array_reg[17] ;
 wire \inst_to_wrap_tx_fifo_array_reg[18] ;
 wire \inst_to_wrap_tx_fifo_array_reg[19] ;
 wire \inst_to_wrap_tx_fifo_array_reg[1] ;
 wire \inst_to_wrap_tx_fifo_array_reg[20] ;
 wire \inst_to_wrap_tx_fifo_array_reg[21] ;
 wire \inst_to_wrap_tx_fifo_array_reg[22] ;
 wire \inst_to_wrap_tx_fifo_array_reg[23] ;
 wire \inst_to_wrap_tx_fifo_array_reg[24] ;
 wire \inst_to_wrap_tx_fifo_array_reg[25] ;
 wire \inst_to_wrap_tx_fifo_array_reg[26] ;
 wire \inst_to_wrap_tx_fifo_array_reg[27] ;
 wire \inst_to_wrap_tx_fifo_array_reg[28] ;
 wire \inst_to_wrap_tx_fifo_array_reg[29] ;
 wire \inst_to_wrap_tx_fifo_array_reg[2] ;
 wire \inst_to_wrap_tx_fifo_array_reg[30] ;
 wire \inst_to_wrap_tx_fifo_array_reg[31] ;
 wire \inst_to_wrap_tx_fifo_array_reg[32] ;
 wire \inst_to_wrap_tx_fifo_array_reg[33] ;
 wire \inst_to_wrap_tx_fifo_array_reg[34] ;
 wire \inst_to_wrap_tx_fifo_array_reg[35] ;
 wire \inst_to_wrap_tx_fifo_array_reg[36] ;
 wire \inst_to_wrap_tx_fifo_array_reg[37] ;
 wire \inst_to_wrap_tx_fifo_array_reg[38] ;
 wire \inst_to_wrap_tx_fifo_array_reg[39] ;
 wire \inst_to_wrap_tx_fifo_array_reg[3] ;
 wire \inst_to_wrap_tx_fifo_array_reg[40] ;
 wire \inst_to_wrap_tx_fifo_array_reg[41] ;
 wire \inst_to_wrap_tx_fifo_array_reg[42] ;
 wire \inst_to_wrap_tx_fifo_array_reg[43] ;
 wire \inst_to_wrap_tx_fifo_array_reg[44] ;
 wire \inst_to_wrap_tx_fifo_array_reg[45] ;
 wire \inst_to_wrap_tx_fifo_array_reg[46] ;
 wire \inst_to_wrap_tx_fifo_array_reg[47] ;
 wire \inst_to_wrap_tx_fifo_array_reg[48] ;
 wire \inst_to_wrap_tx_fifo_array_reg[49] ;
 wire \inst_to_wrap_tx_fifo_array_reg[4] ;
 wire \inst_to_wrap_tx_fifo_array_reg[50] ;
 wire \inst_to_wrap_tx_fifo_array_reg[51] ;
 wire \inst_to_wrap_tx_fifo_array_reg[52] ;
 wire \inst_to_wrap_tx_fifo_array_reg[53] ;
 wire \inst_to_wrap_tx_fifo_array_reg[54] ;
 wire \inst_to_wrap_tx_fifo_array_reg[55] ;
 wire \inst_to_wrap_tx_fifo_array_reg[56] ;
 wire \inst_to_wrap_tx_fifo_array_reg[57] ;
 wire \inst_to_wrap_tx_fifo_array_reg[58] ;
 wire \inst_to_wrap_tx_fifo_array_reg[59] ;
 wire \inst_to_wrap_tx_fifo_array_reg[5] ;
 wire \inst_to_wrap_tx_fifo_array_reg[60] ;
 wire \inst_to_wrap_tx_fifo_array_reg[61] ;
 wire \inst_to_wrap_tx_fifo_array_reg[62] ;
 wire \inst_to_wrap_tx_fifo_array_reg[63] ;
 wire \inst_to_wrap_tx_fifo_array_reg[64] ;
 wire \inst_to_wrap_tx_fifo_array_reg[65] ;
 wire \inst_to_wrap_tx_fifo_array_reg[66] ;
 wire \inst_to_wrap_tx_fifo_array_reg[67] ;
 wire \inst_to_wrap_tx_fifo_array_reg[68] ;
 wire \inst_to_wrap_tx_fifo_array_reg[69] ;
 wire \inst_to_wrap_tx_fifo_array_reg[6] ;
 wire \inst_to_wrap_tx_fifo_array_reg[70] ;
 wire \inst_to_wrap_tx_fifo_array_reg[71] ;
 wire \inst_to_wrap_tx_fifo_array_reg[72] ;
 wire \inst_to_wrap_tx_fifo_array_reg[73] ;
 wire \inst_to_wrap_tx_fifo_array_reg[74] ;
 wire \inst_to_wrap_tx_fifo_array_reg[75] ;
 wire \inst_to_wrap_tx_fifo_array_reg[76] ;
 wire \inst_to_wrap_tx_fifo_array_reg[77] ;
 wire \inst_to_wrap_tx_fifo_array_reg[78] ;
 wire \inst_to_wrap_tx_fifo_array_reg[79] ;
 wire \inst_to_wrap_tx_fifo_array_reg[7] ;
 wire \inst_to_wrap_tx_fifo_array_reg[80] ;
 wire \inst_to_wrap_tx_fifo_array_reg[81] ;
 wire \inst_to_wrap_tx_fifo_array_reg[82] ;
 wire \inst_to_wrap_tx_fifo_array_reg[83] ;
 wire \inst_to_wrap_tx_fifo_array_reg[84] ;
 wire \inst_to_wrap_tx_fifo_array_reg[85] ;
 wire \inst_to_wrap_tx_fifo_array_reg[86] ;
 wire \inst_to_wrap_tx_fifo_array_reg[87] ;
 wire \inst_to_wrap_tx_fifo_array_reg[88] ;
 wire \inst_to_wrap_tx_fifo_array_reg[89] ;
 wire \inst_to_wrap_tx_fifo_array_reg[8] ;
 wire \inst_to_wrap_tx_fifo_array_reg[90] ;
 wire \inst_to_wrap_tx_fifo_array_reg[91] ;
 wire \inst_to_wrap_tx_fifo_array_reg[92] ;
 wire \inst_to_wrap_tx_fifo_array_reg[93] ;
 wire \inst_to_wrap_tx_fifo_array_reg[94] ;
 wire \inst_to_wrap_tx_fifo_array_reg[95] ;
 wire \inst_to_wrap_tx_fifo_array_reg[96] ;
 wire \inst_to_wrap_tx_fifo_array_reg[97] ;
 wire \inst_to_wrap_tx_fifo_array_reg[98] ;
 wire \inst_to_wrap_tx_fifo_array_reg[99] ;
 wire \inst_to_wrap_tx_fifo_array_reg[9] ;
 wire \inst_to_wrap_tx_fifo_r_ptr_reg[0] ;
 wire \inst_to_wrap_tx_fifo_r_ptr_reg[1] ;
 wire \inst_to_wrap_tx_fifo_r_ptr_reg[2] ;
 wire \inst_to_wrap_tx_fifo_r_ptr_reg[3] ;
 wire \inst_to_wrap_tx_fifo_w_ptr_reg[0] ;
 wire \inst_to_wrap_tx_fifo_w_ptr_reg[1] ;
 wire \inst_to_wrap_tx_fifo_w_ptr_reg[2] ;
 wire \inst_to_wrap_tx_fifo_w_ptr_reg[3] ;
 wire \inst_to_wrap_u_usb_cdc_addr[0] ;
 wire \inst_to_wrap_u_usb_cdc_addr[1] ;
 wire \inst_to_wrap_u_usb_cdc_addr[2] ;
 wire \inst_to_wrap_u_usb_cdc_addr[3] ;
 wire \inst_to_wrap_u_usb_cdc_addr[4] ;
 wire \inst_to_wrap_u_usb_cdc_addr[5] ;
 wire \inst_to_wrap_u_usb_cdc_addr[6] ;
 wire inst_to_wrap_u_usb_cdc_bulk_in_valid;
 wire inst_to_wrap_u_usb_cdc_bulk_out_nak;
 wire inst_to_wrap_u_usb_cdc_ctrl_in_req;
 wire \inst_to_wrap_u_usb_cdc_endp[0] ;
 wire \inst_to_wrap_u_usb_cdc_endp[1] ;
 wire \inst_to_wrap_u_usb_cdc_endp[2] ;
 wire \inst_to_wrap_u_usb_cdc_endp[3] ;
 wire inst_to_wrap_u_usb_cdc_in_data_ack;
 wire \inst_to_wrap_u_usb_cdc_out_data[0] ;
 wire \inst_to_wrap_u_usb_cdc_out_data[1] ;
 wire \inst_to_wrap_u_usb_cdc_out_data[2] ;
 wire \inst_to_wrap_u_usb_cdc_out_data[3] ;
 wire \inst_to_wrap_u_usb_cdc_out_data[4] ;
 wire \inst_to_wrap_u_usb_cdc_out_data[5] ;
 wire \inst_to_wrap_u_usb_cdc_out_data[6] ;
 wire \inst_to_wrap_u_usb_cdc_out_data[7] ;
 wire inst_to_wrap_u_usb_cdc_out_err;
 wire \inst_to_wrap_u_usb_cdc_rstn_sq[0] ;
 wire \inst_to_wrap_u_usb_cdc_rstn_sq[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[10] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[11] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[12] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[13] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[14] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[15] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[16] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[17] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[18] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[19] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[20] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[21] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[22] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[23] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[24] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[25] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[26] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[27] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[28] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[29] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[30] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[31] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[32] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[33] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[34] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[35] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[36] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[37] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[38] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[39] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[40] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[41] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[42] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[43] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[44] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[45] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[46] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[47] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[48] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[49] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[50] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[51] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[52] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[53] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[54] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[55] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[56] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[57] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[58] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[59] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[60] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[61] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[62] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[63] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[64] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[65] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[66] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[67] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[68] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[69] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[70] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[71] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[7] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[8] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[9] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[3] ;
 wire inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q;
 wire inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_state_q;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[7] ;
 wire inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_mask_q;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq[1] ;
 wire inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_mask_q;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[10] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[11] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[12] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[13] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[14] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[15] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[16] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[17] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[18] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[19] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[20] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[21] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[22] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[23] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[24] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[25] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[26] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[27] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[28] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[29] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[30] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[31] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[32] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[33] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[34] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[35] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[36] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[37] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[38] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[39] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[40] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[41] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[42] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[43] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[44] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[45] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[46] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[47] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[48] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[49] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[50] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[51] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[52] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[53] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[54] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[55] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[56] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[57] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[58] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[59] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[60] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[61] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[62] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[63] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[64] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[65] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[66] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[67] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[68] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[69] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[70] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[71] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[7] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[8] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[9] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ;
 wire inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_full_o;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[1] ;
 wire inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_mask_q;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq[1] ;
 wire inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_mask_q;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq[1] ;
 wire inst_to_wrap_u_usb_cdc_u_ctrl_endp_N109;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ;
 wire inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ;
 wire inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q;
 wire inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_endp_q;
 wire inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[1] ;
 wire inst_to_wrap_u_usb_cdc_u_ctrl_endp_usb_reset_q;
 wire \inst_to_wrap_u_usb_cdc_u_sie_addr_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_addr_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_addr_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_addr_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_addr_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_addr_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_addr_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[10] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[11] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[12] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[13] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[14] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[15] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[7] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[8] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_crc16_q[9] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[3] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_out_eop_q;
 wire \inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_pid_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_pid_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_pid_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_N51;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[10] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[11] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[12] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[13] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[14] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[15] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[16] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[17] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[7] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[8] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[9] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_0_;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_fq;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[2] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_N30;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_N31;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[3] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[4] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[5] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[6] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[7] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[1] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[2] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ;
 wire \inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[1] ;
 wire inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q;
 wire net59;
 wire \last_HADDR[0] ;
 wire \last_HADDR[10] ;
 wire \last_HADDR[11] ;
 wire \last_HADDR[12] ;
 wire \last_HADDR[13] ;
 wire \last_HADDR[14] ;
 wire \last_HADDR[15] ;
 wire \last_HADDR[1] ;
 wire \last_HADDR[2] ;
 wire \last_HADDR[3] ;
 wire \last_HADDR[4] ;
 wire \last_HADDR[5] ;
 wire \last_HADDR[6] ;
 wire \last_HADDR[7] ;
 wire \last_HADDR[8] ;
 wire \last_HADDR[9] ;
 wire last_HSEL;
 wire last_HTRANS_1_;
 wire last_HWRITE;
 wire n1576;
 wire n1577;
 wire n1578;
 wire n1580;
 wire n1581;
 wire n1582;
 wire n1583;
 wire n1584;
 wire n1585;
 wire n1586;
 wire n1587;
 wire n1588;
 wire n1589;
 wire n1590;
 wire n1591;
 wire n1592;
 wire n1593;
 wire n1594;
 wire n1595;
 wire n1596;
 wire n1597;
 wire n1598;
 wire n1599;
 wire n1600;
 wire n1601;
 wire n1602;
 wire n1603;
 wire n1604;
 wire n1605;
 wire n1606;
 wire n1607;
 wire n1608;
 wire n1609;
 wire n1610;
 wire n1611;
 wire n1612;
 wire n1613;
 wire n1614;
 wire n1615;
 wire n1616;
 wire n1617;
 wire n1618;
 wire n1619;
 wire n1620;
 wire n1621;
 wire n1622;
 wire n1623;
 wire n1624;
 wire n1625;
 wire n1626;
 wire n1627;
 wire n1628;
 wire n1629;
 wire n1630;
 wire n1631;
 wire n1632;
 wire n1633;
 wire n1634;
 wire n1635;
 wire n1636;
 wire n1637;
 wire n1638;
 wire n1639;
 wire n1640;
 wire n1641;
 wire n1642;
 wire n1643;
 wire n1644;
 wire n1645;
 wire n1646;
 wire n1647;
 wire n1648;
 wire n1649;
 wire n1650;
 wire n1651;
 wire n1652;
 wire n1653;
 wire n1654;
 wire n1655;
 wire n1656;
 wire n1657;
 wire n1658;
 wire n1659;
 wire n1660;
 wire n1661;
 wire n1662;
 wire n1663;
 wire n1664;
 wire n1665;
 wire n1666;
 wire n1667;
 wire n1668;
 wire n1669;
 wire n1670;
 wire n1671;
 wire n1672;
 wire n1673;
 wire n1674;
 wire n1675;
 wire n1676;
 wire n1677;
 wire n1678;
 wire n1679;
 wire n1680;
 wire n1681;
 wire n1682;
 wire n1683;
 wire n1684;
 wire n1685;
 wire n1686;
 wire n1687;
 wire n1688;
 wire n1689;
 wire n1690;
 wire n1691;
 wire n1692;
 wire n1693;
 wire n1694;
 wire n1695;
 wire n1696;
 wire n1697;
 wire n1698;
 wire n1699;
 wire n1700;
 wire n1701;
 wire n1702;
 wire n1703;
 wire n1704;
 wire n1705;
 wire n1706;
 wire n1707;
 wire n1708;
 wire n1709;
 wire n1710;
 wire n1711;
 wire n1712;
 wire n1713;
 wire n1714;
 wire n1715;
 wire n1716;
 wire n1717;
 wire n1718;
 wire n1719;
 wire n1720;
 wire n1721;
 wire n1722;
 wire n1723;
 wire n1724;
 wire n1725;
 wire n1726;
 wire n1727;
 wire n1728;
 wire n1729;
 wire n1730;
 wire n1731;
 wire n1732;
 wire n1733;
 wire n1734;
 wire n1735;
 wire n1736;
 wire n1737;
 wire n1738;
 wire n1739;
 wire n1740;
 wire n1741;
 wire n1742;
 wire n1743;
 wire n1744;
 wire n1745;
 wire n1746;
 wire n1747;
 wire n1748;
 wire n1749;
 wire n1750;
 wire n1751;
 wire n1752;
 wire n1753;
 wire n1754;
 wire n1755;
 wire n1756;
 wire n1757;
 wire n1758;
 wire n1759;
 wire n1760;
 wire n1761;
 wire n1762;
 wire n1763;
 wire n1764;
 wire n1765;
 wire n1766;
 wire n1767;
 wire n1768;
 wire n1769;
 wire n1770;
 wire n1771;
 wire n1772;
 wire n1773;
 wire n1774;
 wire n1775;
 wire n1776;
 wire n1777;
 wire n1778;
 wire n1779;
 wire n1780;
 wire n1781;
 wire n1782;
 wire n1783;
 wire n1784;
 wire n1785;
 wire n1786;
 wire n1787;
 wire n1788;
 wire n1789;
 wire n1790;
 wire n1791;
 wire n1792;
 wire n1793;
 wire n1794;
 wire n1795;
 wire n1796;
 wire n1797;
 wire n1798;
 wire n1799;
 wire n1800;
 wire n1801;
 wire n1802;
 wire n1803;
 wire n1804;
 wire n1805;
 wire n1806;
 wire n1807;
 wire n1808;
 wire n1809;
 wire n1810;
 wire n1811;
 wire n1812;
 wire n1813;
 wire n1814;
 wire n1815;
 wire n1816;
 wire n1817;
 wire n1818;
 wire n1819;
 wire n1820;
 wire n1821;
 wire n1822;
 wire n1823;
 wire n1824;
 wire n1825;
 wire n1826;
 wire n1827;
 wire n1828;
 wire n1829;
 wire n1830;
 wire n1831;
 wire n1832;
 wire n1833;
 wire n1834;
 wire n1835;
 wire n1836;
 wire n1837;
 wire n1838;
 wire n1839;
 wire n1840;
 wire n1841;
 wire n1842;
 wire n1843;
 wire n1844;
 wire n1845;
 wire n1846;
 wire n1847;
 wire n1848;
 wire n1849;
 wire n1850;
 wire n1851;
 wire n1852;
 wire n1853;
 wire n1854;
 wire n1855;
 wire n1856;
 wire n1857;
 wire n1858;
 wire n1859;
 wire n1860;
 wire n1861;
 wire n1862;
 wire n1863;
 wire n1864;
 wire n1865;
 wire n1866;
 wire n1867;
 wire n1868;
 wire n1869;
 wire n1870;
 wire n1871;
 wire n1872;
 wire n1873;
 wire n1874;
 wire n1875;
 wire n1876;
 wire n1877;
 wire n1878;
 wire n1879;
 wire n1880;
 wire n1881;
 wire n1882;
 wire n1883;
 wire n1884;
 wire n1885;
 wire n1886;
 wire n1887;
 wire n1888;
 wire n1889;
 wire n1890;
 wire n1891;
 wire n1892;
 wire n1893;
 wire n1894;
 wire n1895;
 wire n1896;
 wire n1897;
 wire n1898;
 wire n1899;
 wire n1900;
 wire n1901;
 wire n1902;
 wire n1903;
 wire n1904;
 wire n1905;
 wire n1906;
 wire n1907;
 wire n1908;
 wire n1909;
 wire n1910;
 wire n1911;
 wire n1912;
 wire n1913;
 wire n1914;
 wire n1915;
 wire n1916;
 wire n1917;
 wire n1918;
 wire n1919;
 wire n1920;
 wire n1921;
 wire n1922;
 wire n1923;
 wire n1924;
 wire n1925;
 wire n1926;
 wire n1927;
 wire n1928;
 wire n1929;
 wire n1930;
 wire n1931;
 wire n1932;
 wire n1933;
 wire n1934;
 wire n1935;
 wire n1936;
 wire n1937;
 wire n1938;
 wire n1939;
 wire n1940;
 wire n1941;
 wire n1942;
 wire n1943;
 wire n1944;
 wire n1945;
 wire n1946;
 wire n1947;
 wire n1948;
 wire n1949;
 wire n1950;
 wire n1951;
 wire n1952;
 wire n1953;
 wire n1954;
 wire n1955;
 wire n1956;
 wire n1957;
 wire n1958;
 wire n1959;
 wire n1960;
 wire n1961;
 wire n1962;
 wire n1963;
 wire n1964;
 wire n1965;
 wire n1966;
 wire n1967;
 wire n1968;
 wire n1969;
 wire n1970;
 wire n1971;
 wire n1972;
 wire n1973;
 wire n1974;
 wire n1975;
 wire n1976;
 wire n1977;
 wire n1978;
 wire n1979;
 wire n1980;
 wire n1981;
 wire n1982;
 wire n1983;
 wire n1984;
 wire n1985;
 wire n1986;
 wire n1987;
 wire n1988;
 wire n1989;
 wire n1990;
 wire n1991;
 wire n1992;
 wire n1993;
 wire n1994;
 wire n1995;
 wire n1996;
 wire n1997;
 wire n1998;
 wire n1999;
 wire n2000;
 wire n2001;
 wire n2002;
 wire n2003;
 wire n2004;
 wire n2005;
 wire n2006;
 wire n2007;
 wire n2008;
 wire n2009;
 wire n2010;
 wire n2011;
 wire n2012;
 wire n2013;
 wire n2014;
 wire n2015;
 wire n2016;
 wire n2017;
 wire n2018;
 wire n2019;
 wire n2020;
 wire n2021;
 wire n2022;
 wire n2023;
 wire n2024;
 wire n2025;
 wire n2026;
 wire n2027;
 wire n2028;
 wire n2029;
 wire n2030;
 wire n2031;
 wire n2032;
 wire n2033;
 wire n2034;
 wire n2035;
 wire n2036;
 wire n2037;
 wire n2038;
 wire n2039;
 wire n2040;
 wire n2041;
 wire n2042;
 wire n2043;
 wire n2044;
 wire n2045;
 wire n2046;
 wire n2047;
 wire n2048;
 wire n2049;
 wire n2050;
 wire n2051;
 wire n2052;
 wire n2053;
 wire n2054;
 wire n2055;
 wire n2056;
 wire n2057;
 wire n2058;
 wire n2059;
 wire n2060;
 wire n2061;
 wire n2062;
 wire n2063;
 wire n2064;
 wire n2065;
 wire n2066;
 wire n2067;
 wire n2068;
 wire n2069;
 wire n2070;
 wire n2071;
 wire n2072;
 wire n2073;
 wire n2074;
 wire n2075;
 wire n2076;
 wire n2077;
 wire n2078;
 wire n2079;
 wire n2080;
 wire n2081;
 wire n2082;
 wire n2083;
 wire n2084;
 wire n2085;
 wire n2086;
 wire n2087;
 wire n2088;
 wire n2089;
 wire n2090;
 wire n2091;
 wire n2092;
 wire n2093;
 wire n2094;
 wire n2095;
 wire n2096;
 wire n2097;
 wire n2098;
 wire n2099;
 wire n2100;
 wire n2101;
 wire n2102;
 wire n2103;
 wire n2104;
 wire n2105;
 wire n2106;
 wire n2107;
 wire n2108;
 wire n2109;
 wire n2110;
 wire n2111;
 wire n2112;
 wire n2113;
 wire n2114;
 wire n2115;
 wire n2116;
 wire n2117;
 wire n2118;
 wire n2119;
 wire n2120;
 wire n2121;
 wire n2122;
 wire n2123;
 wire n2124;
 wire n2125;
 wire n2126;
 wire n2127;
 wire n2128;
 wire n2129;
 wire n2130;
 wire n2131;
 wire n2132;
 wire n2133;
 wire n2134;
 wire n2135;
 wire n2136;
 wire n2137;
 wire n2138;
 wire n2139;
 wire n2140;
 wire n2141;
 wire n2142;
 wire n2143;
 wire n2144;
 wire n2145;
 wire n2146;
 wire n2147;
 wire n2148;
 wire n2149;
 wire n2150;
 wire n2151;
 wire n2152;
 wire n2153;
 wire n2154;
 wire n2155;
 wire n2156;
 wire n2157;
 wire n2158;
 wire n2159;
 wire n2160;
 wire n2161;
 wire n2162;
 wire n2163;
 wire n2164;
 wire n2165;
 wire n2166;
 wire n2167;
 wire n2168;
 wire n2169;
 wire n2170;
 wire n2171;
 wire n2172;
 wire n2173;
 wire n2174;
 wire n2175;
 wire n2176;
 wire n2177;
 wire n2178;
 wire n2179;
 wire n2180;
 wire n2181;
 wire n2182;
 wire n2183;
 wire n2184;
 wire n2185;
 wire n2186;
 wire n2187;
 wire n2188;
 wire n2189;
 wire n2190;
 wire n2191;
 wire n2192;
 wire n2193;
 wire n2194;
 wire n2195;
 wire n2196;
 wire n2197;
 wire n2198;
 wire n2199;
 wire n2200;
 wire n2201;
 wire n2202;
 wire n2203;
 wire n2204;
 wire n2205;
 wire n2206;
 wire n2207;
 wire n2208;
 wire n2209;
 wire n2210;
 wire n2211;
 wire n2212;
 wire n2213;
 wire n2214;
 wire n2215;
 wire n2216;
 wire n2217;
 wire n2218;
 wire n2219;
 wire n2220;
 wire n2221;
 wire n2222;
 wire n2223;
 wire n2224;
 wire n2225;
 wire n2226;
 wire n2227;
 wire n2228;
 wire n2229;
 wire n2230;
 wire n2231;
 wire n2232;
 wire n2233;
 wire n2234;
 wire n2235;
 wire n2236;
 wire n2237;
 wire n2238;
 wire n2239;
 wire n2240;
 wire n2241;
 wire n2242;
 wire n2243;
 wire n2244;
 wire n2245;
 wire n2246;
 wire n2247;
 wire n2248;
 wire n2249;
 wire n2250;
 wire n2251;
 wire n2252;
 wire n2253;
 wire n2254;
 wire n2255;
 wire n2256;
 wire n2257;
 wire n2258;
 wire n2259;
 wire n2260;
 wire n2261;
 wire n2262;
 wire n2263;
 wire n2264;
 wire n2265;
 wire n2266;
 wire n2267;
 wire n2268;
 wire n2269;
 wire net62;
 wire clknet_leaf_0_HCLK;
 wire n2283;
 wire n2284;
 wire n2285;
 wire n2286;
 wire n2288;
 wire n2289;
 wire n2290;
 wire n2291;
 wire n2293;
 wire n2294;
 wire n2295;
 wire n2296;
 wire n2297;
 wire n2298;
 wire n2299;
 wire n2300;
 wire n2301;
 wire n2302;
 wire n2303;
 wire n2304;
 wire n2305;
 wire n2306;
 wire n2307;
 wire n2308;
 wire n2309;
 wire n2310;
 wire n2311;
 wire n2312;
 wire n2313;
 wire n2314;
 wire n2315;
 wire n2316;
 wire n2317;
 wire n2318;
 wire n2319;
 wire n2320;
 wire n2321;
 wire n2322;
 wire n2323;
 wire n2325;
 wire n2326;
 wire n2327;
 wire n2328;
 wire n2329;
 wire n2330;
 wire n2331;
 wire n2332;
 wire n2333;
 wire n2334;
 wire n2335;
 wire n2336;
 wire n2337;
 wire n2338;
 wire n2339;
 wire n2340;
 wire n2341;
 wire n2342;
 wire n2343;
 wire n2344;
 wire n2345;
 wire n2346;
 wire n2347;
 wire n2348;
 wire n2349;
 wire n2350;
 wire n2351;
 wire n2352;
 wire n2353;
 wire n2354;
 wire n2355;
 wire n2356;
 wire n2357;
 wire n2358;
 wire n2359;
 wire n2360;
 wire n2361;
 wire n2362;
 wire n2363;
 wire n2364;
 wire n2365;
 wire n2366;
 wire n2367;
 wire n2368;
 wire n2369;
 wire n2370;
 wire n2371;
 wire n2372;
 wire n2373;
 wire n2374;
 wire n2375;
 wire n2376;
 wire n2377;
 wire n2378;
 wire n2379;
 wire n2380;
 wire n2381;
 wire n2382;
 wire n2383;
 wire n2384;
 wire n2385;
 wire n2386;
 wire n2387;
 wire n2388;
 wire n2389;
 wire n2390;
 wire n2391;
 wire n2392;
 wire n2393;
 wire n2394;
 wire n2395;
 wire n2396;
 wire n2397;
 wire n2398;
 wire n2399;
 wire n2400;
 wire n2401;
 wire n2402;
 wire n2404;
 wire n2405;
 wire n2406;
 wire n2407;
 wire n2408;
 wire n2409;
 wire n2410;
 wire n2411;
 wire n2412;
 wire n2413;
 wire n2414;
 wire n2415;
 wire n2416;
 wire n2417;
 wire n2418;
 wire n2419;
 wire n2420;
 wire n2421;
 wire n2422;
 wire n2423;
 wire n2424;
 wire n2425;
 wire n2426;
 wire n2427;
 wire n2428;
 wire n2429;
 wire n2430;
 wire n2431;
 wire n2432;
 wire n2433;
 wire n2434;
 wire n2435;
 wire n2436;
 wire n2437;
 wire n2438;
 wire n2439;
 wire n2440;
 wire n2441;
 wire n2442;
 wire n2443;
 wire n2444;
 wire n2445;
 wire n2446;
 wire n2447;
 wire n2448;
 wire n2449;
 wire n2450;
 wire n2451;
 wire n2452;
 wire n2453;
 wire n2454;
 wire n2455;
 wire n2456;
 wire n2457;
 wire n2458;
 wire n2459;
 wire n2460;
 wire n2461;
 wire n2462;
 wire n2463;
 wire n2464;
 wire n2465;
 wire n2466;
 wire n2467;
 wire n2468;
 wire n2469;
 wire n2470;
 wire n2471;
 wire n2472;
 wire n2473;
 wire n2474;
 wire n2475;
 wire n2476;
 wire n2477;
 wire n2478;
 wire n2479;
 wire n2480;
 wire n2481;
 wire n2482;
 wire n2483;
 wire n2484;
 wire n2485;
 wire n2486;
 wire n2487;
 wire n2488;
 wire n2489;
 wire n2490;
 wire n2491;
 wire n2492;
 wire n2493;
 wire n2494;
 wire n2495;
 wire n2496;
 wire n2497;
 wire n2498;
 wire n2499;
 wire n2500;
 wire n2501;
 wire n2502;
 wire n2503;
 wire n2504;
 wire n2505;
 wire n2506;
 wire n2507;
 wire n2508;
 wire n2509;
 wire n2510;
 wire n2511;
 wire n2512;
 wire n2513;
 wire n2514;
 wire n2515;
 wire n2516;
 wire n2517;
 wire n2518;
 wire n2519;
 wire n2520;
 wire n2521;
 wire n2522;
 wire n2523;
 wire n2524;
 wire n2525;
 wire n2526;
 wire n2527;
 wire n2528;
 wire n2529;
 wire n2530;
 wire n2531;
 wire n2532;
 wire n2533;
 wire n2534;
 wire n2535;
 wire n2536;
 wire n2537;
 wire n2538;
 wire n2539;
 wire n2540;
 wire n2541;
 wire n2542;
 wire n2543;
 wire n2544;
 wire n2545;
 wire n2546;
 wire n2547;
 wire n2548;
 wire n2549;
 wire n2550;
 wire n2551;
 wire n2552;
 wire n2553;
 wire n2554;
 wire n2555;
 wire n2556;
 wire n2557;
 wire n2558;
 wire n2559;
 wire n2560;
 wire n2561;
 wire n2562;
 wire n2563;
 wire n2564;
 wire n2565;
 wire n2566;
 wire n2567;
 wire n2568;
 wire n2569;
 wire n2570;
 wire n2571;
 wire n2572;
 wire n2573;
 wire n2574;
 wire n2575;
 wire n2576;
 wire n2577;
 wire n2578;
 wire n2579;
 wire n2580;
 wire n2581;
 wire n2582;
 wire n2583;
 wire n2584;
 wire n2585;
 wire n2586;
 wire n2587;
 wire n2588;
 wire n2589;
 wire n2590;
 wire n2591;
 wire n2592;
 wire n2593;
 wire n2594;
 wire n2595;
 wire n2596;
 wire n2597;
 wire n2598;
 wire n2599;
 wire n2600;
 wire n2601;
 wire n2602;
 wire n2603;
 wire n2604;
 wire n2605;
 wire n2606;
 wire n2607;
 wire n2608;
 wire n2609;
 wire n2610;
 wire n2611;
 wire n2612;
 wire n2613;
 wire n2614;
 wire n2615;
 wire n2616;
 wire n2617;
 wire n2618;
 wire n2619;
 wire n2620;
 wire n2621;
 wire n2622;
 wire n2623;
 wire n2624;
 wire n2625;
 wire n2626;
 wire n2627;
 wire n2628;
 wire n2629;
 wire n2630;
 wire n2631;
 wire n2632;
 wire n2633;
 wire n2634;
 wire n2635;
 wire n2636;
 wire n2637;
 wire n2638;
 wire n2639;
 wire n2640;
 wire n2641;
 wire n2642;
 wire n2643;
 wire n2644;
 wire n2645;
 wire n2646;
 wire n2647;
 wire n2648;
 wire n2649;
 wire n2650;
 wire n2651;
 wire n2652;
 wire n2653;
 wire n2654;
 wire n2655;
 wire n2656;
 wire n2657;
 wire n2658;
 wire n2659;
 wire n2660;
 wire n2661;
 wire n2662;
 wire n2663;
 wire n2664;
 wire n2665;
 wire n2666;
 wire n2667;
 wire n2668;
 wire n2669;
 wire n2670;
 wire n2671;
 wire n2672;
 wire n2673;
 wire n2674;
 wire n2675;
 wire n2676;
 wire n2677;
 wire n2678;
 wire n2680;
 wire n2681;
 wire n2682;
 wire n2683;
 wire n2684;
 wire n2685;
 wire n2686;
 wire n2687;
 wire n2688;
 wire n2689;
 wire n2690;
 wire n2691;
 wire n2692;
 wire n2693;
 wire n2694;
 wire n2695;
 wire n2696;
 wire n2697;
 wire n2698;
 wire n2700;
 wire n2701;
 wire n2702;
 wire n2703;
 wire n2704;
 wire n2705;
 wire n2706;
 wire n2707;
 wire n2708;
 wire n2709;
 wire n2711;
 wire n2712;
 wire n2713;
 wire n2714;
 wire n2715;
 wire n2716;
 wire n2717;
 wire n2718;
 wire n2719;
 wire n2720;
 wire n2721;
 wire n2722;
 wire n2723;
 wire n2724;
 wire n2725;
 wire n2726;
 wire n2727;
 wire n2728;
 wire n2729;
 wire n2730;
 wire n2731;
 wire n2732;
 wire n2733;
 wire n2734;
 wire n2735;
 wire n2736;
 wire n2737;
 wire n2738;
 wire n2739;
 wire n2740;
 wire n2741;
 wire n2742;
 wire n2743;
 wire n2744;
 wire n2745;
 wire n2746;
 wire n2747;
 wire n2748;
 wire n2749;
 wire n2750;
 wire n2751;
 wire n2752;
 wire n2753;
 wire n2754;
 wire n2755;
 wire n2756;
 wire n2757;
 wire n2758;
 wire n2759;
 wire n2760;
 wire n2761;
 wire n2762;
 wire n2763;
 wire n2764;
 wire n2765;
 wire n2766;
 wire n2767;
 wire n2768;
 wire n2769;
 wire n2770;
 wire n2771;
 wire n2772;
 wire n2773;
 wire n2774;
 wire n2775;
 wire n2776;
 wire n2777;
 wire n2778;
 wire n2779;
 wire n2780;
 wire n2781;
 wire n2782;
 wire n2783;
 wire n2784;
 wire n2785;
 wire n2786;
 wire n2787;
 wire n2788;
 wire n2789;
 wire n2790;
 wire n2791;
 wire n2792;
 wire n2793;
 wire n2794;
 wire n2795;
 wire n2796;
 wire n2797;
 wire n2798;
 wire n2799;
 wire n2800;
 wire n2801;
 wire n2802;
 wire n2803;
 wire n2804;
 wire n2805;
 wire n2806;
 wire n2807;
 wire n2808;
 wire n2809;
 wire n2810;
 wire n2811;
 wire n2812;
 wire n2813;
 wire n2814;
 wire n2815;
 wire n2816;
 wire n2817;
 wire n2818;
 wire n2819;
 wire n2820;
 wire n2821;
 wire n2822;
 wire n2823;
 wire n2824;
 wire n2825;
 wire n2826;
 wire n2827;
 wire n2828;
 wire n2829;
 wire n2830;
 wire n2831;
 wire n2832;
 wire n2833;
 wire n2834;
 wire n2835;
 wire n2836;
 wire n2837;
 wire n2838;
 wire n2839;
 wire n2840;
 wire n2841;
 wire n2842;
 wire n2843;
 wire n2844;
 wire n2845;
 wire n2846;
 wire n2847;
 wire n2848;
 wire n2849;
 wire n2850;
 wire n2851;
 wire n2852;
 wire n2853;
 wire n2854;
 wire n2855;
 wire n2856;
 wire n2857;
 wire n2858;
 wire n2859;
 wire n2860;
 wire n2861;
 wire n2862;
 wire n2863;
 wire n2864;
 wire n2865;
 wire n2866;
 wire n2867;
 wire n2868;
 wire n2869;
 wire n2870;
 wire n2872;
 wire n2873;
 wire n2874;
 wire n2875;
 wire n2876;
 wire n2877;
 wire n2878;
 wire n2879;
 wire n2880;
 wire n2881;
 wire n2882;
 wire n2883;
 wire n2884;
 wire n2885;
 wire n2886;
 wire n2887;
 wire n2888;
 wire n2889;
 wire n2890;
 wire n2891;
 wire n2892;
 wire n2893;
 wire n2894;
 wire n2895;
 wire n2896;
 wire n2897;
 wire n2898;
 wire n2899;
 wire n2900;
 wire n2901;
 wire n2902;
 wire n2903;
 wire n2904;
 wire n2905;
 wire n2906;
 wire n2907;
 wire n2908;
 wire n2909;
 wire n2910;
 wire n2911;
 wire n2912;
 wire n2913;
 wire n2914;
 wire n2915;
 wire n2916;
 wire n2917;
 wire n2918;
 wire n2919;
 wire n2920;
 wire n2921;
 wire n2922;
 wire n2923;
 wire n2924;
 wire n2925;
 wire n2926;
 wire n2927;
 wire n2928;
 wire n2929;
 wire n2930;
 wire n2931;
 wire n2932;
 wire n2933;
 wire n2934;
 wire n2935;
 wire n2936;
 wire n2937;
 wire n2938;
 wire n2939;
 wire n2940;
 wire n2941;
 wire n2942;
 wire n2943;
 wire n2944;
 wire n2945;
 wire n2946;
 wire n2947;
 wire n2948;
 wire n2949;
 wire n2950;
 wire n2951;
 wire n2952;
 wire n2953;
 wire n2954;
 wire n2955;
 wire n2956;
 wire n2957;
 wire n2958;
 wire n2959;
 wire n2960;
 wire n2961;
 wire n2962;
 wire n2963;
 wire n2964;
 wire n2965;
 wire n2966;
 wire n2967;
 wire n2968;
 wire n2969;
 wire n2970;
 wire n2971;
 wire n2972;
 wire n2973;
 wire n2974;
 wire n2975;
 wire n2976;
 wire n2977;
 wire n2978;
 wire n2979;
 wire n2980;
 wire n2981;
 wire n2982;
 wire n2983;
 wire n2984;
 wire n2985;
 wire n2986;
 wire n2987;
 wire n2988;
 wire n2989;
 wire n2990;
 wire n2991;
 wire n2992;
 wire n2993;
 wire n2994;
 wire n2995;
 wire n2996;
 wire n2997;
 wire n2998;
 wire n2999;
 wire n3000;
 wire n3001;
 wire n3002;
 wire n3003;
 wire n3004;
 wire n3005;
 wire n3006;
 wire n3007;
 wire n3008;
 wire n3009;
 wire n3010;
 wire n3011;
 wire n3012;
 wire n3013;
 wire n3014;
 wire n3015;
 wire n3016;
 wire n3017;
 wire n3018;
 wire n3019;
 wire n3020;
 wire n3021;
 wire n3022;
 wire n3023;
 wire n3024;
 wire n3025;
 wire n3026;
 wire n3027;
 wire n3028;
 wire n3029;
 wire n3030;
 wire n3031;
 wire n3032;
 wire n3033;
 wire n3034;
 wire n3035;
 wire n3036;
 wire n3037;
 wire n3038;
 wire n3039;
 wire n3040;
 wire n3041;
 wire n3042;
 wire n3043;
 wire n3044;
 wire n3045;
 wire n3046;
 wire n3047;
 wire n3048;
 wire n3049;
 wire n3050;
 wire n3051;
 wire n3052;
 wire n3053;
 wire n3054;
 wire n3055;
 wire n3056;
 wire n3057;
 wire n3058;
 wire n3059;
 wire n3060;
 wire n3061;
 wire n3062;
 wire n3063;
 wire n3064;
 wire n3065;
 wire n3066;
 wire n3067;
 wire n3068;
 wire n3069;
 wire n3070;
 wire n3071;
 wire n3072;
 wire n3073;
 wire n3074;
 wire n3075;
 wire n3076;
 wire n3077;
 wire n3078;
 wire n3079;
 wire n3080;
 wire n3081;
 wire n3082;
 wire n3083;
 wire n3084;
 wire n3085;
 wire n3086;
 wire n3087;
 wire n3088;
 wire n3089;
 wire n3090;
 wire n3091;
 wire n3092;
 wire n3093;
 wire n3094;
 wire n3095;
 wire n3096;
 wire n3097;
 wire n3098;
 wire n3099;
 wire n3100;
 wire n3101;
 wire n3102;
 wire n3103;
 wire n3104;
 wire n3105;
 wire n3106;
 wire n3107;
 wire n3108;
 wire n3109;
 wire n3110;
 wire n3111;
 wire n3112;
 wire n3113;
 wire n3114;
 wire n3115;
 wire n3116;
 wire n3117;
 wire n3118;
 wire n3119;
 wire n3120;
 wire n3121;
 wire n3122;
 wire n3123;
 wire n3124;
 wire n3125;
 wire n3126;
 wire n3127;
 wire n3128;
 wire n3129;
 wire n3130;
 wire n3131;
 wire n3132;
 wire n3133;
 wire n3134;
 wire n3135;
 wire n3136;
 wire n3137;
 wire n3138;
 wire n3139;
 wire n3140;
 wire n3141;
 wire n3142;
 wire n3143;
 wire n3144;
 wire n3145;
 wire n3146;
 wire n3147;
 wire n3148;
 wire n3149;
 wire n3150;
 wire n3151;
 wire n3152;
 wire n3153;
 wire n3154;
 wire n3155;
 wire n3156;
 wire n3157;
 wire n3158;
 wire n3159;
 wire n3160;
 wire n3161;
 wire n3162;
 wire n3163;
 wire n3164;
 wire n3165;
 wire n3166;
 wire n3167;
 wire n3168;
 wire n3169;
 wire n3170;
 wire n3171;
 wire n3172;
 wire n3173;
 wire n3174;
 wire n3175;
 wire n3176;
 wire n3177;
 wire n3178;
 wire n3179;
 wire n3180;
 wire n3181;
 wire n3182;
 wire n3183;
 wire n3184;
 wire n3185;
 wire n3186;
 wire n3187;
 wire n3188;
 wire n3189;
 wire n3190;
 wire n3191;
 wire n3192;
 wire n3193;
 wire n3194;
 wire n3195;
 wire n3196;
 wire n3197;
 wire n3198;
 wire n3199;
 wire n3200;
 wire n3201;
 wire n3202;
 wire n3203;
 wire n3204;
 wire n3205;
 wire n3206;
 wire n3207;
 wire n3208;
 wire n3209;
 wire n3210;
 wire n3211;
 wire n3212;
 wire n3213;
 wire n3214;
 wire n3215;
 wire n3216;
 wire n3217;
 wire n3218;
 wire n3219;
 wire n3220;
 wire n3221;
 wire n3222;
 wire n3223;
 wire n3224;
 wire n3225;
 wire n3226;
 wire n3227;
 wire n3228;
 wire n3229;
 wire n3230;
 wire n3231;
 wire n3232;
 wire n3233;
 wire n3234;
 wire n3235;
 wire n3236;
 wire n3237;
 wire n3238;
 wire n3239;
 wire n3240;
 wire n3241;
 wire n3242;
 wire n3243;
 wire n3244;
 wire n3245;
 wire n3246;
 wire n3247;
 wire n3248;
 wire n3249;
 wire n3250;
 wire n3251;
 wire n3252;
 wire n3253;
 wire n3254;
 wire n3255;
 wire n3256;
 wire n3257;
 wire n3258;
 wire n3259;
 wire n3260;
 wire n3261;
 wire n3262;
 wire n3263;
 wire n3264;
 wire n3265;
 wire n3266;
 wire n3267;
 wire n3268;
 wire n3269;
 wire n3270;
 wire n3271;
 wire n3272;
 wire n3273;
 wire n3274;
 wire n3275;
 wire n3276;
 wire n3277;
 wire n3278;
 wire n3279;
 wire n3280;
 wire n3281;
 wire n3282;
 wire n3283;
 wire n3284;
 wire n3285;
 wire n3286;
 wire n3287;
 wire n3288;
 wire n3289;
 wire n3290;
 wire n3291;
 wire n3292;
 wire n3293;
 wire n3294;
 wire n3295;
 wire n3296;
 wire n3297;
 wire n3298;
 wire n3299;
 wire n3300;
 wire n3301;
 wire n3302;
 wire n3303;
 wire n3304;
 wire n3305;
 wire n3306;
 wire n3307;
 wire n3308;
 wire n3309;
 wire n3310;
 wire n3311;
 wire n3312;
 wire n3313;
 wire n3314;
 wire n3315;
 wire n3316;
 wire n3317;
 wire n3318;
 wire n3319;
 wire n3320;
 wire n3321;
 wire n3322;
 wire n3323;
 wire n3324;
 wire n3325;
 wire n3326;
 wire n3327;
 wire n3328;
 wire n3329;
 wire n3330;
 wire n3331;
 wire n3332;
 wire n3333;
 wire n3334;
 wire n3335;
 wire n3336;
 wire n3337;
 wire n3338;
 wire n3339;
 wire n3340;
 wire n3341;
 wire n3342;
 wire n3343;
 wire n3344;
 wire n3345;
 wire n3346;
 wire n3347;
 wire n3348;
 wire n3349;
 wire n3350;
 wire n3351;
 wire n3352;
 wire n3353;
 wire n3354;
 wire n3355;
 wire n3356;
 wire n3357;
 wire n3358;
 wire n3359;
 wire n3360;
 wire n3361;
 wire n3362;
 wire n3363;
 wire n3364;
 wire n3365;
 wire n3366;
 wire n3367;
 wire n3368;
 wire n3369;
 wire n3370;
 wire n3371;
 wire n3372;
 wire n3373;
 wire n3374;
 wire n3375;
 wire n3376;
 wire n3377;
 wire n3378;
 wire n3379;
 wire n3380;
 wire n3381;
 wire n3382;
 wire n3383;
 wire n3384;
 wire n3385;
 wire n3386;
 wire n3387;
 wire n3388;
 wire n3389;
 wire n3390;
 wire n3391;
 wire n3392;
 wire n3393;
 wire n3394;
 wire n3395;
 wire n3396;
 wire n3397;
 wire n3398;
 wire n3399;
 wire n3400;
 wire n3401;
 wire n3402;
 wire n3403;
 wire n3404;
 wire n3405;
 wire n3406;
 wire n3407;
 wire n3408;
 wire n3409;
 wire n3410;
 wire n3411;
 wire n3412;
 wire n3413;
 wire n3414;
 wire n3415;
 wire n3416;
 wire n3417;
 wire n3418;
 wire n3419;
 wire n3420;
 wire n3421;
 wire n3422;
 wire n3423;
 wire n3424;
 wire n3425;
 wire n3426;
 wire n3427;
 wire n3428;
 wire n3429;
 wire n3430;
 wire n3431;
 wire n3432;
 wire n3433;
 wire n3434;
 wire n3435;
 wire n3436;
 wire n3437;
 wire n3438;
 wire n3439;
 wire n3440;
 wire n3441;
 wire n3442;
 wire n3443;
 wire n3444;
 wire n3445;
 wire n3446;
 wire n3447;
 wire n3448;
 wire n3449;
 wire n3450;
 wire n3451;
 wire n3452;
 wire n3453;
 wire n3454;
 wire n3455;
 wire n3456;
 wire n3457;
 wire n3458;
 wire n3459;
 wire n3460;
 wire n3461;
 wire n3462;
 wire n3463;
 wire n3464;
 wire n3465;
 wire n3466;
 wire n3467;
 wire n3468;
 wire n3469;
 wire n3470;
 wire n3471;
 wire n3472;
 wire n3473;
 wire n3474;
 wire n3475;
 wire n3476;
 wire n3477;
 wire n3478;
 wire n3479;
 wire n3480;
 wire n3481;
 wire n3482;
 wire n3483;
 wire n3484;
 wire n3485;
 wire n3486;
 wire n3487;
 wire n3488;
 wire n3489;
 wire n3490;
 wire n3491;
 wire n3492;
 wire n3493;
 wire n3494;
 wire n3495;
 wire n3496;
 wire n3497;
 wire n3498;
 wire n3499;
 wire n3500;
 wire n3501;
 wire n3502;
 wire n3503;
 wire n3504;
 wire n3505;
 wire n3506;
 wire n3507;
 wire n3508;
 wire n3509;
 wire n3510;
 wire n3511;
 wire n3512;
 wire n3513;
 wire n3514;
 wire n3515;
 wire n3516;
 wire n3517;
 wire n3518;
 wire n3519;
 wire n3520;
 wire n3521;
 wire n3522;
 wire n3523;
 wire n3524;
 wire n3525;
 wire n3526;
 wire n3527;
 wire n3528;
 wire n3529;
 wire n3530;
 wire n3531;
 wire n3532;
 wire n3533;
 wire n3535;
 wire n3536;
 wire n3537;
 wire n3538;
 wire n3539;
 wire n3540;
 wire n3541;
 wire n3542;
 wire n3543;
 wire n3544;
 wire n3545;
 wire n3546;
 wire n3547;
 wire n3548;
 wire n3549;
 wire n3550;
 wire n3551;
 wire n3552;
 wire n3553;
 wire n3554;
 wire n3555;
 wire n3556;
 wire n3557;
 wire n3558;
 wire n3559;
 wire n3560;
 wire n3561;
 wire n3562;
 wire n3563;
 wire n3564;
 wire n3565;
 wire n3566;
 wire n3567;
 wire n3568;
 wire n3569;
 wire n3570;
 wire n3571;
 wire n3572;
 wire n3573;
 wire n3574;
 wire n3575;
 wire n3576;
 wire n3577;
 wire n3578;
 wire n3579;
 wire n3580;
 wire n3581;
 wire n3582;
 wire n3583;
 wire n3584;
 wire n3585;
 wire n3586;
 wire n3587;
 wire n3588;
 wire n3589;
 wire n3590;
 wire n3591;
 wire n3592;
 wire n3593;
 wire n3594;
 wire n3595;
 wire n3596;
 wire n3597;
 wire n3598;
 wire n3599;
 wire n3600;
 wire n3601;
 wire n3602;
 wire n3603;
 wire n3604;
 wire n3605;
 wire n3606;
 wire n3607;
 wire n3608;
 wire n3609;
 wire n3610;
 wire n3611;
 wire n3612;
 wire n3613;
 wire n3614;
 wire n3615;
 wire n3616;
 wire n3617;
 wire n3618;
 wire n3619;
 wire n3620;
 wire n3621;
 wire n3622;
 wire n3623;
 wire n3624;
 wire n3625;
 wire n3626;
 wire n3627;
 wire n3628;
 wire n3629;
 wire n3630;
 wire n3631;
 wire n3632;
 wire n3633;
 wire n3634;
 wire n3635;
 wire n3636;
 wire n3637;
 wire n3638;
 wire n3639;
 wire n3640;
 wire n3641;
 wire n3642;
 wire n3643;
 wire n3644;
 wire n3645;
 wire n3646;
 wire n3647;
 wire n3648;
 wire n3649;
 wire n3650;
 wire n3651;
 wire n3652;
 wire n3653;
 wire n3654;
 wire n3655;
 wire n3656;
 wire n3657;
 wire n3658;
 wire n3659;
 wire n3660;
 wire n3661;
 wire n3662;
 wire n3663;
 wire n3664;
 wire n3665;
 wire n3666;
 wire n3667;
 wire n3668;
 wire n3669;
 wire n3670;
 wire n3671;
 wire n3672;
 wire n3673;
 wire n3674;
 wire n3675;
 wire n3676;
 wire n3677;
 wire n3678;
 wire n3679;
 wire n3680;
 wire n3681;
 wire n3682;
 wire n3683;
 wire n3684;
 wire n3685;
 wire n3686;
 wire n3687;
 wire n3688;
 wire n3689;
 wire n3690;
 wire n3691;
 wire n3692;
 wire n3693;
 wire n3694;
 wire n3695;
 wire n3696;
 wire n3697;
 wire n3698;
 wire n3699;
 wire n3700;
 wire n3701;
 wire n3702;
 wire n3703;
 wire n3704;
 wire n3705;
 wire n3706;
 wire n3707;
 wire n3708;
 wire n3709;
 wire n3710;
 wire n3711;
 wire n3712;
 wire n3713;
 wire n3714;
 wire n3715;
 wire n3716;
 wire n3717;
 wire n3718;
 wire n3719;
 wire n3720;
 wire n3721;
 wire n3722;
 wire n3723;
 wire n3724;
 wire n3725;
 wire n3726;
 wire n3727;
 wire n3728;
 wire n3729;
 wire n3730;
 wire n3731;
 wire n3732;
 wire n3733;
 wire n3734;
 wire n3735;
 wire n3736;
 wire n3737;
 wire n3738;
 wire n3739;
 wire n3740;
 wire n3741;
 wire n3742;
 wire n3743;
 wire n3744;
 wire n3745;
 wire n3746;
 wire n3747;
 wire n3748;
 wire n3749;
 wire n3750;
 wire n3751;
 wire n3752;
 wire n3753;
 wire n3754;
 wire n3755;
 wire n3756;
 wire n3757;
 wire n3758;
 wire n3759;
 wire n3760;
 wire n3761;
 wire n3762;
 wire n3763;
 wire n3764;
 wire n3765;
 wire n3766;
 wire n3767;
 wire n3768;
 wire n3769;
 wire n3770;
 wire n3771;
 wire n3772;
 wire n3773;
 wire n3774;
 wire n3775;
 wire n3776;
 wire n3777;
 wire n3778;
 wire n3779;
 wire n3780;
 wire n3781;
 wire n3782;
 wire n3783;
 wire n3784;
 wire n3785;
 wire n3786;
 wire n3787;
 wire n3788;
 wire n3789;
 wire n3790;
 wire n3791;
 wire n3792;
 wire n3793;
 wire n3794;
 wire n3795;
 wire n3796;
 wire n3797;
 wire n3798;
 wire n3799;
 wire n3800;
 wire n3801;
 wire n3802;
 wire n3803;
 wire n3804;
 wire n3805;
 wire n3806;
 wire n3807;
 wire n3808;
 wire n3809;
 wire n3810;
 wire n3811;
 wire n3812;
 wire n3813;
 wire n3814;
 wire n3815;
 wire n3816;
 wire n3817;
 wire n3818;
 wire n3819;
 wire n3820;
 wire n3821;
 wire n3822;
 wire n3823;
 wire n3824;
 wire n3825;
 wire n3826;
 wire n3827;
 wire n3828;
 wire n3829;
 wire n3830;
 wire n3831;
 wire n3832;
 wire n3833;
 wire n3834;
 wire n3835;
 wire n3836;
 wire n3837;
 wire n3838;
 wire n3839;
 wire n3840;
 wire n3841;
 wire n3852;
 wire n3859;
 wire n3860;
 wire n3861;
 wire n3862;
 wire n3863;
 wire n3864;
 wire n3865;
 wire n3866;
 wire n3867;
 wire n3868;
 wire n3869;
 wire n3870;
 wire n3871;
 wire n_RX_EMPTY_FLAG_FLAG_;
 wire n_RX_FULL_FLAG_FLAG_;
 wire n_TX_EMPTY_FLAG_FLAG_;
 wire n_TX_FULL_FLAG_FLAG_;
 wire \rx_fifo_th[0] ;
 wire \rx_fifo_th[1] ;
 wire \rx_fifo_th[2] ;
 wire \rx_fifo_th[3] ;
 wire net60;
 wire \tx_fifo_th[0] ;
 wire \tx_fifo_th[1] ;
 wire \tx_fifo_th[2] ;
 wire \tx_fifo_th[3] ;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net61;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire clknet_leaf_1_HCLK;
 wire clknet_leaf_2_HCLK;
 wire clknet_leaf_3_HCLK;
 wire clknet_leaf_4_HCLK;
 wire clknet_leaf_5_HCLK;
 wire clknet_leaf_6_HCLK;
 wire clknet_leaf_7_HCLK;
 wire clknet_leaf_8_HCLK;
 wire clknet_0_HCLK;
 wire clknet_1_0__leaf_HCLK;
 wire clknet_1_1__leaf_HCLK;
 wire clknet_leaf_0_usb_cdc_clk_48MHz;
 wire clknet_leaf_1_usb_cdc_clk_48MHz;
 wire clknet_leaf_2_usb_cdc_clk_48MHz;
 wire clknet_leaf_3_usb_cdc_clk_48MHz;
 wire clknet_leaf_4_usb_cdc_clk_48MHz;
 wire clknet_leaf_5_usb_cdc_clk_48MHz;
 wire clknet_leaf_6_usb_cdc_clk_48MHz;
 wire clknet_leaf_7_usb_cdc_clk_48MHz;
 wire clknet_leaf_8_usb_cdc_clk_48MHz;
 wire clknet_leaf_9_usb_cdc_clk_48MHz;
 wire clknet_0_usb_cdc_clk_48MHz;
 wire clknet_1_0__leaf_usb_cdc_clk_48MHz;
 wire clknet_1_1__leaf_usb_cdc_clk_48MHz;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;

 sky130_fd_sc_hd__dfrtp_1 CG_REG_reg_0_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1605),
    .RESET_B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(CG_REG_0_));
 sky130_fd_sc_hd__dfrtp_1 CONTROL_REG_reg_0_ (.CLK(clknet_leaf_0_HCLK),
    .D(n1612),
    .RESET_B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(CONTROL_REG_0_));
 sky130_fd_sc_hd__dfrtp_1 ICR_REG_reg_0_ (.CLK(clknet_leaf_1_HCLK),
    .D(N26),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ICR_REG[0] ));
 sky130_fd_sc_hd__dfrtp_1 ICR_REG_reg_1_ (.CLK(clknet_leaf_1_HCLK),
    .D(N27),
    .RESET_B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ICR_REG[1] ));
 sky130_fd_sc_hd__dfrtp_1 ICR_REG_reg_2_ (.CLK(clknet_leaf_1_HCLK),
    .D(N28),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ICR_REG[2] ));
 sky130_fd_sc_hd__dfrtp_1 ICR_REG_reg_3_ (.CLK(clknet_leaf_1_HCLK),
    .D(N29),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ICR_REG[3] ));
 sky130_fd_sc_hd__dfrtp_1 ICR_REG_reg_4_ (.CLK(clknet_leaf_0_HCLK),
    .D(N30),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ICR_REG[4] ));
 sky130_fd_sc_hd__dfrtp_1 ICR_REG_reg_5_ (.CLK(clknet_leaf_0_HCLK),
    .D(N31),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\ICR_REG[5] ));
 sky130_fd_sc_hd__dfrtp_1 IM_REG_reg_0_ (.CLK(clknet_leaf_0_HCLK),
    .D(n1606),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\IM_REG[0] ));
 sky130_fd_sc_hd__dfrtp_1 IM_REG_reg_1_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1607),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\IM_REG[1] ));
 sky130_fd_sc_hd__dfrtp_1 IM_REG_reg_2_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1608),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\IM_REG[2] ));
 sky130_fd_sc_hd__dfrtp_1 IM_REG_reg_3_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1609),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\IM_REG[3] ));
 sky130_fd_sc_hd__dfrtp_1 IM_REG_reg_4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n1610),
    .RESET_B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\IM_REG[4] ));
 sky130_fd_sc_hd__dfrtp_1 IM_REG_reg_5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n1611),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\IM_REG[5] ));
 sky130_fd_sc_hd__dfrtp_1 RIS_REG_reg_0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2127),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RIS_REG[0] ));
 sky130_fd_sc_hd__dfrtp_1 RIS_REG_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2133),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RIS_REG[1] ));
 sky130_fd_sc_hd__dfrtp_1 RIS_REG_reg_2_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1847),
    .RESET_B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RIS_REG[2] ));
 sky130_fd_sc_hd__dfrtp_1 RIS_REG_reg_3_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1849),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RIS_REG[3] ));
 sky130_fd_sc_hd__dfrtp_1 RIS_REG_reg_4_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1846),
    .RESET_B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RIS_REG[4] ));
 sky130_fd_sc_hd__dfrtp_1 RIS_REG_reg_5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2138),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RIS_REG[5] ));
 sky130_fd_sc_hd__dfrtp_1 RXFIFOT_REG_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1613),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\rx_fifo_th[0] ));
 sky130_fd_sc_hd__dfrtp_1 RXFIFOT_REG_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1614),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\rx_fifo_th[1] ));
 sky130_fd_sc_hd__dfrtp_1 RXFIFOT_REG_reg_2_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1615),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\rx_fifo_th[2] ));
 sky130_fd_sc_hd__dfrtp_1 RXFIFOT_REG_reg_3_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1616),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\rx_fifo_th[3] ));
 sky130_fd_sc_hd__dfrtp_1 TXFIFOT_REG_reg_0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n1617),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tx_fifo_th[0] ));
 sky130_fd_sc_hd__dfrtp_1 TXFIFOT_REG_reg_1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n1618),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tx_fifo_th[1] ));
 sky130_fd_sc_hd__dfrtp_1 TXFIFOT_REG_reg_2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n1619),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tx_fifo_th[2] ));
 sky130_fd_sc_hd__dfrtp_1 TXFIFOT_REG_reg_3_ (.CLK(clknet_leaf_7_HCLK),
    .D(n1620),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\tx_fifo_th[3] ));
 sky130_fd_sc_hd__o2bb2ai_1 U2261 (.A1_N(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[3] ),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2299));
 sky130_fd_sc_hd__o2bb2ai_1 U2262 (.A1_N(n3443),
    .A2_N(n2998),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .B2(n2297),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2308));
 sky130_fd_sc_hd__o2bb2ai_1 U2263 (.A1_N(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ),
    .A2_N(n3331),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ),
    .B2(n3331),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3332));
 sky130_fd_sc_hd__o2bb2ai_1 U2264 (.A1_N(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .A2_N(n2669),
    .B1(inst_to_wrap_u_usb_cdc_in_data_ack),
    .B2(n2670),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3350));
 sky130_fd_sc_hd__o2bb2ai_1 U2265 (.A1_N(\IM_REG[0] ),
    .A2_N(n3709),
    .B1(n3143),
    .B2(n2425),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2426));
 sky130_fd_sc_hd__o2bb2ai_4 U2266 (.A1_N(n2803),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[12] ),
    .B1(n2803),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2846));
 sky130_fd_sc_hd__o2bb2ai_1 U2267 (.A1_N(n3050),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[14] ),
    .B1(n3050),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2838));
 sky130_fd_sc_hd__nand4bb_1 U2268 (.A_N(n2776),
    .B_N(n2775),
    .C(n2774),
    .D(n2773),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3033));
 sky130_fd_sc_hd__mux2_1 U2269 (.A0(\RXFIFOLEVEL_REG[3] ),
    .A1(n3541),
    .S(n3533),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1850));
 sky130_fd_sc_hd__o2bb2ai_1 U2270 (.A1_N(\inst_to_wrap_rx_fifo_w_ptr_reg[2] ),
    .A2_N(n3610),
    .B1(\inst_to_wrap_rx_fifo_w_ptr_reg[2] ),
    .B2(n3610),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3546));
 sky130_fd_sc_hd__and3b_2 U2271 (.A_N(n3442),
    .B(n2701),
    .C(n2700),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3438));
 sky130_fd_sc_hd__o2bb2ai_1 U2272 (.A1_N(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ),
    .A2_N(n3177),
    .B1(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ),
    .B2(n3177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3153));
 sky130_fd_sc_hd__o2bb2ai_1 U2273 (.A1_N(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .A2_N(n3357),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .B2(n3357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2320));
 sky130_fd_sc_hd__o2bb2ai_1 U2274 (.A1_N(n2621),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[3] ),
    .B1(n2600),
    .B2(n2599),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2601));
 sky130_fd_sc_hd__o2bb2ai_1 U2275 (.A1_N(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[7] ),
    .A2_N(n2621),
    .B1(n2623),
    .B2(n2622),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2624));
 sky130_fd_sc_hd__and3b_1 U2276 (.A_N(n3081),
    .B(n3083),
    .C(n3082),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3092));
 sky130_fd_sc_hd__o2bb2ai_1 U2277 (.A1_N(n3563),
    .A2_N(\inst_to_wrap_rx_fifo_r_ptr_reg[3] ),
    .B1(n3563),
    .B2(n3517),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1842));
 sky130_fd_sc_hd__o2bb2ai_1 U2278 (.A1_N(n3301),
    .A2_N(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ),
    .B1(net209),
    .B2(n3168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2126));
 sky130_fd_sc_hd__o2bb2ai_1 U2279 (.A1_N(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ),
    .A2_N(n3043),
    .B1(n2336),
    .B2(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2173));
 sky130_fd_sc_hd__o2bb2ai_1 U2280 (.A1_N(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[1] ),
    .A2_N(n3840),
    .B1(n3826),
    .B2(n2414),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_N51));
 sky130_fd_sc_hd__o2bb2ai_1 U2281 (.A1_N(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[6] ),
    .A2_N(n3743),
    .B1(n3740),
    .B2(n3826),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1598));
 sky130_fd_sc_hd__or2_1 U2282 (.A(n2331),
    .B(n2330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2663));
 sky130_fd_sc_hd__nor2b_1 U2283 (.A(n2752),
    .B_N(n2758),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2753));
 sky130_fd_sc_hd__and3b_1 U2284 (.A_N(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_mask_q),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq[0] ),
    .C(n3508),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3567));
 sky130_fd_sc_hd__and3b_1 U2285 (.A_N(n3811),
    .B(n3801),
    .C(n3800),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3803));
 sky130_fd_sc_hd__and3b_1 U2286 (.A_N(n2548),
    .B(n3713),
    .C(n3708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3706));
 sky130_fd_sc_hd__and3b_1 U2287 (.A_N(n3776),
    .B(n3778),
    .C(n3777),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3788));
 sky130_fd_sc_hd__nor2b_2 U2288 (.A(n2662),
    .B_N(\inst_to_wrap_u_usb_cdc_endp[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2806));
 sky130_fd_sc_hd__nor2b_1 U2289 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ),
    .B_N(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2716));
 sky130_fd_sc_hd__nor2b_4 U2290 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[1] ),
    .B_N(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3825));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_HCLK (.A(clknet_1_0__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_HCLK));
 sky130_fd_sc_hd__inv_2 U2292 (.A(net61),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(HREADYOUT));
 sky130_fd_sc_hd__inv_2 U2293 (.A(net62),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(eco_net_7_0));
 sky130_fd_sc_hd__inv_2 U2294 (.A(net63),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(eco_net_13_0));
 sky130_fd_sc_hd__inv_2 U2295 (.A(net64),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(eco_net_16_0));
 sky130_fd_sc_hd__inv_2 U2296 (.A(net65),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(eco_net_19_0));
 sky130_fd_sc_hd__inv_2 U2297 (.A(net66),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(eco_net_21_0));
 sky130_fd_sc_hd__inv_2 U2298 (.A(net67),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(eco_net_23_0));
 sky130_fd_sc_hd__inv_2 U2299 (.A(net68),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(eco_net_28_0));
 sky130_fd_sc_hd__nor4_1 U2300 (.A(n3348),
    .B(n2884),
    .C(n3439),
    .D(n2680),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2732));
 sky130_fd_sc_hd__a21oi_1 U2301 (.A1(n3836),
    .A2(n3715),
    .B1(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net56));
 sky130_fd_sc_hd__clkbuf_1 U2302 (.A(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3862));
 sky130_fd_sc_hd__or3b_1 U2303 (.A(n3499),
    .B(n3348),
    .C_N(n3349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2670));
 sky130_fd_sc_hd__or4_1 U2304 (.A(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[5] ),
    .C(n2863),
    .D(n2327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2328));
 sky130_fd_sc_hd__or2_1 U2305 (.A(n3466),
    .B(n2670),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2761));
 sky130_fd_sc_hd__or4_1 U2306 (.A(n2853),
    .B(n2830),
    .C(n2329),
    .D(n2328),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2330));
 sky130_fd_sc_hd__or2_1 U2307 (.A(n2663),
    .B(n3051),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2778));
 sky130_fd_sc_hd__and4_4 U2308 (.A(n2996),
    .B(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .D(n2885),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3023));
 sky130_fd_sc_hd__or2_2 U2309 (.A(n2743),
    .B(n2778),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3087));
 sky130_fd_sc_hd__or4_1 U2310 (.A(n3467),
    .B(n3466),
    .C(n3465),
    .D(n3464),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3470));
 sky130_fd_sc_hd__or4_2 U2311 (.A(n3466),
    .B(n3477),
    .C(n2698),
    .D(n3465),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3442));
 sky130_fd_sc_hd__or4_2 U2312 (.A(n2821),
    .B(n3052),
    .C(n2335),
    .D(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3043));
 sky130_fd_sc_hd__clkbuf_1 U2313 (.A(eco_net_18_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_20_0));
 sky130_fd_sc_hd__nand2_1 U2314 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2283));
 sky130_fd_sc_hd__inv_2 U2315 (.A(n2283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3389));
 sky130_fd_sc_hd__inv_2 U2316 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3777));
 sky130_fd_sc_hd__inv_2 U2317 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3778));
 sky130_fd_sc_hd__o22ai_1 U2318 (.A1(n3777),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[1] ),
    .B1(n3778),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2284));
 sky130_fd_sc_hd__a221o_1 U2319 (.A1(n3777),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[1] ),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[1] ),
    .B2(n3778),
    .C1(n2284),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2414));
 sky130_fd_sc_hd__nor2_1 U2320 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[0] ),
    .B(n2414),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3840));
 sky130_fd_sc_hd__or3_2 U2321 (.A(\inst_to_wrap_u_usb_cdc_endp[3] ),
    .B(\inst_to_wrap_u_usb_cdc_endp[1] ),
    .C(\inst_to_wrap_u_usb_cdc_endp[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2662));
 sky130_fd_sc_hd__inv_2 U2322 (.A(n2806),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3094));
 sky130_fd_sc_hd__inv_2 U2323 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2820));
 sky130_fd_sc_hd__or3_2 U2324 (.A(n2820),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2774));
 sky130_fd_sc_hd__inv_2 U2325 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3760));
 sky130_fd_sc_hd__or2_2 U2326 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3784));
 sky130_fd_sc_hd__nor2_4 U2327 (.A(n3760),
    .B(n3784),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3089));
 sky130_fd_sc_hd__or2_2 U2328 (.A(n2774),
    .B(n3089),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2908));
 sky130_fd_sc_hd__nor2_1 U2329 (.A(n3094),
    .B(n2908),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3841));
 sky130_fd_sc_hd__inv_2 U2330 (.A(net345),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3839));
 sky130_fd_sc_hd__inv_2 U2331 (.A(net339),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3838));
 sky130_fd_sc_hd__or4_1 U2332 (.A(\last_HADDR[12] ),
    .B(\last_HADDR[13] ),
    .C(\last_HADDR[14] ),
    .D(\last_HADDR[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2286));
 sky130_fd_sc_hd__or4_1 U2333 (.A(\last_HADDR[0] ),
    .B(\last_HADDR[1] ),
    .C(\last_HADDR[5] ),
    .D(\last_HADDR[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2285));
 sky130_fd_sc_hd__or2_2 U2334 (.A(n2990),
    .B(n3095),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3465));
 sky130_fd_sc_hd__nand4_1 U2335 (.A(n2995),
    .B(n2709),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ),
    .D(net211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3377));
 sky130_fd_sc_hd__nor2_1 U2336 (.A(\last_HADDR[7] ),
    .B(n2288),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2356));
 sky130_fd_sc_hd__inv_2 U2337 (.A(n2356),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2354));
 sky130_fd_sc_hd__or4b_1 U2338 (.A(\last_HADDR[3] ),
    .B(\last_HADDR[2] ),
    .C(n2288),
    .D_N(\last_HADDR[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2427));
 sky130_fd_sc_hd__inv_2 U2339 (.A(\last_HADDR[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2355));
 sky130_fd_sc_hd__or4_1 U2340 (.A(\last_HADDR[8] ),
    .B(\last_HADDR[9] ),
    .C(\last_HADDR[10] ),
    .D(\last_HADDR[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2289));
 sky130_fd_sc_hd__or3_1 U2341 (.A(\last_HADDR[7] ),
    .B(n2290),
    .C(n2289),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2548));
 sky130_fd_sc_hd__or3_1 U2342 (.A(\last_HADDR[4] ),
    .B(n2355),
    .C(n2548),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2425));
 sky130_fd_sc_hd__inv_2 U2343 (.A(\last_HADDR[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3708));
 sky130_fd_sc_hd__inv_2 U2344 (.A(\last_HADDR[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2353));
 sky130_fd_sc_hd__a221o_1 U2345 (.A1(\last_HADDR[2] ),
    .A2(\last_HADDR[3] ),
    .B1(n3708),
    .B2(n2353),
    .C1(n2548),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2291));
 sky130_fd_sc_hd__and4_2 U2346 (.A(n2354),
    .B(n2427),
    .C(n2425),
    .D(n2291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_8_0));
 sky130_fd_sc_hd__clkbuf_2 U2347 (.A(eco_net_8_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_9_0));
 sky130_fd_sc_hd__buf_1 U2348 (.A(eco_net_8_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_11_0));
 sky130_fd_sc_hd__clkbuf_1 U2349 (.A(eco_net_11_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_30_0));
 sky130_fd_sc_hd__clkbuf_1 U2350 (.A(eco_net_11_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_10_0));
 sky130_fd_sc_hd__clkbuf_1 U2351 (.A(eco_net_8_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_14_0));
 sky130_fd_sc_hd__clkbuf_1 U2352 (.A(eco_net_14_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_15_0));
 sky130_fd_sc_hd__clkbuf_1 U2353 (.A(eco_net_14_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_12_0));
 sky130_fd_sc_hd__buf_1 U2354 (.A(eco_net_8_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_18_0));
 sky130_fd_sc_hd__clkbuf_1 U2355 (.A(eco_net_18_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_17_0));
 sky130_fd_sc_hd__buf_1 U2356 (.A(eco_net_8_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_24_0));
 sky130_fd_sc_hd__clkbuf_1 U2357 (.A(eco_net_24_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_22_0));
 sky130_fd_sc_hd__clkbuf_1 U2358 (.A(eco_net_24_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_25_0));
 sky130_fd_sc_hd__buf_1 U2359 (.A(eco_net_8_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_27_0));
 sky130_fd_sc_hd__clkbuf_1 U2360 (.A(eco_net_27_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_26_0));
 sky130_fd_sc_hd__clkbuf_1 U2361 (.A(eco_net_27_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_29_0));
 sky130_fd_sc_hd__inv_2 U2362 (.A(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2584));
 sky130_fd_sc_hd__nor2_1 U2363 (.A(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[1] ),
    .B(n2584),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3060));
 sky130_fd_sc_hd__and3_1 U2364 (.A(n3060),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[2] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3057));
 sky130_fd_sc_hd__nor2_1 U2365 (.A(inst_to_wrap_u_usb_cdc_out_err),
    .B(n3057),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3351));
 sky130_fd_sc_hd__inv_2 U2366 (.A(n3351),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3466));
 sky130_fd_sc_hd__nor2_1 U2367 (.A(inst_to_wrap_u_usb_cdc_out_err),
    .B(inst_to_wrap_u_usb_cdc_u_sie_out_eop_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2294));
 sky130_fd_sc_hd__and3_1 U2368 (.A(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3457));
 sky130_fd_sc_hd__nand2_1 U2369 (.A(n3457),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3456));
 sky130_fd_sc_hd__inv_2 U2370 (.A(n3456),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2661));
 sky130_fd_sc_hd__nand2_1 U2371 (.A(n2661),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3454));
 sky130_fd_sc_hd__inv_2 U2372 (.A(n3089),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3083));
 sky130_fd_sc_hd__inv_2 U2373 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3079));
 sky130_fd_sc_hd__inv_2 U2374 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2744));
 sky130_fd_sc_hd__nor2_2 U2375 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[3] ),
    .B(n2744),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2772));
 sky130_fd_sc_hd__and3_1 U2376 (.A(n3079),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .C(n2772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2779));
 sky130_fd_sc_hd__inv_2 U2377 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_fq),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3781));
 sky130_fd_sc_hd__inv_2 U2378 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3765));
 sky130_fd_sc_hd__o22a_2 U2379 (.A1(n3781),
    .A2(n3765),
    .B1(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_fq),
    .B2(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3051));
 sky130_fd_sc_hd__and3_2 U2380 (.A(n3083),
    .B(n2779),
    .C(n3051),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3499));
 sky130_fd_sc_hd__inv_2 U2381 (.A(n3499),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3477));
 sky130_fd_sc_hd__inv_2 U2382 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3771));
 sky130_fd_sc_hd__inv_2 U2383 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3774));
 sky130_fd_sc_hd__or3_1 U2384 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[0] ),
    .B(n3771),
    .C(n3774),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3734));
 sky130_fd_sc_hd__nand2_1 U2385 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_0_),
    .B(n3734),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3776));
 sky130_fd_sc_hd__inv_2 U2386 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3779));
 sky130_fd_sc_hd__inv_2 U2387 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3736));
 sky130_fd_sc_hd__clkinv_2 U2388 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3752));
 sky130_fd_sc_hd__nor2_1 U2389 (.A(n3752),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3731));
 sky130_fd_sc_hd__inv_2 U2390 (.A(n3731),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3780));
 sky130_fd_sc_hd__or4_1 U2391 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .B(n3779),
    .C(n3736),
    .D(n3780),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2293));
 sky130_fd_sc_hd__clkinv_4 U2392 (.A(n3825),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3826));
 sky130_fd_sc_hd__a31o_1 U2393 (.A1(n3083),
    .A2(n3776),
    .A3(n2293),
    .B1(n3826),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2333));
 sky130_fd_sc_hd__o22a_1 U2394 (.A1(n2294),
    .A2(n3454),
    .B1(n3477),
    .B2(n2333),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3091));
 sky130_fd_sc_hd__inv_2 U2395 (.A(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2754));
 sky130_fd_sc_hd__inv_2 U2396 (.A(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2759));
 sky130_fd_sc_hd__inv_2 U2397 (.A(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2757));
 sky130_fd_sc_hd__or2_1 U2398 (.A(n2759),
    .B(n2757),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2752));
 sky130_fd_sc_hd__or2_4 U2399 (.A(\inst_to_wrap_u_usb_cdc_endp[0] ),
    .B(n2662),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2990));
 sky130_fd_sc_hd__inv_2 U2400 (.A(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2814));
 sky130_fd_sc_hd__nand2_1 U2401 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2673));
 sky130_fd_sc_hd__nor2_1 U2402 (.A(n3466),
    .B(n2673),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3467));
 sky130_fd_sc_hd__inv_2 U2403 (.A(n3467),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2316));
 sky130_fd_sc_hd__nor2_1 U2404 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .B(n2316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2667));
 sky130_fd_sc_hd__or4_1 U2405 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[6] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[5] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[4] ),
    .D(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2296));
 sky130_fd_sc_hd__or4_1 U2406 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[0] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[1] ),
    .D(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2295));
 sky130_fd_sc_hd__or2_1 U2407 (.A(n2296),
    .B(n2295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2671));
 sky130_fd_sc_hd__inv_2 U2408 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2685));
 sky130_fd_sc_hd__and3_1 U2409 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[1] ),
    .C(n2685),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3387));
 sky130_fd_sc_hd__nor2_2 U2410 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3012));
 sky130_fd_sc_hd__nor2_1 U2411 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3002));
 sky130_fd_sc_hd__inv_2 U2412 (.A(n3002),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2688));
 sky130_fd_sc_hd__nor2_2 U2413 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .B(n2688),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2959));
 sky130_fd_sc_hd__inv_2 U2414 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3368));
 sky130_fd_sc_hd__nor2_1 U2415 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .B(n3368),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3372));
 sky130_fd_sc_hd__and3_1 U2416 (.A(n3012),
    .B(n2959),
    .C(n3372),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2909));
 sky130_fd_sc_hd__a21boi_1 U2417 (.A1(n3387),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .B1_N(n2909),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2672));
 sky130_fd_sc_hd__nand2b_1 U2418 (.A_N(n2671),
    .B(n2672),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3348));
 sky130_fd_sc_hd__inv_2 U2419 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2697));
 sky130_fd_sc_hd__nor2_1 U2420 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ),
    .B(n2697),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3349));
 sky130_fd_sc_hd__nand2b_1 U2421 (.A_N(n2667),
    .B(n2761),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2318));
 sky130_fd_sc_hd__and3_1 U2422 (.A(n2814),
    .B(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q),
    .C(n2318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2314));
 sky130_fd_sc_hd__inv_2 U2423 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3394));
 sky130_fd_sc_hd__or4_2 U2424 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[2] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .D(n3394),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2687));
 sky130_fd_sc_hd__inv_2 U2425 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2786));
 sky130_fd_sc_hd__and3_1 U2426 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[2] ),
    .B(n3394),
    .C(n2786),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2885));
 sky130_fd_sc_hd__clkinv_2 U2427 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3359));
 sky130_fd_sc_hd__inv_2 U2428 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2884));
 sky130_fd_sc_hd__clkinv_2 U2429 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3440));
 sky130_fd_sc_hd__inv_2 U2430 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3361));
 sky130_fd_sc_hd__nor2_1 U2431 (.A(n3440),
    .B(n3361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3027));
 sky130_fd_sc_hd__inv_2 U2432 (.A(n3027),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3363));
 sky130_fd_sc_hd__nor2_2 U2433 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .B(n3363),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3418));
 sky130_fd_sc_hd__inv_2 U2434 (.A(n3418),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2962));
 sky130_fd_sc_hd__or4_1 U2435 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .B(n3359),
    .C(n2884),
    .D(n2962),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2297));
 sky130_fd_sc_hd__inv_2 U2436 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3010));
 sky130_fd_sc_hd__and3_1 U2437 (.A(n3010),
    .B(n3361),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3416));
 sky130_fd_sc_hd__inv_2 U2438 (.A(n3416),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2886));
 sky130_fd_sc_hd__nor2_1 U2439 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(n2886),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3443));
 sky130_fd_sc_hd__inv_2 U2440 (.A(n3012),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2956));
 sky130_fd_sc_hd__clkinv_2 U2441 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3005));
 sky130_fd_sc_hd__nor2_1 U2442 (.A(n2956),
    .B(n3005),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2998));
 sky130_fd_sc_hd__inv_2 U2443 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2306));
 sky130_fd_sc_hd__inv_2 U2444 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2923));
 sky130_fd_sc_hd__a22oi_1 U2445 (.A1(n3361),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[0] ),
    .B1(n3440),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2298));
 sky130_fd_sc_hd__o221a_1 U2446 (.A1(n3440),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[1] ),
    .B1(n3361),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[0] ),
    .C1(n2298),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2304));
 sky130_fd_sc_hd__inv_1 U2447 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2300));
 sky130_fd_sc_hd__o221a_1 U2448 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[2] ),
    .A2(n3010),
    .B1(n2300),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .C1(n2299),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2303));
 sky130_fd_sc_hd__a22oi_1 U2449 (.A1(n3359),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[6] ),
    .B1(n3005),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2301));
 sky130_fd_sc_hd__o221a_1 U2450 (.A1(n3359),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[6] ),
    .B1(n3005),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[4] ),
    .C1(n2301),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2302));
 sky130_fd_sc_hd__and3_1 U2451 (.A(n2304),
    .B(n2303),
    .C(n2302),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2305));
 sky130_fd_sc_hd__o221a_1 U2452 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .A2(n2306),
    .B1(n2923),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[5] ),
    .C1(n2305),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2307));
 sky130_fd_sc_hd__a31o_1 U2453 (.A1(n2885),
    .A2(n3368),
    .A3(n2308),
    .B1(n2307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2309));
 sky130_fd_sc_hd__nor2_1 U2454 (.A(n3499),
    .B(n2309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2317));
 sky130_fd_sc_hd__and3_1 U2455 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ),
    .C(n2317),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2669));
 sky130_fd_sc_hd__and3_1 U2456 (.A(n2814),
    .B(n3351),
    .C(n2669),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2996));
 sky130_fd_sc_hd__o211a_1 U2457 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ),
    .A2(n2687),
    .B1(n2996),
    .C1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2310));
 sky130_fd_sc_hd__a211o_1 U2458 (.A1(n2806),
    .A2(inst_to_wrap_u_usb_cdc_bulk_in_valid),
    .B1(n2314),
    .C1(n2310),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2311));
 sky130_fd_sc_hd__o31a_1 U2459 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[3] ),
    .A2(n2754),
    .A3(n2752),
    .B1(n2311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3071));
 sky130_fd_sc_hd__or2_4 U2460 (.A(n2774),
    .B(n2744),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3070));
 sky130_fd_sc_hd__clkinv_2 U2461 (.A(n3070),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2821));
 sky130_fd_sc_hd__nand2_1 U2462 (.A(n3071),
    .B(n2821),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2745));
 sky130_fd_sc_hd__nor2_2 U2463 (.A(n2774),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3047));
 sky130_fd_sc_hd__inv_2 U2464 (.A(n2311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2313));
 sky130_fd_sc_hd__inv_2 U2465 (.A(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2751));
 sky130_fd_sc_hd__or4_1 U2466 (.A(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[2] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[1] ),
    .D(n2751),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2312));
 sky130_fd_sc_hd__and3_2 U2467 (.A(n2814),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ),
    .C(n2697),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3038));
 sky130_fd_sc_hd__a211oi_2 U2468 (.A1(n2313),
    .A2(n2312),
    .B1(n3038),
    .C1(n2662),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3046));
 sky130_fd_sc_hd__nand2_1 U2469 (.A(n3047),
    .B(n3046),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3072));
 sky130_fd_sc_hd__nor2_1 U2470 (.A(n2314),
    .B(n2313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3073));
 sky130_fd_sc_hd__nand2b_1 U2471 (.A_N(n3072),
    .B(n3073),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2746));
 sky130_fd_sc_hd__inv_2 U2472 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2575));
 sky130_fd_sc_hd__inv_2 U2473 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3792));
 sky130_fd_sc_hd__nand2_2 U2474 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3793));
 sky130_fd_sc_hd__a31o_4 U2475 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[1] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[2] ),
    .A3(n3792),
    .B1(n3793),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2626));
 sky130_fd_sc_hd__or3_1 U2476 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[0] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2583));
 sky130_fd_sc_hd__or2_1 U2477 (.A(n2626),
    .B(n2583),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3830));
 sky130_fd_sc_hd__or2_1 U2478 (.A(n2575),
    .B(n3830),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2562));
 sky130_fd_sc_hd__inv_2 U2479 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2567));
 sky130_fd_sc_hd__nand2_1 U2480 (.A(n2567),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3716));
 sky130_fd_sc_hd__inv_2 U2481 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2565));
 sky130_fd_sc_hd__nand2_1 U2482 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[1] ),
    .B(n2565),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2581));
 sky130_fd_sc_hd__and2_1 U2483 (.A(n3716),
    .B(n2581),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2334));
 sky130_fd_sc_hd__or2_1 U2484 (.A(n3089),
    .B(n2334),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2572));
 sky130_fd_sc_hd__nor2_1 U2485 (.A(n2562),
    .B(n2572),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2595));
 sky130_fd_sc_hd__inv_2 U2486 (.A(n2595),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2599));
 sky130_fd_sc_hd__a32o_1 U2487 (.A1(n3091),
    .A2(n2745),
    .A3(n2746),
    .B1(n3091),
    .B2(n2599),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3095));
 sky130_fd_sc_hd__a22o_1 U2488 (.A1(n3499),
    .A2(n3349),
    .B1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q),
    .B2(n2669),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2315));
 sky130_fd_sc_hd__or4b_2 U2489 (.A(n3466),
    .B(n3465),
    .C(n2667),
    .D_N(n2315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3365));
 sky130_fd_sc_hd__nor2_2 U2490 (.A(n3010),
    .B(n3363),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3004));
 sky130_fd_sc_hd__and3_1 U2491 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .C(n3004),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3357));
 sky130_fd_sc_hd__a21oi_1 U2492 (.A1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q),
    .A2(n2317),
    .B1(n2316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2319));
 sky130_fd_sc_hd__or3_2 U2493 (.A(n2319),
    .B(n3465),
    .C(n2318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3367));
 sky130_fd_sc_hd__a2bb2o_1 U2494 (.A1_N(n3365),
    .A2_N(n2320),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .B2(n3367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1917));
 sky130_fd_sc_hd__inv_2 U2495 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2803));
 sky130_fd_sc_hd__inv_2 U2496 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3065));
 sky130_fd_sc_hd__inv_2 U2497 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2616));
 sky130_fd_sc_hd__clkinv_2 U2498 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3049));
 sky130_fd_sc_hd__inv_2 U2499 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2639));
 sky130_fd_sc_hd__inv_2 U2500 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2644));
 sky130_fd_sc_hd__clkinv_2 U2501 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3050));
 sky130_fd_sc_hd__inv_2 U2502 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2611));
 sky130_fd_sc_hd__a22o_1 U2503 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[5] ),
    .B1(n3050),
    .B2(n2611),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2321));
 sky130_fd_sc_hd__a221o_1 U2504 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[3] ),
    .B1(n2644),
    .B2(n2803),
    .C1(n2321),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2322));
 sky130_fd_sc_hd__a221o_1 U2505 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[4] ),
    .B1(n3049),
    .B2(n2639),
    .C1(n2322),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2323));
 sky130_fd_sc_hd__a221o_1 U2506 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[6] ),
    .B1(n3065),
    .B2(n2616),
    .C1(n2323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3048));
 sky130_fd_sc_hd__or3b_2 U2507 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ),
    .C_N(n2772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2819));
 sky130_fd_sc_hd__nand2_1 U2508 (.A(n2402),
    .B(n3869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2404));
 sky130_fd_sc_hd__or2_1 U2509 (.A(n3048),
    .B(n2819),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3081));
 sky130_fd_sc_hd__inv_2 U2510 (.A(n3038),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2596));
 sky130_fd_sc_hd__inv_2 U2511 (.A(inst_to_wrap_u_usb_cdc_bulk_out_nak),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3495));
 sky130_fd_sc_hd__nor2_1 U2512 (.A(n3094),
    .B(n3495),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2767));
 sky130_fd_sc_hd__inv_2 U2513 (.A(n2767),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2765));
 sky130_fd_sc_hd__inv_2 U2514 (.A(n2779),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2743));
 sky130_fd_sc_hd__mux2_1 U2515 (.A0(n3065),
    .A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .S(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2840));
 sky130_fd_sc_hd__inv_2 U2516 (.A(n2840),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2841));
 sky130_fd_sc_hd__a2bb2o_1 U2517 (.A1_N(n3049),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[15] ),
    .B1(n3049),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2831));
 sky130_fd_sc_hd__inv_2 U2518 (.A(n2831),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2830));
 sky130_fd_sc_hd__inv_2 U2519 (.A(n2838),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2837));
 sky130_fd_sc_hd__mux2_1 U2520 (.A0(n2830),
    .A1(n2831),
    .S(n2837),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2835));
 sky130_fd_sc_hd__inv_2 U2521 (.A(n2835),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2833));
 sky130_fd_sc_hd__mux2_1 U2522 (.A0(n2840),
    .A1(n2841),
    .S(n2833),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2325));
 sky130_fd_sc_hd__nand2_1 U2523 (.A(n2325),
    .B(n2846),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2331));
 sky130_fd_sc_hd__o2bb2a_1 U2524 (.A1_N(n2616),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[9] ),
    .B1(n2616),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2851));
 sky130_fd_sc_hd__inv_2 U2525 (.A(n2851),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2853));
 sky130_fd_sc_hd__inv_2 U2526 (.A(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2829));
 sky130_fd_sc_hd__or4_1 U2527 (.A(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[3] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[2] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[4] ),
    .D(n2829),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2329));
 sky130_fd_sc_hd__o2bb2a_1 U2528 (.A1_N(n2639),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[11] ),
    .B1(n2639),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2843));
 sky130_fd_sc_hd__inv_2 U2529 (.A(n2843),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2845));
 sky130_fd_sc_hd__o2bb2a_1 U2530 (.A1_N(n2611),
    .A2_N(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[10] ),
    .B1(n2611),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2850));
 sky130_fd_sc_hd__mux2_1 U2531 (.A0(n2843),
    .A1(n2845),
    .S(n2850),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2848));
 sky130_fd_sc_hd__fa_1 U2532 (.A(n2325),
    .B(n2846),
    .CIN(n2848),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2856));
 sky130_fd_sc_hd__inv_2 U2533 (.A(n2856),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2855));
 sky130_fd_sc_hd__mux2_1 U2534 (.A0(n2853),
    .A1(n2851),
    .S(n2855),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2860));
 sky130_fd_sc_hd__fa_2 U2535 (.A(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[8] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ),
    .CIN(n2860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2863));
 sky130_fd_sc_hd__or2_1 U2536 (.A(n2843),
    .B(n2850),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2326));
 sky130_fd_sc_hd__or4_1 U2537 (.A(n2835),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[6] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[7] ),
    .D(n2326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2327));
 sky130_fd_sc_hd__a21o_1 U2538 (.A1(n2596),
    .A2(n2765),
    .B1(n3087),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2332));
 sky130_fd_sc_hd__a22o_1 U2539 (.A1(n2806),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[1] ),
    .B1(n2814),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2805));
 sky130_fd_sc_hd__inv_2 U2540 (.A(n2805),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2816));
 sky130_fd_sc_hd__nand2_1 U2541 (.A(n3046),
    .B(n2816),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2569));
 sky130_fd_sc_hd__nand2_1 U2542 (.A(n3047),
    .B(n2569),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2602));
 sky130_fd_sc_hd__o211a_1 U2543 (.A1(n2803),
    .A2(n3081),
    .B1(n2332),
    .C1(n2602),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2336));
 sky130_fd_sc_hd__o21a_2 U2544 (.A1(n2334),
    .A2(n2562),
    .B1(n2333),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3029));
 sky130_fd_sc_hd__nor2_2 U2545 (.A(n3089),
    .B(n3029),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3045));
 sky130_fd_sc_hd__clkinv_4 U2546 (.A(n3045),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3074));
 sky130_fd_sc_hd__inv_2 U2547 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3056));
 sky130_fd_sc_hd__or3_1 U2548 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[3] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2748));
 sky130_fd_sc_hd__nor2_1 U2549 (.A(n3056),
    .B(n2748),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3052));
 sky130_fd_sc_hd__and2_1 U2550 (.A(n2778),
    .B(n2779),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2335));
 sky130_fd_sc_hd__or2_1 U2551 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[3] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2741));
 sky130_fd_sc_hd__o221a_1 U2552 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .A2(n2741),
    .B1(n3056),
    .B2(n2820),
    .C1(n3045),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2773));
 sky130_fd_sc_hd__nand2_1 U2553 (.A(n2773),
    .B(n3079),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2866));
 sky130_fd_sc_hd__clkbuf_8 U2554 (.A(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3852));
 sky130_fd_sc_hd__a21boi_1 U2555 (.A1(net293),
    .A2(net303),
    .B1_N(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1576));
 sky130_fd_sc_hd__clkbuf_1 U2556 (.A(net294),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3864));
 sky130_fd_sc_hd__buf_8 U2557 (.A(net297),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3861));
 sky130_fd_sc_hd__clkbuf_1 U2558 (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3868));
 sky130_fd_sc_hd__clkbuf_8 U2559 (.A(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3860));
 sky130_fd_sc_hd__buf_6 U2560 (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3859));
 sky130_fd_sc_hd__clkbuf_1 U2561 (.A(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3866));
 sky130_fd_sc_hd__clkbuf_1 U2562 (.A(n1576),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3867));
 sky130_fd_sc_hd__clkbuf_1 U2563 (.A(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3863));
 sky130_fd_sc_hd__buf_1 U2564 (.A(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3865));
 sky130_fd_sc_hd__inv_2 U2565 (.A(n_RX_FULL_FLAG_FLAG_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3513));
 sky130_fd_sc_hd__and3_4 U2566 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq[0] ),
    .B(n3838),
    .C(n3513),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3524));
 sky130_fd_sc_hd__clkinv_2 U2567 (.A(n3524),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3609));
 sky130_fd_sc_hd__nand2_1 U2568 (.A(last_HTRANS_1_),
    .B(last_HSEL),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2337));
 sky130_fd_sc_hd__or4_1 U2569 (.A(\last_HADDR[4] ),
    .B(\last_HADDR[3] ),
    .C(n3708),
    .D(n2548),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2342));
 sky130_fd_sc_hd__or3_2 U2570 (.A(last_HWRITE),
    .B(n2337),
    .C(n2342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3520));
 sky130_fd_sc_hd__a21o_1 U2571 (.A1(n_RX_EMPTY_FLAG_FLAG_),
    .A2(n3609),
    .B1(n3520),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3563));
 sky130_fd_sc_hd__inv_2 U2572 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3549));
 sky130_fd_sc_hd__and3_1 U2573 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .B(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .C(n3549),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2481));
 sky130_fd_sc_hd__and3_1 U2574 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .B(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .C(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2338));
 sky130_fd_sc_hd__o2bb2a_1 U2575 (.A1_N(net207),
    .A2_N(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B1(n2338),
    .B2(n3549),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3517));
 sky130_fd_sc_hd__a22o_1 U2576 (.A1(\RIS_REG[1] ),
    .A2(\IM_REG[1] ),
    .B1(\RIS_REG[3] ),
    .B2(\IM_REG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2341));
 sky130_fd_sc_hd__a22o_1 U2577 (.A1(\RIS_REG[0] ),
    .A2(\IM_REG[0] ),
    .B1(\IM_REG[4] ),
    .B2(\RIS_REG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2340));
 sky130_fd_sc_hd__a22o_1 U2578 (.A1(\RIS_REG[2] ),
    .A2(\IM_REG[2] ),
    .B1(\RIS_REG[5] ),
    .B2(\IM_REG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2339));
 sky130_fd_sc_hd__or3_1 U2579 (.A(n2341),
    .B(n2340),
    .C(n2339),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net59));
 sky130_fd_sc_hd__clkinv_2 U2580 (.A(n2342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2494));
 sky130_fd_sc_hd__and3_4 U2581 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .B(\inst_to_wrap_rx_fifo_r_ptr_reg[3] ),
    .C(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2479));
 sky130_fd_sc_hd__clkinv_2 U2582 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3547));
 sky130_fd_sc_hd__and3_4 U2583 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .B(n3549),
    .C(n3547),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2478));
 sky130_fd_sc_hd__a22o_1 U2584 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[121] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2352));
 sky130_fd_sc_hd__clkinv_2 U2585 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3559));
 sky130_fd_sc_hd__clkinv_2 U2586 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3560));
 sky130_fd_sc_hd__and3_4 U2587 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[3] ),
    .B(n3560),
    .C(n3547),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2480));
 sky130_fd_sc_hd__a22o_1 U2588 (.A1(n2481),
    .A2(\inst_to_wrap_rx_fifo_array_reg[57] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2345));
 sky130_fd_sc_hd__and3_4 U2589 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[3] ),
    .B(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .C(n3560),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2483));
 sky130_fd_sc_hd__and3_4 U2590 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[3] ),
    .B(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .C(n3547),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2482));
 sky130_fd_sc_hd__a22o_1 U2591 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[105] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2344));
 sky130_fd_sc_hd__and3_4 U2592 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .B(n3560),
    .C(n3549),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2485));
 sky130_fd_sc_hd__and3_4 U2593 (.A(n3560),
    .B(n3549),
    .C(n3547),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2484));
 sky130_fd_sc_hd__a22o_1 U2594 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[41] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2343));
 sky130_fd_sc_hd__or4_1 U2595 (.A(n3559),
    .B(n2345),
    .C(n2344),
    .D(n2343),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2351));
 sky130_fd_sc_hd__a22o_1 U2596 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[113] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2350));
 sky130_fd_sc_hd__a22o_1 U2597 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[49] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2348));
 sky130_fd_sc_hd__a22o_1 U2598 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[97] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2347));
 sky130_fd_sc_hd__a22o_1 U2599 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[33] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2346));
 sky130_fd_sc_hd__or4_1 U2600 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2348),
    .C(n2347),
    .D(n2346),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2349));
 sky130_fd_sc_hd__o22a_1 U2601 (.A1(n2352),
    .A2(n2351),
    .B1(n2350),
    .B2(n2349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2363));
 sky130_fd_sc_hd__and3_2 U2602 (.A(\last_HADDR[2] ),
    .B(n2356),
    .C(n2355),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2460));
 sky130_fd_sc_hd__or3_1 U2603 (.A(\last_HADDR[3] ),
    .B(n2353),
    .C(n2548),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2357));
 sky130_fd_sc_hd__nor2_1 U2604 (.A(n3708),
    .B(n2357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3703));
 sky130_fd_sc_hd__a22o_1 U2605 (.A1(n2460),
    .A2(\RIS_REG[1] ),
    .B1(n3703),
    .B2(\rx_fifo_th[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2362));
 sky130_fd_sc_hd__nor2_2 U2606 (.A(n2355),
    .B(n2354),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3709));
 sky130_fd_sc_hd__o211a_1 U2607 (.A1(\RIS_REG[1] ),
    .A2(n3708),
    .B1(n3709),
    .C1(\IM_REG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2360));
 sky130_fd_sc_hd__nor2_1 U2608 (.A(n3708),
    .B(n2425),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2429));
 sky130_fd_sc_hd__and3_2 U2609 (.A(n2356),
    .B(n2355),
    .C(n3708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2495));
 sky130_fd_sc_hd__a22o_1 U2610 (.A1(\RXFIFOLEVEL_REG[1] ),
    .A2(n2429),
    .B1(n2495),
    .B2(\ICR_REG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2359));
 sky130_fd_sc_hd__nor2_1 U2611 (.A(\last_HADDR[2] ),
    .B(n2425),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2390));
 sky130_fd_sc_hd__nor2_1 U2612 (.A(\last_HADDR[2] ),
    .B(n2357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3700));
 sky130_fd_sc_hd__a22o_1 U2613 (.A1(\TXFIFOLEVEL_REG[1] ),
    .A2(n2390),
    .B1(n3700),
    .B2(\tx_fifo_th[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2358));
 sky130_fd_sc_hd__or4_1 U2614 (.A(eco_net_9_0),
    .B(n2360),
    .C(n2359),
    .D(n2358),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2361));
 sky130_fd_sc_hd__a211o_1 U2615 (.A1(n2494),
    .A2(n2363),
    .B1(n2362),
    .C1(n2361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_0));
 sky130_fd_sc_hd__a22o_1 U2616 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[123] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2373));
 sky130_fd_sc_hd__a22o_1 U2617 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[59] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2366));
 sky130_fd_sc_hd__a22o_1 U2618 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[107] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2365));
 sky130_fd_sc_hd__a22o_1 U2619 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[43] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2364));
 sky130_fd_sc_hd__or4_1 U2620 (.A(n3559),
    .B(n2366),
    .C(n2365),
    .D(n2364),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2372));
 sky130_fd_sc_hd__a22o_1 U2621 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[115] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2371));
 sky130_fd_sc_hd__a22o_1 U2622 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[51] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2369));
 sky130_fd_sc_hd__a22o_1 U2623 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[99] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2368));
 sky130_fd_sc_hd__a22o_1 U2624 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[35] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2367));
 sky130_fd_sc_hd__or4_1 U2625 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2369),
    .C(n2368),
    .D(n2367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2370));
 sky130_fd_sc_hd__o22a_1 U2626 (.A1(n2373),
    .A2(n2372),
    .B1(n2371),
    .B2(n2370),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2379));
 sky130_fd_sc_hd__a22o_1 U2627 (.A1(n2460),
    .A2(\RIS_REG[3] ),
    .B1(n3703),
    .B2(\rx_fifo_th[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2378));
 sky130_fd_sc_hd__o211a_1 U2628 (.A1(\RIS_REG[3] ),
    .A2(n3708),
    .B1(n3709),
    .C1(\IM_REG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2376));
 sky130_fd_sc_hd__a22o_1 U2629 (.A1(\RXFIFOLEVEL_REG[3] ),
    .A2(n2429),
    .B1(n2495),
    .B2(\ICR_REG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2375));
 sky130_fd_sc_hd__a22o_1 U2630 (.A1(\TXFIFOLEVEL_REG[3] ),
    .A2(n2390),
    .B1(n3700),
    .B2(\tx_fifo_th[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2374));
 sky130_fd_sc_hd__or4_1 U2631 (.A(eco_net_9_0),
    .B(n2376),
    .C(n2375),
    .D(n2374),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2377));
 sky130_fd_sc_hd__a211o_1 U2632 (.A1(n2494),
    .A2(n2379),
    .B1(n2378),
    .C1(n2377),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_2_0));
 sky130_fd_sc_hd__a22o_1 U2633 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[122] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2389));
 sky130_fd_sc_hd__a22o_1 U2634 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[58] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2382));
 sky130_fd_sc_hd__a22o_1 U2635 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[106] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2381));
 sky130_fd_sc_hd__a22o_1 U2636 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[42] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2380));
 sky130_fd_sc_hd__or4_1 U2637 (.A(n3559),
    .B(n2382),
    .C(n2381),
    .D(n2380),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2388));
 sky130_fd_sc_hd__a22o_1 U2638 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[114] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2387));
 sky130_fd_sc_hd__a22o_1 U2639 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[50] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2385));
 sky130_fd_sc_hd__a22o_1 U2640 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[98] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2384));
 sky130_fd_sc_hd__a22o_1 U2641 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[34] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2383));
 sky130_fd_sc_hd__or4_1 U2642 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2385),
    .C(n2384),
    .D(n2383),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2386));
 sky130_fd_sc_hd__o22a_1 U2643 (.A1(n2389),
    .A2(n2388),
    .B1(n2387),
    .B2(n2386),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2396));
 sky130_fd_sc_hd__a22o_1 U2644 (.A1(n2460),
    .A2(\RIS_REG[2] ),
    .B1(n3703),
    .B2(\rx_fifo_th[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2395));
 sky130_fd_sc_hd__o211a_1 U2645 (.A1(\RIS_REG[2] ),
    .A2(n3708),
    .B1(n3709),
    .C1(\IM_REG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2393));
 sky130_fd_sc_hd__a22o_1 U2646 (.A1(\RXFIFOLEVEL_REG[2] ),
    .A2(n2429),
    .B1(n2495),
    .B2(\ICR_REG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2392));
 sky130_fd_sc_hd__a22o_1 U2647 (.A1(\TXFIFOLEVEL_REG[2] ),
    .A2(n2390),
    .B1(n3700),
    .B2(\tx_fifo_th[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2391));
 sky130_fd_sc_hd__or4_1 U2648 (.A(eco_net_9_0),
    .B(n2393),
    .C(n2392),
    .D(n2391),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2394));
 sky130_fd_sc_hd__a211o_1 U2649 (.A1(n2494),
    .A2(n2396),
    .B1(n2395),
    .C1(n2394),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_1_0));
 sky130_fd_sc_hd__and3_1 U2650 (.A(n3825),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[17] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2547));
 sky130_fd_sc_hd__or2_1 U2651 (.A(n2547),
    .B(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2250));
 sky130_fd_sc_hd__nor2_2 U2652 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3722));
 sky130_fd_sc_hd__inv_4 U2653 (.A(n3722),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(net60));
 sky130_fd_sc_hd__inv_2 U2654 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3333));
 sky130_fd_sc_hd__inv_2 U2655 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3331));
 sky130_fd_sc_hd__inv_2 U2656 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3336));
 sky130_fd_sc_hd__nor2_1 U2657 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2398));
 sky130_fd_sc_hd__nand2_1 U2658 (.A(n3336),
    .B(n2398),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2399));
 sky130_fd_sc_hd__o21a_1 U2659 (.A1(n3336),
    .A2(n2398),
    .B1(n2399),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2401));
 sky130_fd_sc_hd__or2_1 U2660 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ),
    .B(n2399),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2405));
 sky130_fd_sc_hd__inv_1 U2661 (.A(n2405),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2397));
 sky130_fd_sc_hd__or4_2 U2662 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .C(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ),
    .D(n3333),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3116));
 sky130_fd_sc_hd__a22o_1 U2663 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .A2(n2401),
    .B1(n2397),
    .B2(n3116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2409));
 sky130_fd_sc_hd__a21oi_1 U2664 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .B1(n2398),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2400));
 sky130_fd_sc_hd__a22o_1 U2665 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ),
    .B2(n2400),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2408));
 sky130_fd_sc_hd__and2_1 U2666 (.A(n2399),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2406));
 sky130_fd_sc_hd__o22a_1 U2667 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .A2(n2401),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ),
    .B2(n2400),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2402));
 sky130_fd_sc_hd__o22a_1 U2668 (.A1(n2406),
    .A2(n3333),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3869));
 sky130_fd_sc_hd__inv_2 U2669 (.A(n3836),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3870));
 sky130_fd_sc_hd__a22o_1 U2670 (.A1(n2406),
    .A2(n3333),
    .B1(n2405),
    .B2(n2404),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2407));
 sky130_fd_sc_hd__o31a_1 U2671 (.A1(n2409),
    .A2(n2408),
    .A3(n2407),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2410));
 sky130_fd_sc_hd__and4_1 U2672 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[1] ),
    .C(n2410),
    .D(n3839),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3123));
 sky130_fd_sc_hd__clkinv_2 U2673 (.A(n3123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3121));
 sky130_fd_sc_hd__nor2_1 U2674 (.A(n3331),
    .B(n3121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3118));
 sky130_fd_sc_hd__and2_1 U2675 (.A(n3333),
    .B(n3118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3120));
 sky130_fd_sc_hd__and3_2 U2676 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .C(n3120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3320));
 sky130_fd_sc_hd__clkinv_2 U2677 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3337));
 sky130_fd_sc_hd__clkinv_2 U2678 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3325));
 sky130_fd_sc_hd__a221o_1 U2679 (.A1(n3116),
    .A2(n3325),
    .B1(n3116),
    .B2(n3331),
    .C1(n3121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3117));
 sky130_fd_sc_hd__a32o_1 U2680 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[3] ),
    .A2(n3337),
    .A3(n3116),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[3] ),
    .B2(n3117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2411));
 sky130_fd_sc_hd__or2_1 U2681 (.A(n3320),
    .B(n2411),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2153));
 sky130_fd_sc_hd__or2_1 U2682 (.A(n2820),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2412));
 sky130_fd_sc_hd__and3_1 U2683 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ),
    .C(n2772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2592));
 sky130_fd_sc_hd__clkinv_2 U2684 (.A(n2592),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2617));
 sky130_fd_sc_hd__a21oi_1 U2685 (.A1(n2412),
    .A2(n2617),
    .B1(n3089),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3790));
 sky130_fd_sc_hd__or2_1 U2686 (.A(n3790),
    .B(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2413));
 sky130_fd_sc_hd__nor2b_1 U2687 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[0] ),
    .B_N(n2413),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_N30));
 sky130_fd_sc_hd__o211a_1 U2688 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[0] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[1] ),
    .B1(n2413),
    .C1(n3793),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_N31));
 sky130_fd_sc_hd__inv_2 U2689 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_usb_reset_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2738));
 sky130_fd_sc_hd__a32o_1 U2690 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ),
    .A2(n2738),
    .A3(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q),
    .B1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_usb_reset_q),
    .B2(n3465),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(inst_to_wrap_u_usb_cdc_u_ctrl_endp_N109));
 sky130_fd_sc_hd__nor2_1 U2691 (.A(n2567),
    .B(n2565),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3836));
 sky130_fd_sc_hd__inv_2 U2692 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3715));
 sky130_fd_sc_hd__nor2_1 U2693 (.A(n2908),
    .B(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(inst_to_wrap_u_usb_cdc_ctrl_in_req));
 sky130_fd_sc_hd__a22o_1 U2694 (.A1(\inst_to_wrap_rx_fifo_array_reg[120] ),
    .A2(n2479),
    .B1(\inst_to_wrap_rx_fifo_array_reg[24] ),
    .B2(n2478),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2424));
 sky130_fd_sc_hd__a22o_1 U2695 (.A1(\inst_to_wrap_rx_fifo_array_reg[56] ),
    .A2(net207),
    .B1(\inst_to_wrap_rx_fifo_array_reg[72] ),
    .B2(n2480),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2417));
 sky130_fd_sc_hd__a22o_1 U2696 (.A1(\inst_to_wrap_rx_fifo_array_reg[104] ),
    .A2(n2483),
    .B1(\inst_to_wrap_rx_fifo_array_reg[88] ),
    .B2(n2482),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2416));
 sky130_fd_sc_hd__a22o_1 U2697 (.A1(\inst_to_wrap_rx_fifo_array_reg[40] ),
    .A2(n2485),
    .B1(\inst_to_wrap_rx_fifo_array_reg[8] ),
    .B2(n2484),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2415));
 sky130_fd_sc_hd__or4_1 U2698 (.A(n2417),
    .B(n2416),
    .C(n3559),
    .D(n2415),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2423));
 sky130_fd_sc_hd__a22o_1 U2699 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[112] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2422));
 sky130_fd_sc_hd__a22o_1 U2700 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[48] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2420));
 sky130_fd_sc_hd__a22o_1 U2701 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[96] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2419));
 sky130_fd_sc_hd__a22o_1 U2702 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[32] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2418));
 sky130_fd_sc_hd__or4_1 U2703 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2420),
    .C(n2419),
    .D(n2418),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2421));
 sky130_fd_sc_hd__o22a_1 U2704 (.A1(n2424),
    .A2(n2423),
    .B1(n2422),
    .B2(n2421),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2435));
 sky130_fd_sc_hd__a32o_1 U2705 (.A1(\RIS_REG[0] ),
    .A2(\IM_REG[0] ),
    .A3(n3709),
    .B1(\RIS_REG[0] ),
    .B2(n2460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2434));
 sky130_fd_sc_hd__inv_2 U2706 (.A(\TXFIFOLEVEL_REG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3143));
 sky130_fd_sc_hd__a31o_1 U2707 (.A1(\last_HADDR[4] ),
    .A2(\last_HADDR[3] ),
    .A3(CONTROL_REG_0_),
    .B1(n2426),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2432));
 sky130_fd_sc_hd__inv_2 U2708 (.A(n2427),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3712));
 sky130_fd_sc_hd__a22o_1 U2709 (.A1(n3712),
    .A2(CG_REG_0_),
    .B1(\rx_fifo_th[0] ),
    .B2(n3703),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2428));
 sky130_fd_sc_hd__a211o_1 U2710 (.A1(\RXFIFOLEVEL_REG[0] ),
    .A2(n2429),
    .B1(eco_net_9_0),
    .C1(n2428),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2431));
 sky130_fd_sc_hd__a22o_1 U2711 (.A1(\ICR_REG[0] ),
    .A2(n2495),
    .B1(\tx_fifo_th[0] ),
    .B2(n3700),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2430));
 sky130_fd_sc_hd__a211o_1 U2712 (.A1(n3708),
    .A2(n2432),
    .B1(n2431),
    .C1(n2430),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2433));
 sky130_fd_sc_hd__a211o_1 U2713 (.A1(n2494),
    .A2(n2435),
    .B1(n2434),
    .C1(n2433),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net));
 sky130_fd_sc_hd__a22o_1 U2714 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[124] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2445));
 sky130_fd_sc_hd__a22o_1 U2715 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[60] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2438));
 sky130_fd_sc_hd__a22o_1 U2716 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[108] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2437));
 sky130_fd_sc_hd__a22o_1 U2717 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[44] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2436));
 sky130_fd_sc_hd__or4_1 U2718 (.A(n3559),
    .B(n2438),
    .C(n2437),
    .D(n2436),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2444));
 sky130_fd_sc_hd__a22o_1 U2719 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[116] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2443));
 sky130_fd_sc_hd__a22o_1 U2720 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[52] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2441));
 sky130_fd_sc_hd__a22o_1 U2721 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[100] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2440));
 sky130_fd_sc_hd__a22o_1 U2722 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[36] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2439));
 sky130_fd_sc_hd__or4_1 U2723 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2441),
    .C(n2440),
    .D(n2439),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2442));
 sky130_fd_sc_hd__o22a_1 U2724 (.A1(n2445),
    .A2(n2444),
    .B1(n2443),
    .B2(n2442),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2448));
 sky130_fd_sc_hd__o211a_1 U2725 (.A1(\RIS_REG[4] ),
    .A2(n3708),
    .B1(n3709),
    .C1(\IM_REG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2447));
 sky130_fd_sc_hd__a22o_1 U2726 (.A1(n2460),
    .A2(\RIS_REG[4] ),
    .B1(n2495),
    .B2(\ICR_REG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2446));
 sky130_fd_sc_hd__a211o_1 U2727 (.A1(n2448),
    .A2(n2494),
    .B1(n2447),
    .C1(n2446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_3_0));
 sky130_fd_sc_hd__a22o_1 U2728 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[125] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2458));
 sky130_fd_sc_hd__a22o_1 U2729 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[61] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2451));
 sky130_fd_sc_hd__a22o_1 U2730 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[109] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2450));
 sky130_fd_sc_hd__a22o_1 U2731 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[45] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2449));
 sky130_fd_sc_hd__or4_1 U2732 (.A(n3559),
    .B(n2451),
    .C(n2450),
    .D(n2449),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2457));
 sky130_fd_sc_hd__a22o_1 U2733 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[117] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2456));
 sky130_fd_sc_hd__a22o_1 U2734 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[53] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2454));
 sky130_fd_sc_hd__a22o_1 U2735 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[101] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2453));
 sky130_fd_sc_hd__a22o_1 U2736 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[37] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2452));
 sky130_fd_sc_hd__or4_1 U2737 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2454),
    .C(n2453),
    .D(n2452),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2455));
 sky130_fd_sc_hd__o22a_1 U2738 (.A1(n2458),
    .A2(n2457),
    .B1(n2456),
    .B2(n2455),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2463));
 sky130_fd_sc_hd__or2_1 U2739 (.A(\RIS_REG[5] ),
    .B(n3708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2459));
 sky130_fd_sc_hd__a31o_1 U2740 (.A1(n3709),
    .A2(\IM_REG[5] ),
    .A3(n2459),
    .B1(eco_net_9_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2462));
 sky130_fd_sc_hd__a22o_1 U2741 (.A1(n2460),
    .A2(\RIS_REG[5] ),
    .B1(n2495),
    .B2(\ICR_REG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2461));
 sky130_fd_sc_hd__a211o_1 U2742 (.A1(n2494),
    .A2(n2463),
    .B1(n2462),
    .C1(n2461),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_4_0));
 sky130_fd_sc_hd__a22o_1 U2743 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[126] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2473));
 sky130_fd_sc_hd__a22o_1 U2744 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[62] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2466));
 sky130_fd_sc_hd__a22o_1 U2745 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[110] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2465));
 sky130_fd_sc_hd__a22o_1 U2746 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[46] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2464));
 sky130_fd_sc_hd__or4_1 U2747 (.A(n3559),
    .B(n2466),
    .C(n2465),
    .D(n2464),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2472));
 sky130_fd_sc_hd__a22o_1 U2748 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[118] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2471));
 sky130_fd_sc_hd__a22o_1 U2749 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[54] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2469));
 sky130_fd_sc_hd__a22o_1 U2750 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[102] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2468));
 sky130_fd_sc_hd__a22o_1 U2751 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[38] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2467));
 sky130_fd_sc_hd__or4_1 U2752 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2469),
    .C(n2468),
    .D(n2467),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2470));
 sky130_fd_sc_hd__o22a_1 U2753 (.A1(n2473),
    .A2(n2472),
    .B1(n2471),
    .B2(n2470),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2474));
 sky130_fd_sc_hd__a21o_1 U2754 (.A1(n2494),
    .A2(n2474),
    .B1(eco_net_9_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_5_0));
 sky130_fd_sc_hd__a22o_1 U2755 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[127] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2492));
 sky130_fd_sc_hd__a22o_1 U2756 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[63] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2477));
 sky130_fd_sc_hd__a22o_1 U2757 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[111] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2476));
 sky130_fd_sc_hd__a22o_1 U2758 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[47] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2475));
 sky130_fd_sc_hd__or4_1 U2759 (.A(n3559),
    .B(n2477),
    .C(n2476),
    .D(n2475),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2491));
 sky130_fd_sc_hd__a22o_1 U2760 (.A1(n2479),
    .A2(\inst_to_wrap_rx_fifo_array_reg[119] ),
    .B1(n2478),
    .B2(\inst_to_wrap_rx_fifo_array_reg[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2490));
 sky130_fd_sc_hd__a22o_1 U2761 (.A1(net207),
    .A2(\inst_to_wrap_rx_fifo_array_reg[55] ),
    .B1(n2480),
    .B2(\inst_to_wrap_rx_fifo_array_reg[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2488));
 sky130_fd_sc_hd__a22o_1 U2762 (.A1(n2483),
    .A2(\inst_to_wrap_rx_fifo_array_reg[103] ),
    .B1(n2482),
    .B2(\inst_to_wrap_rx_fifo_array_reg[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2487));
 sky130_fd_sc_hd__a22o_1 U2763 (.A1(n2485),
    .A2(\inst_to_wrap_rx_fifo_array_reg[39] ),
    .B1(n2484),
    .B2(\inst_to_wrap_rx_fifo_array_reg[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2486));
 sky130_fd_sc_hd__or4_1 U2764 (.A(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B(n2488),
    .C(n2487),
    .D(n2486),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2489));
 sky130_fd_sc_hd__o22a_1 U2765 (.A1(n2492),
    .A2(n2491),
    .B1(n2490),
    .B2(n2489),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2493));
 sky130_fd_sc_hd__a21o_1 U2766 (.A1(n2494),
    .A2(n2493),
    .B1(eco_net_9_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(eco_net_6_0));
 sky130_fd_sc_hd__and3_2 U2767 (.A(last_HTRANS_1_),
    .B(last_HSEL),
    .C(last_HWRITE),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3713));
 sky130_fd_sc_hd__nand2_2 U2768 (.A(n3713),
    .B(n2495),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2496));
 sky130_fd_sc_hd__nor2b_1 U2769 (.A(n2496),
    .B_N(net237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(N26));
 sky130_fd_sc_hd__nor2b_1 U2770 (.A(n2496),
    .B_N(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(N27));
 sky130_fd_sc_hd__nor2b_1 U2771 (.A(n2496),
    .B_N(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(N28));
 sky130_fd_sc_hd__nor2b_1 U2772 (.A(n2496),
    .B_N(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(N29));
 sky130_fd_sc_hd__nor2b_1 U2773 (.A(n2496),
    .B_N(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(N30));
 sky130_fd_sc_hd__nor2b_1 U2774 (.A(n2496),
    .B_N(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(N31));
 sky130_fd_sc_hd__inv_2 U2775 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3746));
 sky130_fd_sc_hd__nand2_2 U2776 (.A(n3746),
    .B(n3752),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3756));
 sky130_fd_sc_hd__inv_2 U2777 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2532));
 sky130_fd_sc_hd__o221a_1 U2778 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ),
    .A2(n3756),
    .B1(n2532),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[2] ),
    .C1(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2497));
 sky130_fd_sc_hd__a31o_2 U2779 (.A1(n2497),
    .A2(n3746),
    .A3(n3752),
    .B1(n3826),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2542));
 sky130_fd_sc_hd__inv_2 U2780 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2543));
 sky130_fd_sc_hd__or2_4 U2781 (.A(n2497),
    .B(n3826),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2530));
 sky130_fd_sc_hd__inv_2 U2782 (.A(n2530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2546));
 sky130_fd_sc_hd__a22o_1 U2783 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[0] ),
    .A2(n2542),
    .B1(n2543),
    .B2(n2546),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2269));
 sky130_fd_sc_hd__inv_1 U2784 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2499));
 sky130_fd_sc_hd__and4_1 U2785 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[3] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[1] ),
    .D(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2534));
 sky130_fd_sc_hd__and3_1 U2786 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[4] ),
    .C(n2534),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2527));
 sky130_fd_sc_hd__and3_1 U2787 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[6] ),
    .B(n2527),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2522));
 sky130_fd_sc_hd__and3_1 U2788 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[9] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[8] ),
    .C(n2522),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2517));
 sky130_fd_sc_hd__and3_1 U2789 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[10] ),
    .B(n2517),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2512));
 sky130_fd_sc_hd__and3_1 U2790 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[12] ),
    .B(n2512),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2507));
 sky130_fd_sc_hd__and3_1 U2791 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[14] ),
    .B(n2507),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2502));
 sky130_fd_sc_hd__nand2_1 U2792 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[16] ),
    .B(n2502),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2498));
 sky130_fd_sc_hd__mux2_1 U2793 (.A0(n2499),
    .A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[17] ),
    .S(n2498),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2500));
 sky130_fd_sc_hd__a22o_1 U2794 (.A1(n2546),
    .A2(n2500),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[17] ),
    .B2(n2542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2268));
 sky130_fd_sc_hd__inv_1 U2795 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2503));
 sky130_fd_sc_hd__inv_2 U2796 (.A(n2542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2529));
 sky130_fd_sc_hd__o21ai_1 U2797 (.A1(n2502),
    .A2(n2530),
    .B1(n2529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2501));
 sky130_fd_sc_hd__a32o_1 U2798 (.A1(n2546),
    .A2(n2503),
    .A3(n2502),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[16] ),
    .B2(n2501),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2267));
 sky130_fd_sc_hd__nor2_1 U2799 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[14] ),
    .B(n2530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2506));
 sky130_fd_sc_hd__o21ai_1 U2800 (.A1(n2507),
    .A2(n2530),
    .B1(n2529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2508));
 sky130_fd_sc_hd__inv_1 U2801 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2505));
 sky130_fd_sc_hd__and3_1 U2802 (.A(n2546),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[14] ),
    .C(n2507),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2504));
 sky130_fd_sc_hd__o32a_1 U2803 (.A1(n2506),
    .A2(n2508),
    .A3(n2505),
    .B1(n2504),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2266));
 sky130_fd_sc_hd__a22o_1 U2804 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[14] ),
    .A2(n2508),
    .B1(n2507),
    .B2(n2506),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2265));
 sky130_fd_sc_hd__nor2_1 U2805 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[12] ),
    .B(n2530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2511));
 sky130_fd_sc_hd__o21ai_1 U2806 (.A1(n2512),
    .A2(n2530),
    .B1(n2529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2513));
 sky130_fd_sc_hd__inv_1 U2807 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2510));
 sky130_fd_sc_hd__and3_1 U2808 (.A(n2546),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[12] ),
    .C(n2512),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2509));
 sky130_fd_sc_hd__o32a_1 U2809 (.A1(n2511),
    .A2(n2513),
    .A3(n2510),
    .B1(n2509),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2264));
 sky130_fd_sc_hd__a22o_1 U2810 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[12] ),
    .A2(n2513),
    .B1(n2512),
    .B2(n2511),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2263));
 sky130_fd_sc_hd__nor2_1 U2811 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[10] ),
    .B(n2530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2516));
 sky130_fd_sc_hd__o21ai_1 U2812 (.A1(n2517),
    .A2(n2530),
    .B1(n2529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2518));
 sky130_fd_sc_hd__inv_1 U2813 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2515));
 sky130_fd_sc_hd__and3_1 U2814 (.A(n2546),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[10] ),
    .C(n2517),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2514));
 sky130_fd_sc_hd__o32a_1 U2815 (.A1(n2516),
    .A2(n2518),
    .A3(n2515),
    .B1(n2514),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2262));
 sky130_fd_sc_hd__a22o_1 U2816 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[10] ),
    .A2(n2518),
    .B1(n2517),
    .B2(n2516),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2261));
 sky130_fd_sc_hd__nor2_1 U2817 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[8] ),
    .B(n2530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2521));
 sky130_fd_sc_hd__o21ai_1 U2818 (.A1(n2522),
    .A2(n2530),
    .B1(n2529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2523));
 sky130_fd_sc_hd__inv_1 U2819 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2520));
 sky130_fd_sc_hd__and3_1 U2820 (.A(n2546),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[8] ),
    .C(n2522),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2519));
 sky130_fd_sc_hd__o32a_1 U2821 (.A1(n2521),
    .A2(n2523),
    .A3(n2520),
    .B1(n2519),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2260));
 sky130_fd_sc_hd__a22o_1 U2822 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[8] ),
    .A2(n2523),
    .B1(n2522),
    .B2(n2521),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2259));
 sky130_fd_sc_hd__nor2_1 U2823 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[6] ),
    .B(n2530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2526));
 sky130_fd_sc_hd__o21ai_1 U2824 (.A1(n2527),
    .A2(n2530),
    .B1(n2529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2528));
 sky130_fd_sc_hd__inv_1 U2825 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2525));
 sky130_fd_sc_hd__and3_1 U2826 (.A(n2546),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[6] ),
    .C(n2527),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2524));
 sky130_fd_sc_hd__o32a_1 U2827 (.A1(n2526),
    .A2(n2528),
    .A3(n2525),
    .B1(n2524),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2258));
 sky130_fd_sc_hd__a22o_1 U2828 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[6] ),
    .A2(n2528),
    .B1(n2527),
    .B2(n2526),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2257));
 sky130_fd_sc_hd__nor2_1 U2829 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[4] ),
    .B(n2530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2533));
 sky130_fd_sc_hd__o21ai_1 U2830 (.A1(n2534),
    .A2(n2530),
    .B1(n2529),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2535));
 sky130_fd_sc_hd__and3_1 U2831 (.A(n2546),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[4] ),
    .C(n2534),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2531));
 sky130_fd_sc_hd__o32a_1 U2832 (.A1(n2533),
    .A2(n2535),
    .A3(n2532),
    .B1(n2531),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2256));
 sky130_fd_sc_hd__a22o_1 U2833 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[4] ),
    .A2(n2535),
    .B1(n2534),
    .B2(n2533),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2255));
 sky130_fd_sc_hd__inv_1 U2834 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2538));
 sky130_fd_sc_hd__and3_1 U2835 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2537));
 sky130_fd_sc_hd__inv_2 U2836 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2541));
 sky130_fd_sc_hd__inv_2 U2837 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2545));
 sky130_fd_sc_hd__o32a_1 U2838 (.A1(n2542),
    .A2(n2545),
    .A3(n2543),
    .B1(n2542),
    .B2(n2546),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2539));
 sky130_fd_sc_hd__a21o_1 U2839 (.A1(n2541),
    .A2(n2546),
    .B1(n2539),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2536));
 sky130_fd_sc_hd__a32o_1 U2840 (.A1(n2546),
    .A2(n2538),
    .A3(n2537),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[3] ),
    .B2(n2536),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2254));
 sky130_fd_sc_hd__nor2_1 U2841 (.A(n2545),
    .B(n2543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2540));
 sky130_fd_sc_hd__a32o_1 U2842 (.A1(n2546),
    .A2(n2541),
    .A3(n2540),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[2] ),
    .B2(n2539),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2253));
 sky130_fd_sc_hd__a21o_1 U2843 (.A1(n2543),
    .A2(n2546),
    .B1(n2542),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2544));
 sky130_fd_sc_hd__a32o_1 U2844 (.A1(n2546),
    .A2(n2545),
    .A3(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[0] ),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[1] ),
    .B2(n2544),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2252));
 sky130_fd_sc_hd__a31o_1 U2845 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[9] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[8] ),
    .A3(n2547),
    .B1(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2251));
 sky130_fd_sc_hd__or4b_4 U2846 (.A(n_TX_FULL_FLAG_FLAG_),
    .B(\last_HADDR[4] ),
    .C(\last_HADDR[3] ),
    .D_N(n3706),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3194));
 sky130_fd_sc_hd__inv_2 U2847 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3183));
 sky130_fd_sc_hd__inv_2 U2848 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3193));
 sky130_fd_sc_hd__or3_2 U2849 (.A(n3194),
    .B(n3183),
    .C(n3193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3208));
 sky130_fd_sc_hd__clkinv_2 U2850 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3190));
 sky130_fd_sc_hd__or3b_4 U2851 (.A(n3208),
    .B(n3190),
    .C_N(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3215));
 sky130_fd_sc_hd__clkinv_2 U2852 (.A(n3215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3216));
 sky130_fd_sc_hd__a22o_1 U2853 (.A1(n3216),
    .A2(net27),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2249));
 sky130_fd_sc_hd__or3b_1 U2854 (.A(n_TX_EMPTY_FLAG_FLAG_),
    .B(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_mask_q),
    .C_N(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3301));
 sky130_fd_sc_hd__inv_2 U2855 (.A(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3304));
 sky130_fd_sc_hd__clkinv_2 U2856 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3158));
 sky130_fd_sc_hd__inv_2 U2857 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3127));
 sky130_fd_sc_hd__clkinv_2 U2858 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3157));
 sky130_fd_sc_hd__and3_4 U2859 (.A(n3158),
    .B(n3127),
    .C(n3157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3288));
 sky130_fd_sc_hd__and3_4 U2860 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ),
    .B(n3158),
    .C(n3127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3287));
 sky130_fd_sc_hd__a22o_1 U2861 (.A1(\inst_to_wrap_tx_fifo_array_reg[15] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[47] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2552));
 sky130_fd_sc_hd__and3_4 U2862 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ),
    .B(n3127),
    .C(n3157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3290));
 sky130_fd_sc_hd__and3_1 U2863 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ),
    .B(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ),
    .C(n3127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3289));
 sky130_fd_sc_hd__a22o_1 U2864 (.A1(\inst_to_wrap_tx_fifo_array_reg[31] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[63] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2551));
 sky130_fd_sc_hd__and3_4 U2865 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ),
    .B(n3158),
    .C(n3157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3292));
 sky130_fd_sc_hd__and3_4 U2866 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ),
    .B(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ),
    .C(n3158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3291));
 sky130_fd_sc_hd__a22o_1 U2867 (.A1(\inst_to_wrap_tx_fifo_array_reg[79] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[111] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2550));
 sky130_fd_sc_hd__and3_4 U2868 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ),
    .B(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ),
    .C(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3293));
 sky130_fd_sc_hd__and3_4 U2869 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ),
    .B(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ),
    .C(n3157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3294));
 sky130_fd_sc_hd__a22o_1 U2870 (.A1(\inst_to_wrap_tx_fifo_array_reg[127] ),
    .A2(n3293),
    .B1(\inst_to_wrap_tx_fifo_array_reg[95] ),
    .B2(n3294),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2549));
 sky130_fd_sc_hd__or4_1 U2871 (.A(n2552),
    .B(n2551),
    .C(n2550),
    .D(n2549),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2559));
 sky130_fd_sc_hd__nor2_2 U2872 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .B(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3300));
 sky130_fd_sc_hd__a22o_1 U2873 (.A1(\inst_to_wrap_tx_fifo_array_reg[7] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[39] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2556));
 sky130_fd_sc_hd__a22o_1 U2874 (.A1(\inst_to_wrap_tx_fifo_array_reg[23] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[55] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2555));
 sky130_fd_sc_hd__a22o_1 U2875 (.A1(\inst_to_wrap_tx_fifo_array_reg[71] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[103] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2554));
 sky130_fd_sc_hd__a22o_1 U2876 (.A1(\inst_to_wrap_tx_fifo_array_reg[87] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[119] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2553));
 sky130_fd_sc_hd__or4_1 U2877 (.A(n2556),
    .B(n2555),
    .C(n2554),
    .D(n2553),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2557));
 sky130_fd_sc_hd__a22o_1 U2878 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[7] ),
    .A2(net209),
    .B1(n3300),
    .B2(n2557),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2558));
 sky130_fd_sc_hd__a31o_1 U2879 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n2559),
    .B1(n2558),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2248));
 sky130_fd_sc_hd__or2_4 U2880 (.A(n3116),
    .B(n3121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3321));
 sky130_fd_sc_hd__clkinv_2 U2881 (.A(n3321),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3322));
 sky130_fd_sc_hd__a22o_1 U2882 (.A1(n3322),
    .A2(net91),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2247));
 sky130_fd_sc_hd__nand2_1 U2883 (.A(n2575),
    .B(n3722),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2582));
 sky130_fd_sc_hd__nor2_1 U2884 (.A(n2626),
    .B(n2582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3835));
 sky130_fd_sc_hd__nor2_1 U2885 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[0] ),
    .B(n2626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2580));
 sky130_fd_sc_hd__inv_2 U2886 (.A(n2580),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2579));
 sky130_fd_sc_hd__or2_1 U2887 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[1] ),
    .B(n2579),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2560));
 sky130_fd_sc_hd__inv_2 U2888 (.A(n2560),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2578));
 sky130_fd_sc_hd__inv_1 U2889 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2561));
 sky130_fd_sc_hd__a32o_1 U2890 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ),
    .A2(n2578),
    .A3(n2561),
    .B1(n2560),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2563));
 sky130_fd_sc_hd__or3b_1 U2891 (.A(n3835),
    .B(n2563),
    .C_N(n2562),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2246));
 sky130_fd_sc_hd__o21ai_1 U2892 (.A1(n3716),
    .A2(n2575),
    .B1(n2581),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2585));
 sky130_fd_sc_hd__inv_2 U2893 (.A(n2583),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3717));
 sky130_fd_sc_hd__inv_2 U2894 (.A(n2626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3837));
 sky130_fd_sc_hd__o211a_1 U2895 (.A1(n2575),
    .A2(n2581),
    .B1(n3837),
    .C1(n2582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2566));
 sky130_fd_sc_hd__nand2_1 U2896 (.A(n3717),
    .B(n2566),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2564));
 sky130_fd_sc_hd__mux2_1 U2897 (.A0(n2585),
    .A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[1] ),
    .S(n2564),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2245));
 sky130_fd_sc_hd__o211a_1 U2898 (.A1(n3717),
    .A2(n2567),
    .B1(n2566),
    .C1(n2565),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2568));
 sky130_fd_sc_hd__a21o_1 U2899 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ),
    .A2(n3830),
    .B1(n2568),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2244));
 sky130_fd_sc_hd__or4_4 U2900 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ),
    .C(n2820),
    .D(n3079),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2740));
 sky130_fd_sc_hd__or4_4 U2901 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .B(n2820),
    .C(n3079),
    .D(n2744),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2618));
 sky130_fd_sc_hd__o22a_1 U2902 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[0] ),
    .A2(n2618),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ),
    .B2(n2617),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2571));
 sky130_fd_sc_hd__clkinv_2 U2903 (.A(n3047),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3037));
 sky130_fd_sc_hd__o22a_1 U2904 (.A1(n3070),
    .A2(n2644),
    .B1(n3037),
    .B2(n2569),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2570));
 sky130_fd_sc_hd__o211a_1 U2905 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[8] ),
    .A2(n2740),
    .B1(n2571),
    .C1(n2570),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2573));
 sky130_fd_sc_hd__nor2_1 U2906 (.A(n2573),
    .B(n2572),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2576));
 sky130_fd_sc_hd__inv_1 U2907 (.A(n3830),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2574));
 sky130_fd_sc_hd__o31a_1 U2908 (.A1(n3836),
    .A2(n2576),
    .A3(n2575),
    .B1(n2574),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2577));
 sky130_fd_sc_hd__a211o_1 U2909 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[7] ),
    .A2(n2626),
    .B1(n3835),
    .C1(n2577),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2243));
 sky130_fd_sc_hd__a211o_1 U2910 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[1] ),
    .A2(n2579),
    .B1(n3835),
    .C1(n2578),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2242));
 sky130_fd_sc_hd__a211o_1 U2911 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[0] ),
    .A2(n2626),
    .B1(n2580),
    .C1(n3835),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2241));
 sky130_fd_sc_hd__nor3_2 U2912 (.A(n3830),
    .B(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q),
    .C(n2581),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2625));
 sky130_fd_sc_hd__o211a_2 U2913 (.A1(n3722),
    .A2(n2583),
    .B1(n3837),
    .C1(n2582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2621));
 sky130_fd_sc_hd__a22o_1 U2914 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[1] ),
    .A2(n2621),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[0] ),
    .B2(n2626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2589));
 sky130_fd_sc_hd__o22a_1 U2915 (.A1(n2584),
    .A2(n2617),
    .B1(n3070),
    .B2(n3049),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2587));
 sky130_fd_sc_hd__o22a_1 U2916 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[15] ),
    .A2(n2740),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[7] ),
    .B2(n2618),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2586));
 sky130_fd_sc_hd__inv_2 U2917 (.A(n2585),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3718));
 sky130_fd_sc_hd__or3_2 U2918 (.A(n3089),
    .B(n3718),
    .C(n3830),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2622));
 sky130_fd_sc_hd__a31o_1 U2919 (.A1(n2587),
    .A2(n2586),
    .A3(n3072),
    .B1(n2622),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2588));
 sky130_fd_sc_hd__or3b_1 U2920 (.A(n2625),
    .B(n2589),
    .C_N(n2588),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2240));
 sky130_fd_sc_hd__o22a_1 U2921 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[6] ),
    .A2(n2618),
    .B1(n3070),
    .B2(n3050),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2590));
 sky130_fd_sc_hd__o21ai_1 U2922 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[14] ),
    .A2(n2740),
    .B1(n2590),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2591));
 sky130_fd_sc_hd__a211o_1 U2923 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[1] ),
    .A2(n2592),
    .B1(n3047),
    .C1(n2591),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2594));
 sky130_fd_sc_hd__a22o_1 U2924 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[2] ),
    .A2(n2621),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[1] ),
    .B2(n2626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2593));
 sky130_fd_sc_hd__a21o_1 U2925 (.A1(n2595),
    .A2(n2594),
    .B1(n2593),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2239));
 sky130_fd_sc_hd__inv_2 U2926 (.A(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3059));
 sky130_fd_sc_hd__o22a_1 U2927 (.A1(n3059),
    .A2(n2617),
    .B1(n3070),
    .B2(n3065),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2598));
 sky130_fd_sc_hd__o22a_1 U2928 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[5] ),
    .A2(n2618),
    .B1(n3037),
    .B2(n2596),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2597));
 sky130_fd_sc_hd__o211a_1 U2929 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[13] ),
    .A2(n2740),
    .B1(n2598),
    .C1(n2597),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2600));
 sky130_fd_sc_hd__a21o_1 U2930 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[2] ),
    .A2(n2626),
    .B1(n2601),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2238));
 sky130_fd_sc_hd__a22o_1 U2931 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[4] ),
    .A2(n2621),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[3] ),
    .B2(n2626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2606));
 sky130_fd_sc_hd__inv_2 U2932 (.A(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3058));
 sky130_fd_sc_hd__o22a_1 U2933 (.A1(n3058),
    .A2(n2617),
    .B1(n3070),
    .B2(n2803),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2604));
 sky130_fd_sc_hd__o22a_1 U2934 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[12] ),
    .A2(n2740),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[4] ),
    .B2(n2618),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2603));
 sky130_fd_sc_hd__a31o_1 U2935 (.A1(n2604),
    .A2(n2603),
    .A3(n2602),
    .B1(n2622),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2605));
 sky130_fd_sc_hd__or3b_1 U2936 (.A(n2625),
    .B(n2606),
    .C_N(n2605),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2237));
 sky130_fd_sc_hd__o22a_1 U2937 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[0] ),
    .A2(n2617),
    .B1(n2639),
    .B2(n3070),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2608));
 sky130_fd_sc_hd__o22a_1 U2938 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[11] ),
    .A2(n2740),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[3] ),
    .B2(n2618),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2607));
 sky130_fd_sc_hd__o211a_1 U2939 (.A1(n3046),
    .A2(n3037),
    .B1(n2608),
    .C1(n2607),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2609));
 sky130_fd_sc_hd__a2bb2o_1 U2940 (.A1_N(n2609),
    .A2_N(n2622),
    .B1(n2621),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2610));
 sky130_fd_sc_hd__a211o_1 U2941 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[4] ),
    .A2(n2626),
    .B1(n2625),
    .C1(n2610),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2236));
 sky130_fd_sc_hd__o22a_1 U2942 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[1] ),
    .A2(n2617),
    .B1(n2611),
    .B2(n3070),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2613));
 sky130_fd_sc_hd__o22a_1 U2943 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[10] ),
    .A2(n2740),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[2] ),
    .B2(n2618),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2612));
 sky130_fd_sc_hd__a21oi_1 U2944 (.A1(n2613),
    .A2(n2612),
    .B1(n2622),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2615));
 sky130_fd_sc_hd__a22o_1 U2945 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[6] ),
    .A2(n2621),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[5] ),
    .B2(n2626),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2614));
 sky130_fd_sc_hd__or3_1 U2946 (.A(n2625),
    .B(n2615),
    .C(n2614),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2235));
 sky130_fd_sc_hd__o22a_1 U2947 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[2] ),
    .A2(n2617),
    .B1(n2616),
    .B2(n3070),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2620));
 sky130_fd_sc_hd__o22a_1 U2948 (.A1(n3038),
    .A2(n3037),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[1] ),
    .B2(n2618),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2619));
 sky130_fd_sc_hd__o211a_1 U2949 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[9] ),
    .A2(n2740),
    .B1(n2620),
    .C1(n2619),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2623));
 sky130_fd_sc_hd__a211o_1 U2950 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[6] ),
    .A2(n2626),
    .B1(n2625),
    .C1(n2624),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2234));
 sky130_fd_sc_hd__inv_2 U2951 (.A(\inst_to_wrap_u_usb_cdc_addr[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2792));
 sky130_fd_sc_hd__inv_1 U2952 (.A(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2634));
 sky130_fd_sc_hd__clkinv_2 U2953 (.A(net213),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3428));
 sky130_fd_sc_hd__inv_2 U2954 (.A(\inst_to_wrap_u_usb_cdc_addr[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2798));
 sky130_fd_sc_hd__inv_2 U2955 (.A(\inst_to_wrap_u_usb_cdc_addr[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2795));
 sky130_fd_sc_hd__a22o_1 U2956 (.A1(\inst_to_wrap_u_usb_cdc_out_data[2] ),
    .A2(\inst_to_wrap_u_usb_cdc_addr[2] ),
    .B1(n3405),
    .B2(n2795),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2627));
 sky130_fd_sc_hd__o221a_1 U2957 (.A1(\inst_to_wrap_u_usb_cdc_addr[0] ),
    .A2(n3428),
    .B1(n2798),
    .B2(net213),
    .C1(n2627),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2632));
 sky130_fd_sc_hd__inv_2 U2958 (.A(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3378));
 sky130_fd_sc_hd__inv_2 U2959 (.A(\inst_to_wrap_u_usb_cdc_addr[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2794));
 sky130_fd_sc_hd__inv_2 U2960 (.A(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2635));
 sky130_fd_sc_hd__inv_2 U2961 (.A(\inst_to_wrap_u_usb_cdc_addr[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2788));
 sky130_fd_sc_hd__a22o_1 U2962 (.A1(net215),
    .A2(\inst_to_wrap_u_usb_cdc_addr[6] ),
    .B1(n2635),
    .B2(n2788),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2628));
 sky130_fd_sc_hd__o221a_1 U2963 (.A1(\inst_to_wrap_u_usb_cdc_addr[3] ),
    .A2(n3378),
    .B1(n2794),
    .B2(net218),
    .C1(n2628),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2631));
 sky130_fd_sc_hd__inv_2 U2964 (.A(net211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2712));
 sky130_fd_sc_hd__inv_2 U2965 (.A(\inst_to_wrap_u_usb_cdc_addr[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2797));
 sky130_fd_sc_hd__inv_2 U2966 (.A(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3404));
 sky130_fd_sc_hd__inv_2 U2967 (.A(\inst_to_wrap_u_usb_cdc_addr[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2791));
 sky130_fd_sc_hd__a22o_1 U2968 (.A1(\inst_to_wrap_u_usb_cdc_out_data[5] ),
    .A2(\inst_to_wrap_u_usb_cdc_addr[5] ),
    .B1(n3404),
    .B2(n2791),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2629));
 sky130_fd_sc_hd__o221a_1 U2969 (.A1(\inst_to_wrap_u_usb_cdc_addr[1] ),
    .A2(n2712),
    .B1(n2797),
    .B2(net211),
    .C1(n2629),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2630));
 sky130_fd_sc_hd__and3_1 U2970 (.A(n2632),
    .B(n2631),
    .C(n2630),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2633));
 sky130_fd_sc_hd__o221a_1 U2971 (.A1(\inst_to_wrap_u_usb_cdc_out_data[4] ),
    .A2(n2792),
    .B1(n2634),
    .B2(\inst_to_wrap_u_usb_cdc_addr[4] ),
    .C1(n2633),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2818));
 sky130_fd_sc_hd__nand2_1 U2972 (.A(n3056),
    .B(n2772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3064));
 sky130_fd_sc_hd__nor2_1 U2973 (.A(\inst_to_wrap_u_usb_cdc_out_data[3] ),
    .B(\inst_to_wrap_u_usb_cdc_out_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2717));
 sky130_fd_sc_hd__inv_2 U2974 (.A(n2717),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3424));
 sky130_fd_sc_hd__o21a_1 U2975 (.A1(n3405),
    .A2(n3378),
    .B1(n3424),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2642));
 sky130_fd_sc_hd__inv_2 U2976 (.A(\inst_to_wrap_u_usb_cdc_out_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2693));
 sky130_fd_sc_hd__o22a_1 U2977 (.A1(n2693),
    .A2(net211),
    .B1(\inst_to_wrap_u_usb_cdc_out_data[7] ),
    .B2(n2712),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2646));
 sky130_fd_sc_hd__inv_2 U2978 (.A(n2646),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2637));
 sky130_fd_sc_hd__a22o_1 U2979 (.A1(net213),
    .A2(n2635),
    .B1(n3428),
    .B2(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2648));
 sky130_fd_sc_hd__mux2_1 U2980 (.A0(n3050),
    .A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .S(n2648),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2641));
 sky130_fd_sc_hd__inv_2 U2981 (.A(n2641),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2636));
 sky130_fd_sc_hd__fa_1 U2982 (.A(n2642),
    .B(n2637),
    .CIN(n2636),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2638));
 sky130_fd_sc_hd__mux2_1 U2983 (.A0(n2639),
    .A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[4] ),
    .S(n2638),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2640));
 sky130_fd_sc_hd__a31o_1 U2984 (.A1(n3060),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[2] ),
    .A3(n3058),
    .B1(n2640),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2657));
 sky130_fd_sc_hd__fa_1 U2985 (.A(\inst_to_wrap_u_usb_cdc_out_data[4] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_data_q[6] ),
    .CIN(n2641),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2645));
 sky130_fd_sc_hd__a22o_1 U2986 (.A1(\inst_to_wrap_u_usb_cdc_out_data[5] ),
    .A2(n3049),
    .B1(n3404),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2650));
 sky130_fd_sc_hd__fa_1 U2987 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[5] ),
    .B(n2642),
    .CIN(n2650),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2651));
 sky130_fd_sc_hd__nor2_1 U2988 (.A(\inst_to_wrap_u_usb_cdc_out_data[3] ),
    .B(n2645),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2643));
 sky130_fd_sc_hd__a221o_1 U2989 (.A1(n2645),
    .A2(net218),
    .B1(n2644),
    .B2(n2651),
    .C1(n2643),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2656));
 sky130_fd_sc_hd__fa_1 U2990 (.A(net213),
    .B(net217),
    .CIN(n2646),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2647));
 sky130_fd_sc_hd__fa_1 U2991 (.A(net216),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .CIN(n2647),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2654));
 sky130_fd_sc_hd__fa_1 U2992 (.A(net211),
    .B(net219),
    .CIN(n2648),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2649));
 sky130_fd_sc_hd__fa_1 U2993 (.A(\inst_to_wrap_u_usb_cdc_u_sie_data_q[3] ),
    .B(n2650),
    .CIN(n2649),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .SUM(n2653));
 sky130_fd_sc_hd__nor2_1 U2994 (.A(n2651),
    .B(n2654),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2652));
 sky130_fd_sc_hd__a211o_1 U2995 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ),
    .A2(n2654),
    .B1(n2653),
    .C1(n2652),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2655));
 sky130_fd_sc_hd__or4_1 U2996 (.A(n3051),
    .B(n2657),
    .C(n2656),
    .D(n2655),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2771));
 sky130_fd_sc_hd__or3_2 U2997 (.A(n3079),
    .B(n3064),
    .C(n2771),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3085));
 sky130_fd_sc_hd__nor2_4 U2998 (.A(n3074),
    .B(n3085),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3036));
 sky130_fd_sc_hd__and3_1 U2999 (.A(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ),
    .B(n3036),
    .C(n3059),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2660));
 sky130_fd_sc_hd__clkinv_2 U3000 (.A(n3029),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3080));
 sky130_fd_sc_hd__a31o_1 U3001 (.A1(n3070),
    .A2(n3072),
    .A3(n2740),
    .B1(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2658));
 sky130_fd_sc_hd__o21ai_1 U3002 (.A1(n3080),
    .A2(n2820),
    .B1(n2658),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2659));
 sky130_fd_sc_hd__a31o_1 U3003 (.A1(n3060),
    .A2(n2818),
    .A3(n2660),
    .B1(n2659),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2233));
 sky130_fd_sc_hd__nand2_1 U3004 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2742));
 sky130_fd_sc_hd__nand2_2 U3005 (.A(n2742),
    .B(n2772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3462));
 sky130_fd_sc_hd__o21a_1 U3006 (.A1(n2661),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[4] ),
    .B1(n3462),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2232));
 sky130_fd_sc_hd__inv_2 U3007 (.A(n3462),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3453));
 sky130_fd_sc_hd__nor2_1 U3008 (.A(n3453),
    .B(n3454),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3460));
 sky130_fd_sc_hd__inv_2 U3009 (.A(n3460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3093));
 sky130_fd_sc_hd__clkinv_2 U3010 (.A(n3051),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3068));
 sky130_fd_sc_hd__a22o_1 U3011 (.A1(n2806),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[1] ),
    .B1(n2814),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2764));
 sky130_fd_sc_hd__inv_2 U3012 (.A(n2764),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2763));
 sky130_fd_sc_hd__a221o_1 U3013 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ),
    .A2(n2763),
    .B1(n3058),
    .B2(n2764),
    .C1(n2662),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3086));
 sky130_fd_sc_hd__a221o_1 U3014 (.A1(n3068),
    .A2(n2663),
    .B1(n3068),
    .B2(n3086),
    .C1(n3089),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2664));
 sky130_fd_sc_hd__a22o_1 U3015 (.A1(inst_to_wrap_u_usb_cdc_out_err),
    .A2(n3093),
    .B1(n2664),
    .B2(n2779),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2231));
 sky130_fd_sc_hd__inv_1 U3016 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2666));
 sky130_fd_sc_hd__inv_2 U3017 (.A(inst_to_wrap_u_usb_cdc_in_data_ack),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3344));
 sky130_fd_sc_hd__or2_1 U3018 (.A(n3344),
    .B(n3499),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2680));
 sky130_fd_sc_hd__o21ai_1 U3019 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ),
    .A2(n3477),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3464));
 sky130_fd_sc_hd__a22o_1 U3020 (.A1(inst_to_wrap_u_usb_cdc_out_err),
    .A2(n2697),
    .B1(n3351),
    .B2(n3464),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2665));
 sky130_fd_sc_hd__a31o_1 U3021 (.A1(n2667),
    .A2(n2666),
    .A3(n2680),
    .B1(n2665),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2668));
 sky130_fd_sc_hd__or2_1 U3022 (.A(n3465),
    .B(n2668),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2676));
 sky130_fd_sc_hd__inv_2 U3023 (.A(n2676),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3355));
 sky130_fd_sc_hd__inv_2 U3024 (.A(inst_to_wrap_u_usb_cdc_out_err),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3475));
 sky130_fd_sc_hd__a31o_1 U3025 (.A1(n3349),
    .A2(n2672),
    .A3(n2671),
    .B1(n3350),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2675));
 sky130_fd_sc_hd__inv_2 U3026 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3345));
 sky130_fd_sc_hd__or4_1 U3027 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q),
    .B(n3345),
    .C(n2673),
    .D(n2680),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2674));
 sky130_fd_sc_hd__or3b_1 U3028 (.A(n3057),
    .B(n2675),
    .C_N(n2674),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2677));
 sky130_fd_sc_hd__a32o_1 U3029 (.A1(n3355),
    .A2(n3475),
    .A3(n2677),
    .B1(n2676),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2230));
 sky130_fd_sc_hd__nand2_1 U3030 (.A(n3477),
    .B(n3349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2678));
 sky130_fd_sc_hd__o32a_1 U3031 (.A1(n3465),
    .A2(n3466),
    .A3(n2678),
    .B1(n3465),
    .B2(n2738),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2736));
 sky130_fd_sc_hd__inv_2 U3032 (.A(n2736),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2739));
 sky130_fd_sc_hd__nor2_1 U3033 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2708));
 sky130_fd_sc_hd__inv_2 U3034 (.A(n2708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2760));
 sky130_fd_sc_hd__or2_1 U3035 (.A(n2786),
    .B(n2760),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3439));
 sky130_fd_sc_hd__o21a_1 U3036 (.A1(n3870),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[0] ),
    .B1(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net58));
 sky130_fd_sc_hd__or4b_1 U3037 (.A(\last_HADDR[4] ),
    .B(n2290),
    .C(n3871),
    .D_N(\last_HADDR[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2288));
 sky130_fd_sc_hd__or4_2 U3038 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(n3348),
    .C(n3439),
    .D(n2680),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3468));
 sky130_fd_sc_hd__or4_1 U3039 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[3] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[4] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[5] ),
    .D(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2681));
 sky130_fd_sc_hd__or4_1 U3040 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[2] ),
    .D(n2681),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2734));
 sky130_fd_sc_hd__nor2_1 U3041 (.A(n3468),
    .B(n2734),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2682));
 sky130_fd_sc_hd__a211o_1 U3042 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[0] ),
    .A2(n2732),
    .B1(n2682),
    .C1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_usb_reset_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2684));
 sky130_fd_sc_hd__or3_1 U3043 (.A(n3348),
    .B(n3439),
    .C(n3344),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3469));
 sky130_fd_sc_hd__or2_1 U3044 (.A(n2736),
    .B(n3469),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2683));
 sky130_fd_sc_hd__a22o_1 U3045 (.A1(n2739),
    .A2(n2684),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[0] ),
    .B2(n2683),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2229));
 sky130_fd_sc_hd__and3_2 U3046 (.A(n3361),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3433));
 sky130_fd_sc_hd__inv_2 U3047 (.A(n3433),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3397));
 sky130_fd_sc_hd__a211o_1 U3048 (.A1(n2786),
    .A2(n3397),
    .B1(n2760),
    .C1(n3010),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2690));
 sky130_fd_sc_hd__and3_1 U3049 (.A(n2685),
    .B(n2760),
    .C(n2687),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2686));
 sky130_fd_sc_hd__o22a_1 U3050 (.A1(n2686),
    .A2(n2962),
    .B1(n3010),
    .B2(n3361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2721));
 sky130_fd_sc_hd__inv_2 U3051 (.A(n2687),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2997));
 sky130_fd_sc_hd__nor2_1 U3052 (.A(n2885),
    .B(n2997),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2706));
 sky130_fd_sc_hd__nor2_1 U3053 (.A(n3010),
    .B(n2688),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3434));
 sky130_fd_sc_hd__inv_2 U3054 (.A(n3434),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3395));
 sky130_fd_sc_hd__o22a_1 U3055 (.A1(n3394),
    .A2(n2886),
    .B1(n2706),
    .B2(n3395),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2689));
 sky130_fd_sc_hd__or4_1 U3056 (.A(net214),
    .B(net216),
    .C(net217),
    .D(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3379));
 sky130_fd_sc_hd__or2_1 U3057 (.A(n3379),
    .B(n3424),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2702));
 sky130_fd_sc_hd__nor2_2 U3058 (.A(net211),
    .B(n2702),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3446));
 sky130_fd_sc_hd__nand2_1 U3059 (.A(n3428),
    .B(n3446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2730));
 sky130_fd_sc_hd__a31o_1 U3060 (.A1(n2690),
    .A2(n2721),
    .A3(n2689),
    .B1(n2730),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2701));
 sky130_fd_sc_hd__or2_1 U3061 (.A(n2760),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2723));
 sky130_fd_sc_hd__or2_1 U3062 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(n2723),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3410));
 sky130_fd_sc_hd__inv_2 U3063 (.A(n3410),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3384));
 sky130_fd_sc_hd__a211o_1 U3064 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .A2(n2760),
    .B1(n3387),
    .C1(n3384),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2696));
 sky130_fd_sc_hd__inv_1 U3065 (.A(n3439),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2694));
 sky130_fd_sc_hd__o21ai_1 U3066 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .B1(n2708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2691));
 sky130_fd_sc_hd__o211a_1 U3067 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .A2(n3394),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .C1(n2691),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2692));
 sky130_fd_sc_hd__a31o_1 U3068 (.A1(n3443),
    .A2(n2694),
    .A3(n2693),
    .B1(n2692),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2695));
 sky130_fd_sc_hd__a21oi_1 U3069 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .A2(n2696),
    .B1(n2695),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2700));
 sky130_fd_sc_hd__nor2_2 U3070 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2954));
 sky130_fd_sc_hd__inv_2 U3071 (.A(n2954),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2955));
 sky130_fd_sc_hd__or4_1 U3072 (.A(n3467),
    .B(n2697),
    .C(n2956),
    .D(n2955),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2698));
 sky130_fd_sc_hd__nand3_1 U3073 (.A(\last_HADDR[11] ),
    .B(\last_HADDR[10] ),
    .C(\last_HADDR[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3871));
 sky130_fd_sc_hd__inv_2 U3074 (.A(n3438),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3435));
 sky130_fd_sc_hd__or3_1 U3075 (.A(net213),
    .B(n2712),
    .C(n2702),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3388));
 sky130_fd_sc_hd__inv_2 U3076 (.A(n3446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3393));
 sky130_fd_sc_hd__nor2_1 U3077 (.A(n3428),
    .B(n3393),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3445));
 sky130_fd_sc_hd__inv_2 U3078 (.A(n3445),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3417));
 sky130_fd_sc_hd__a22o_1 U3079 (.A1(n3389),
    .A2(n3388),
    .B1(n2884),
    .B2(n3417),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2707));
 sky130_fd_sc_hd__inv_2 U3080 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2709));
 sky130_fd_sc_hd__o211a_1 U3081 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ),
    .A2(n3428),
    .B1(n3446),
    .C1(n2709),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3390));
 sky130_fd_sc_hd__inv_2 U3082 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2724));
 sky130_fd_sc_hd__or3_1 U3083 (.A(net217),
    .B(net215),
    .C(n3424),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3402));
 sky130_fd_sc_hd__a21oi_1 U3084 (.A1(net213),
    .A2(net211),
    .B1(n3402),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2722));
 sky130_fd_sc_hd__a31o_1 U3085 (.A1(\inst_to_wrap_u_usb_cdc_out_data[7] ),
    .A2(n2722),
    .A3(n3404),
    .B1(n3446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2703));
 sky130_fd_sc_hd__and3_1 U3086 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ),
    .B(n2724),
    .C(n2703),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3391));
 sky130_fd_sc_hd__a221o_1 U3087 (.A1(n2723),
    .A2(n3390),
    .B1(n2723),
    .B2(n2283),
    .C1(n3391),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2704));
 sky130_fd_sc_hd__o211a_1 U3088 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .A2(n3446),
    .B1(n2704),
    .C1(n3439),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2705));
 sky130_fd_sc_hd__a21oi_1 U3089 (.A1(n2706),
    .A2(n2705),
    .B1(n3395),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3432));
 sky130_fd_sc_hd__a221o_1 U3090 (.A1(n3433),
    .A2(n2708),
    .B1(n3433),
    .B2(n2707),
    .C1(n3432),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3415));
 sky130_fd_sc_hd__or2_1 U3091 (.A(n3345),
    .B(n2716),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3380));
 sky130_fd_sc_hd__or4_1 U3092 (.A(net211),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ),
    .D(n3380),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2711));
 sky130_fd_sc_hd__and3_1 U3093 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2995));
 sky130_fd_sc_hd__or2_1 U3094 (.A(n2285),
    .B(n2286),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2290));
 sky130_fd_sc_hd__and3_1 U3096 (.A(net218),
    .B(n2711),
    .C(n3377),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3409));
 sky130_fd_sc_hd__a22o_1 U3097 (.A1(n2717),
    .A2(n3428),
    .B1(net211),
    .B2(n3378),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3406));
 sky130_fd_sc_hd__inv_2 U3098 (.A(net219),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3405));
 sky130_fd_sc_hd__o211a_1 U3099 (.A1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .A2(n2716),
    .B1(net213),
    .C1(n3405),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2715));
 sky130_fd_sc_hd__o21a_1 U3100 (.A1(net213),
    .A2(n2717),
    .B1(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2714));
 sky130_fd_sc_hd__a32o_1 U3101 (.A1(net219),
    .A2(n3428),
    .A3(n2712),
    .B1(net219),
    .B2(\inst_to_wrap_u_usb_cdc_out_data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2713));
 sky130_fd_sc_hd__or3_1 U3102 (.A(n2714),
    .B(n2713),
    .C(n3379),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3407));
 sky130_fd_sc_hd__or4_1 U3103 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q),
    .B(n2715),
    .C(n3410),
    .D(n3407),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3427));
 sky130_fd_sc_hd__or2_1 U3104 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3425));
 sky130_fd_sc_hd__a22o_1 U3105 (.A1(net212),
    .A2(net219),
    .B1(n2717),
    .B2(n2716),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2718));
 sky130_fd_sc_hd__a31o_1 U3106 (.A1(net210),
    .A2(n3378),
    .A3(n3425),
    .B1(n2718),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2719));
 sky130_fd_sc_hd__a211o_1 U3107 (.A1(n3345),
    .A2(n3406),
    .B1(n3427),
    .C1(n2719),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2720));
 sky130_fd_sc_hd__or2_1 U3108 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .B(n3361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2941));
 sky130_fd_sc_hd__nor2_2 U3109 (.A(n2941),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3426));
 sky130_fd_sc_hd__o21a_1 U3110 (.A1(n3409),
    .A2(n2720),
    .B1(n3426),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2727));
 sky130_fd_sc_hd__nand2_1 U3111 (.A(n3417),
    .B(n3388),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3386));
 sky130_fd_sc_hd__inv_2 U3112 (.A(n2959),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3356));
 sky130_fd_sc_hd__o21a_1 U3113 (.A1(n2722),
    .A2(n3356),
    .B1(n2721),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3414));
 sky130_fd_sc_hd__a31o_1 U3114 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ),
    .A2(n3428),
    .A3(n2724),
    .B1(n2723),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2725));
 sky130_fd_sc_hd__a31o_1 U3115 (.A1(n3394),
    .A2(n3446),
    .A3(n2725),
    .B1(n2886),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2726));
 sky130_fd_sc_hd__o211ai_1 U3116 (.A1(n3386),
    .A2(n2962),
    .B1(n3414),
    .C1(n2726),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3430));
 sky130_fd_sc_hd__a211o_1 U3117 (.A1(n3416),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .B1(n2727),
    .C1(n3430),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2728));
 sky130_fd_sc_hd__o32a_1 U3118 (.A1(n3435),
    .A2(n3415),
    .A3(n2728),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ),
    .B2(n3438),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2228));
 sky130_fd_sc_hd__or3_1 U3119 (.A(n3010),
    .B(n3440),
    .C(n3442),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2729));
 sky130_fd_sc_hd__a211o_2 U3120 (.A1(n2885),
    .A2(net214),
    .B1(n3004),
    .C1(n2729),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3451));
 sky130_fd_sc_hd__inv_2 U3121 (.A(n2729),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2731));
 sky130_fd_sc_hd__inv_2 U3122 (.A(n3004),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3369));
 sky130_fd_sc_hd__a32o_2 U3123 (.A1(n2731),
    .A2(n2885),
    .A3(n2730),
    .B1(n2731),
    .B2(n3369),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3452));
 sky130_fd_sc_hd__o22a_1 U3124 (.A1(net218),
    .A2(n3451),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[3] ),
    .B2(n3452),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2227));
 sky130_fd_sc_hd__inv_1 U3125 (.A(n3468),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2735));
 sky130_fd_sc_hd__a22o_1 U3126 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ),
    .A2(n3469),
    .B1(n2732),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2733));
 sky130_fd_sc_hd__a21o_1 U3127 (.A1(n2735),
    .A2(n2734),
    .B1(n2733),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2737));
 sky130_fd_sc_hd__a32o_1 U3128 (.A1(n2739),
    .A2(n2738),
    .A3(n2737),
    .B1(n2736),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2226));
 sky130_fd_sc_hd__or4_2 U3129 (.A(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[3] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ),
    .D(n3079),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2868));
 sky130_fd_sc_hd__o211a_1 U3130 (.A1(n3068),
    .A2(n2868),
    .B1(n3087),
    .C1(n2740),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3076));
 sky130_fd_sc_hd__a221o_1 U3131 (.A1(n2743),
    .A2(n2742),
    .B1(n2743),
    .B2(n2741),
    .C1(n3068),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3069));
 sky130_fd_sc_hd__a32o_1 U3132 (.A1(n3076),
    .A2(n2745),
    .A3(n3069),
    .B1(n3076),
    .B2(n2744),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2747));
 sky130_fd_sc_hd__o211a_1 U3133 (.A1(n3068),
    .A2(n2748),
    .B1(n2747),
    .C1(n2746),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2749));
 sky130_fd_sc_hd__a2bb2o_1 U3134 (.A1_N(n2749),
    .A2_N(n3074),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ),
    .B2(n3029),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2225));
 sky130_fd_sc_hd__nor2_1 U3135 (.A(n3070),
    .B(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2758));
 sky130_fd_sc_hd__or2_2 U3136 (.A(n2774),
    .B(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2870));
 sky130_fd_sc_hd__a221o_1 U3137 (.A1(n2821),
    .A2(n2752),
    .B1(n2821),
    .B2(n2754),
    .C1(n2870),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2750));
 sky130_fd_sc_hd__a32o_1 U3138 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[2] ),
    .A2(n2751),
    .A3(n2753),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[3] ),
    .B2(n2750),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2224));
 sky130_fd_sc_hd__a21o_1 U3139 (.A1(n2821),
    .A2(n2752),
    .B1(n2870),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2755));
 sky130_fd_sc_hd__a22o_1 U3140 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[2] ),
    .A2(n2755),
    .B1(n2754),
    .B2(n2753),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2223));
 sky130_fd_sc_hd__a21o_1 U3141 (.A1(n2759),
    .A2(n2821),
    .B1(n2870),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2756));
 sky130_fd_sc_hd__a32o_1 U3142 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[0] ),
    .A2(n2757),
    .A3(n2758),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[1] ),
    .B2(n2756),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2222));
 sky130_fd_sc_hd__a22o_1 U3143 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[0] ),
    .A2(n2870),
    .B1(n2759),
    .B2(n2758),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2221));
 sky130_fd_sc_hd__or4_2 U3144 (.A(n2884),
    .B(n2761),
    .C(n2760),
    .D(n3344),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2787));
 sky130_fd_sc_hd__a32o_1 U3145 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[1] ),
    .A2(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_endp_q),
    .A3(n2786),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[1] ),
    .B2(n2787),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2768));
 sky130_fd_sc_hd__nor2_1 U3146 (.A(n3094),
    .B(n3086),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2762));
 sky130_fd_sc_hd__mux2_1 U3147 (.A0(n2768),
    .A1(n2763),
    .S(n2762),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2766));
 sky130_fd_sc_hd__nor2_1 U3148 (.A(n3074),
    .B(n3087),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2784));
 sky130_fd_sc_hd__o221a_1 U3149 (.A1(n2767),
    .A2(n2766),
    .B1(n2765),
    .B2(n2764),
    .C1(n2784),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2770));
 sky130_fd_sc_hd__o21a_1 U3150 (.A1(n3089),
    .A2(n3087),
    .B1(n2768),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2769));
 sky130_fd_sc_hd__a211o_1 U3151 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[1] ),
    .A2(n3029),
    .B1(n2770),
    .C1(n2769),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2220));
 sky130_fd_sc_hd__inv_1 U3152 (.A(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2783));
 sky130_fd_sc_hd__or2_1 U3153 (.A(n2990),
    .B(n3086),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2777));
 sky130_fd_sc_hd__inv_1 U3154 (.A(n2777),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2782));
 sky130_fd_sc_hd__nand2_1 U3155 (.A(n3057),
    .B(n2818),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3084));
 sky130_fd_sc_hd__o21ba_1 U3156 (.A1(n3079),
    .A2(n2771),
    .B1_N(n3064),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2776));
 sky130_fd_sc_hd__a21oi_1 U3157 (.A1(n3056),
    .A2(n2772),
    .B1(n3079),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2775));
 sky130_fd_sc_hd__a221o_1 U3158 (.A1(n2779),
    .A2(n2778),
    .B1(n2779),
    .B2(n2777),
    .C1(n3033),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2780));
 sky130_fd_sc_hd__a211o_1 U3159 (.A1(n3056),
    .A2(n3084),
    .B1(n3052),
    .C1(n2780),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2781));
 sky130_fd_sc_hd__a32o_1 U3160 (.A1(n2784),
    .A2(n2783),
    .A3(n2782),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[0] ),
    .B2(n2781),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2219));
 sky130_fd_sc_hd__nor2_1 U3161 (.A(n3089),
    .B(n3081),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2811));
 sky130_fd_sc_hd__inv_2 U3162 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_endp_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2785));
 sky130_fd_sc_hd__o221ai_2 U3163 (.A1(n2787),
    .A2(n2786),
    .B1(n2787),
    .B2(n2785),
    .C1(\inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2810));
 sky130_fd_sc_hd__inv_1 U3164 (.A(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2789));
 sky130_fd_sc_hd__o221a_1 U3165 (.A1(\inst_to_wrap_u_usb_cdc_addr[6] ),
    .A2(n2789),
    .B1(n2788),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[6] ),
    .C1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2802));
 sky130_fd_sc_hd__a22oi_1 U3166 (.A1(n2791),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[5] ),
    .B1(n2792),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2790));
 sky130_fd_sc_hd__o221a_1 U3167 (.A1(n2792),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[4] ),
    .B1(n2791),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[5] ),
    .C1(n2790),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2801));
 sky130_fd_sc_hd__a22oi_1 U3168 (.A1(n2794),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[3] ),
    .B1(n2795),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2793));
 sky130_fd_sc_hd__o221a_1 U3169 (.A1(n2795),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[2] ),
    .B1(n2794),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[3] ),
    .C1(n2793),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2800));
 sky130_fd_sc_hd__a22oi_1 U3170 (.A1(n2797),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[1] ),
    .B1(n2798),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2796));
 sky130_fd_sc_hd__o221a_1 U3171 (.A1(n2798),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[0] ),
    .B1(n2797),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[1] ),
    .C1(n2796),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2799));
 sky130_fd_sc_hd__and4_1 U3172 (.A(n2802),
    .B(n2801),
    .C(n2800),
    .D(n2799),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3063));
 sky130_fd_sc_hd__and3_1 U3173 (.A(n3063),
    .B(n3049),
    .C(n3065),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2804));
 sky130_fd_sc_hd__and3_1 U3174 (.A(n2804),
    .B(n3068),
    .C(n2803),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3082));
 sky130_fd_sc_hd__nand2_1 U3175 (.A(n2806),
    .B(n3082),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2808));
 sky130_fd_sc_hd__or2_1 U3176 (.A(n3074),
    .B(n3081),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2813));
 sky130_fd_sc_hd__a31o_1 U3177 (.A1(n2806),
    .A2(n3082),
    .A3(n2805),
    .B1(n2813),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2807));
 sky130_fd_sc_hd__a21o_1 U3178 (.A1(n2808),
    .A2(n2810),
    .B1(n2807),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2809));
 sky130_fd_sc_hd__o21ai_1 U3179 (.A1(n2811),
    .A2(n2810),
    .B1(n2809),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2812));
 sky130_fd_sc_hd__a21o_1 U3180 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[1] ),
    .A2(n3029),
    .B1(n2812),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2218));
 sky130_fd_sc_hd__inv_2 U3181 (.A(n2813),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3042));
 sky130_fd_sc_hd__and3_1 U3182 (.A(n2814),
    .B(n3042),
    .C(n3082),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2815));
 sky130_fd_sc_hd__mux2_1 U3183 (.A0(\inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[0] ),
    .A1(n2816),
    .S(n2815),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2817));
 sky130_fd_sc_hd__a31o_1 U3184 (.A1(n3057),
    .A2(n2818),
    .A3(n3036),
    .B1(n2817),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2217));
 sky130_fd_sc_hd__a21oi_4 U3185 (.A1(n3037),
    .A2(n2819),
    .B1(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2865));
 sky130_fd_sc_hd__inv_2 U3186 (.A(n2863),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2857));
 sky130_fd_sc_hd__inv_1 U3187 (.A(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2822));
 sky130_fd_sc_hd__and3_1 U3188 (.A(n2820),
    .B(n3079),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3034));
 sky130_fd_sc_hd__o21a_4 U3189 (.A1(n2821),
    .A2(n3034),
    .B1(n3045),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2859));
 sky130_fd_sc_hd__o221a_1 U3190 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[7] ),
    .A2(n2857),
    .B1(n2822),
    .B2(n2863),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2823));
 sky130_fd_sc_hd__a211o_1 U3191 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[15] ),
    .A2(n2866),
    .B1(n2865),
    .C1(n2823),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2216));
 sky130_fd_sc_hd__a22o_1 U3192 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[14] ),
    .A2(net184),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[6] ),
    .B2(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2824));
 sky130_fd_sc_hd__or2_1 U3193 (.A(n2865),
    .B(n2824),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2215));
 sky130_fd_sc_hd__a22o_1 U3194 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[13] ),
    .A2(net184),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[5] ),
    .B2(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2825));
 sky130_fd_sc_hd__or2_1 U3195 (.A(n2865),
    .B(n2825),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2214));
 sky130_fd_sc_hd__a22o_1 U3196 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[12] ),
    .A2(net184),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[4] ),
    .B2(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2826));
 sky130_fd_sc_hd__or2_1 U3197 (.A(n2865),
    .B(n2826),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2213));
 sky130_fd_sc_hd__a22o_1 U3198 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[11] ),
    .A2(net184),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[3] ),
    .B2(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2827));
 sky130_fd_sc_hd__or2_1 U3199 (.A(n2865),
    .B(n2827),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2212));
 sky130_fd_sc_hd__a22o_1 U3200 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[10] ),
    .A2(net184),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[2] ),
    .B2(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2828));
 sky130_fd_sc_hd__or2_1 U3201 (.A(n2865),
    .B(n2828),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2211));
 sky130_fd_sc_hd__o221a_1 U3202 (.A1(n2831),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[1] ),
    .B1(n2830),
    .B2(n2829),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2832));
 sky130_fd_sc_hd__a211o_1 U3203 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[9] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2832),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2210));
 sky130_fd_sc_hd__inv_1 U3204 (.A(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2834));
 sky130_fd_sc_hd__o221a_1 U3205 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[0] ),
    .A2(n2835),
    .B1(n2834),
    .B2(n2833),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2836));
 sky130_fd_sc_hd__a211o_1 U3206 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[8] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2836),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2209));
 sky130_fd_sc_hd__o221a_1 U3207 (.A1(n2838),
    .A2(n2841),
    .B1(n2837),
    .B2(n2840),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2839));
 sky130_fd_sc_hd__a211o_1 U3208 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[7] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2839),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2208));
 sky130_fd_sc_hd__inv_2 U3209 (.A(n2846),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2844));
 sky130_fd_sc_hd__o221a_1 U3210 (.A1(n2841),
    .A2(n2846),
    .B1(n2840),
    .B2(n2844),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2842));
 sky130_fd_sc_hd__a211o_1 U3211 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[6] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2842),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2207));
 sky130_fd_sc_hd__o221a_1 U3212 (.A1(n2846),
    .A2(n2845),
    .B1(n2844),
    .B2(n2843),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2847));
 sky130_fd_sc_hd__a211o_1 U3213 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[5] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2847),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2206));
 sky130_fd_sc_hd__a22o_1 U3214 (.A1(n2848),
    .A2(n2859),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[4] ),
    .B2(net184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2849));
 sky130_fd_sc_hd__or2_1 U3215 (.A(n2865),
    .B(n2849),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2205));
 sky130_fd_sc_hd__inv_1 U3216 (.A(n2850),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2852));
 sky130_fd_sc_hd__o221a_1 U3217 (.A1(n2853),
    .A2(n2852),
    .B1(n2851),
    .B2(n2850),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2854));
 sky130_fd_sc_hd__a211o_1 U3218 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[3] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2854),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2204));
 sky130_fd_sc_hd__o221a_1 U3219 (.A1(n2857),
    .A2(n2856),
    .B1(n2863),
    .B2(n2855),
    .C1(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2858));
 sky130_fd_sc_hd__a211o_1 U3220 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[2] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2858),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2203));
 sky130_fd_sc_hd__inv_2 U3221 (.A(n2859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2862));
 sky130_fd_sc_hd__nor2_1 U3222 (.A(n2860),
    .B(n2862),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2861));
 sky130_fd_sc_hd__a211o_1 U3223 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[1] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2202));
 sky130_fd_sc_hd__nor2_1 U3224 (.A(n2863),
    .B(n2862),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2864));
 sky130_fd_sc_hd__a211o_1 U3225 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[0] ),
    .A2(net184),
    .B1(n2865),
    .C1(n2864),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2201));
 sky130_fd_sc_hd__inv_2 U3226 (.A(n3034),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2867));
 sky130_fd_sc_hd__a21oi_4 U3227 (.A1(n2868),
    .A2(n2867),
    .B1(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2869));
 sky130_fd_sc_hd__a22o_1 U3228 (.A1(\inst_to_wrap_u_usb_cdc_out_data[7] ),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2200));
 sky130_fd_sc_hd__a22o_1 U3229 (.A1(net215),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[6] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2199));
 sky130_fd_sc_hd__a22o_1 U3230 (.A1(net216),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[5] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2198));
 sky130_fd_sc_hd__a22o_1 U3231 (.A1(net217),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[4] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2197));
 sky130_fd_sc_hd__a22o_1 U3232 (.A1(net218),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[3] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2196));
 sky130_fd_sc_hd__a22o_1 U3233 (.A1(net219),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2195));
 sky130_fd_sc_hd__a22o_1 U3234 (.A1(net210),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2194));
 sky130_fd_sc_hd__a22o_1 U3235 (.A1(net212),
    .A2(net185),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ),
    .B2(n2869),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2193));
 sky130_fd_sc_hd__inv_2 U3236 (.A(n2870),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3032));
 sky130_fd_sc_hd__nor2_2 U3239 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ),
    .B(n2923),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3007));
 sky130_fd_sc_hd__and2_1 U3240 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .B(n3007),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2963));
 sky130_fd_sc_hd__and3_1 U3241 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .B(n3433),
    .C(n2963),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2872));
 sky130_fd_sc_hd__a31o_1 U3242 (.A1(n3004),
    .A2(n2954),
    .A3(n3359),
    .B1(n2872),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2881));
 sky130_fd_sc_hd__inv_2 U3243 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3328));
 sky130_fd_sc_hd__or4_2 U3244 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .C(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .D(n3328),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3101));
 sky130_fd_sc_hd__clkinv_2 U3245 (.A(n3101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2981));
 sky130_fd_sc_hd__clkinv_2 U3246 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3330));
 sky130_fd_sc_hd__nor2_1 U3247 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .B(n3330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3109));
 sky130_fd_sc_hd__inv_2 U3248 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3326));
 sky130_fd_sc_hd__and3_2 U3249 (.A(n3109),
    .B(n3328),
    .C(n3326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2980));
 sky130_fd_sc_hd__a22o_1 U3250 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[71] ),
    .B1(n2980),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2879));
 sky130_fd_sc_hd__nor2_1 U3251 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2873));
 sky130_fd_sc_hd__inv_2 U3252 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3323));
 sky130_fd_sc_hd__and3_2 U3253 (.A(n2873),
    .B(n3330),
    .C(n3323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2983));
 sky130_fd_sc_hd__nor2_1 U3254 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ),
    .B(n3326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2874));
 sky130_fd_sc_hd__and2_2 U3255 (.A(n2874),
    .B(n3109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2982));
 sky130_fd_sc_hd__a22o_1 U3256 (.A1(n2983),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[7] ),
    .B1(n2982),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2878));
 sky130_fd_sc_hd__and3_2 U3257 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .C(n2874),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3103));
 sky130_fd_sc_hd__and3_2 U3258 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .B(n2873),
    .C(n3330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2985));
 sky130_fd_sc_hd__and3_2 U3259 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .B(n2874),
    .C(n3330),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2984));
 sky130_fd_sc_hd__a22o_1 U3260 (.A1(n2985),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[39] ),
    .B1(n2984),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2876));
 sky130_fd_sc_hd__and3_2 U3261 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .C(n2873),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2987));
 sky130_fd_sc_hd__and3_2 U3262 (.A(n2874),
    .B(n3330),
    .C(n3323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2986));
 sky130_fd_sc_hd__a22o_1 U3263 (.A1(n2987),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[55] ),
    .B1(n2986),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2875));
 sky130_fd_sc_hd__a211o_1 U3264 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[63] ),
    .B1(n2876),
    .C1(n2875),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2877));
 sky130_fd_sc_hd__o31a_1 U3265 (.A1(n2879),
    .A2(n2878),
    .A3(n2877),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2880));
 sky130_fd_sc_hd__nand2_1 U3266 (.A(n3007),
    .B(n3005),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2961));
 sky130_fd_sc_hd__clkinv_2 U3267 (.A(n2961),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3011));
 sky130_fd_sc_hd__and3_1 U3268 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .B(n3418),
    .C(n3011),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2946));
 sky130_fd_sc_hd__and2_1 U3269 (.A(n2946),
    .B(n3023),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2931));
 sky130_fd_sc_hd__a211o_1 U3270 (.A1(n3023),
    .A2(n2881),
    .B1(n2880),
    .C1(n2931),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2883));
 sky130_fd_sc_hd__and2_1 U3271 (.A(n2908),
    .B(n3080),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3028));
 sky130_fd_sc_hd__a22o_1 U3272 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ),
    .A2(net185),
    .B1(n3028),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2882));
 sky130_fd_sc_hd__a21o_1 U3273 (.A1(n3032),
    .A2(n2883),
    .B1(n2882),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2192));
 sky130_fd_sc_hd__inv_2 U3274 (.A(n2941),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3019));
 sky130_fd_sc_hd__a21oi_1 U3275 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .A2(n3361),
    .B1(n3019),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2911));
 sky130_fd_sc_hd__and4_1 U3276 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .B(n2885),
    .C(n2996),
    .D(n2884),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3021));
 sky130_fd_sc_hd__and3_1 U3277 (.A(n3372),
    .B(n3021),
    .C(n3010),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3026));
 sky130_fd_sc_hd__nor2_1 U3278 (.A(n2956),
    .B(n2886),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2942));
 sky130_fd_sc_hd__a22o_1 U3279 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[70] ),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[22] ),
    .B2(n2980),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2891));
 sky130_fd_sc_hd__a22o_1 U3280 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[6] ),
    .A2(n2983),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[30] ),
    .B2(n2982),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2890));
 sky130_fd_sc_hd__a22o_1 U3281 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[38] ),
    .A2(n2985),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[46] ),
    .B2(n2984),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2888));
 sky130_fd_sc_hd__a22o_1 U3282 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[54] ),
    .A2(n2987),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[14] ),
    .B2(n2986),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2887));
 sky130_fd_sc_hd__a211o_1 U3283 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[62] ),
    .B1(n2888),
    .C1(n2887),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2889));
 sky130_fd_sc_hd__o31a_1 U3284 (.A1(n2891),
    .A2(n2890),
    .A3(n2889),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2892));
 sky130_fd_sc_hd__a31o_1 U3285 (.A1(n3023),
    .A2(n2954),
    .A3(n2942),
    .B1(n2892),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2893));
 sky130_fd_sc_hd__a211o_1 U3286 (.A1(n2911),
    .A2(n3026),
    .B1(n2931),
    .C1(n2893),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2894));
 sky130_fd_sc_hd__a22o_1 U3287 (.A1(net185),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[6] ),
    .B1(n3032),
    .B2(n2894),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2895));
 sky130_fd_sc_hd__a31o_1 U3288 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[6] ),
    .A2(n2908),
    .A3(n3080),
    .B1(n2895),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2191));
 sky130_fd_sc_hd__a22o_1 U3289 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[69] ),
    .B1(n2980),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2900));
 sky130_fd_sc_hd__a22o_1 U3290 (.A1(n2983),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[5] ),
    .B1(n2982),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2899));
 sky130_fd_sc_hd__a22o_1 U3291 (.A1(n2985),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[37] ),
    .B1(n2984),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2897));
 sky130_fd_sc_hd__a22o_1 U3292 (.A1(n2987),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[53] ),
    .B1(n2986),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2896));
 sky130_fd_sc_hd__a211o_1 U3293 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[61] ),
    .B1(n2897),
    .C1(n2896),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2898));
 sky130_fd_sc_hd__o31a_1 U3294 (.A1(n2900),
    .A2(n2899),
    .A3(n2898),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2905));
 sky130_fd_sc_hd__nor2_1 U3295 (.A(n2956),
    .B(n3356),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2902));
 sky130_fd_sc_hd__and3_1 U3296 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .B(n2998),
    .C(n3019),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2910));
 sky130_fd_sc_hd__a22o_1 U3297 (.A1(n3418),
    .A2(n2998),
    .B1(n3426),
    .B2(n3011),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2901));
 sky130_fd_sc_hd__o32a_1 U3298 (.A1(n2902),
    .A2(n2910),
    .A3(n3368),
    .B1(n2901),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2903));
 sky130_fd_sc_hd__a22o_1 U3299 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .A2(n3026),
    .B1(n3023),
    .B2(n2903),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2904));
 sky130_fd_sc_hd__or3_1 U3300 (.A(n2931),
    .B(n2905),
    .C(n2904),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2906));
 sky130_fd_sc_hd__a22o_1 U3301 (.A1(net185),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[5] ),
    .B1(n3032),
    .B2(n2906),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2907));
 sky130_fd_sc_hd__a31o_1 U3302 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[5] ),
    .A2(n2908),
    .A3(n3080),
    .B1(n2907),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2190));
 sky130_fd_sc_hd__a32o_1 U3303 (.A1(n3023),
    .A2(n2910),
    .A3(n3368),
    .B1(n3023),
    .B2(n2909),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2921));
 sky130_fd_sc_hd__inv_2 U3304 (.A(n2911),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3362));
 sky130_fd_sc_hd__a22o_1 U3305 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[68] ),
    .B1(n2980),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2916));
 sky130_fd_sc_hd__a22o_1 U3306 (.A1(n2983),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[4] ),
    .B1(n2982),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2915));
 sky130_fd_sc_hd__a22o_1 U3307 (.A1(n2985),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[36] ),
    .B1(n2984),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2913));
 sky130_fd_sc_hd__a22o_1 U3308 (.A1(n2987),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[52] ),
    .B1(n2986),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2912));
 sky130_fd_sc_hd__a211o_1 U3309 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[60] ),
    .B1(n2913),
    .C1(n2912),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2914));
 sky130_fd_sc_hd__o31a_1 U3310 (.A1(n2916),
    .A2(n2915),
    .A3(n2914),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2917));
 sky130_fd_sc_hd__a211o_1 U3311 (.A1(n3026),
    .A2(n3362),
    .B1(n2917),
    .C1(n2931),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2918));
 sky130_fd_sc_hd__a31o_1 U3312 (.A1(n2959),
    .A2(n3021),
    .A3(n3005),
    .B1(n2918),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2920));
 sky130_fd_sc_hd__a22o_1 U3313 (.A1(net185),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[4] ),
    .B1(n3028),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2919));
 sky130_fd_sc_hd__a221o_1 U3314 (.A1(n3032),
    .A2(n2921),
    .B1(n3032),
    .B2(n2920),
    .C1(n2919),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2189));
 sky130_fd_sc_hd__a22o_1 U3315 (.A1(n3007),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .B1(n3372),
    .B2(n3359),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2958));
 sky130_fd_sc_hd__and3_1 U3316 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .B(n3434),
    .C(n3011),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2922));
 sky130_fd_sc_hd__a31o_1 U3317 (.A1(n2959),
    .A2(n2954),
    .A3(n2923),
    .B1(n2922),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2924));
 sky130_fd_sc_hd__a32o_1 U3318 (.A1(n3023),
    .A2(n3426),
    .A3(n2958),
    .B1(n3023),
    .B2(n2924),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2935));
 sky130_fd_sc_hd__a22o_1 U3319 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[67] ),
    .B1(n2980),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2929));
 sky130_fd_sc_hd__a22o_1 U3320 (.A1(n2983),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[3] ),
    .B1(n2982),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2928));
 sky130_fd_sc_hd__a22o_1 U3321 (.A1(n2985),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[35] ),
    .B1(n2984),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2926));
 sky130_fd_sc_hd__a22o_1 U3322 (.A1(n2987),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[51] ),
    .B1(n2986),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2925));
 sky130_fd_sc_hd__a211o_1 U3323 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[59] ),
    .B1(n2926),
    .C1(n2925),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2927));
 sky130_fd_sc_hd__o31a_1 U3324 (.A1(n2929),
    .A2(n2928),
    .A3(n2927),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2930));
 sky130_fd_sc_hd__a211o_1 U3325 (.A1(n3019),
    .A2(n3026),
    .B1(n2931),
    .C1(n2930),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2932));
 sky130_fd_sc_hd__a31o_1 U3326 (.A1(n3004),
    .A2(n2954),
    .A3(n3021),
    .B1(n2932),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2934));
 sky130_fd_sc_hd__a22o_1 U3327 (.A1(net185),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[3] ),
    .B1(n3028),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2933));
 sky130_fd_sc_hd__a221o_1 U3328 (.A1(n3032),
    .A2(n2935),
    .B1(n3032),
    .B2(n2934),
    .C1(n2933),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2188));
 sky130_fd_sc_hd__a22o_1 U3329 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[66] ),
    .B1(n2980),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2940));
 sky130_fd_sc_hd__a22o_1 U3330 (.A1(n2983),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[2] ),
    .B1(n2982),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2939));
 sky130_fd_sc_hd__a22o_1 U3331 (.A1(n2985),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[34] ),
    .B1(n2984),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2937));
 sky130_fd_sc_hd__a22o_1 U3332 (.A1(n2987),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[50] ),
    .B1(n2986),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2936));
 sky130_fd_sc_hd__a211o_1 U3333 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[58] ),
    .B1(n2937),
    .C1(n2936),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2938));
 sky130_fd_sc_hd__o31a_1 U3334 (.A1(n2940),
    .A2(n2939),
    .A3(n2938),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2951));
 sky130_fd_sc_hd__nor2_1 U3335 (.A(n3010),
    .B(n2941),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3003));
 sky130_fd_sc_hd__nor2_1 U3336 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ),
    .B(n3005),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3008));
 sky130_fd_sc_hd__a22o_1 U3337 (.A1(n2959),
    .A2(n2998),
    .B1(n2942),
    .B2(n3005),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2943));
 sky130_fd_sc_hd__a31o_1 U3338 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .A2(n3008),
    .A3(n3440),
    .B1(n2943),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2948));
 sky130_fd_sc_hd__or2_1 U3339 (.A(n3027),
    .B(n3416),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2944));
 sky130_fd_sc_hd__a22o_1 U3340 (.A1(n2998),
    .A2(n2944),
    .B1(n3433),
    .B2(n3007),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2945));
 sky130_fd_sc_hd__a31o_1 U3341 (.A1(n3011),
    .A2(n3010),
    .A3(n3363),
    .B1(n2945),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2947));
 sky130_fd_sc_hd__a31o_1 U3342 (.A1(n3007),
    .A2(n3003),
    .A3(n3368),
    .B1(n2946),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3013));
 sky130_fd_sc_hd__a221o_1 U3343 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .A2(n2948),
    .B1(n3368),
    .B2(n2947),
    .C1(n3013),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2949));
 sky130_fd_sc_hd__a32o_1 U3344 (.A1(n3023),
    .A2(n3011),
    .A3(n3003),
    .B1(n3023),
    .B2(n2949),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2950));
 sky130_fd_sc_hd__a211o_1 U3345 (.A1(n3026),
    .A2(n3019),
    .B1(n2951),
    .C1(n2950),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2953));
 sky130_fd_sc_hd__a22o_1 U3346 (.A1(net185),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .B1(n3028),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2952));
 sky130_fd_sc_hd__a21o_1 U3347 (.A1(n3032),
    .A2(n2953),
    .B1(n2952),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2187));
 sky130_fd_sc_hd__o211a_1 U3348 (.A1(n3002),
    .A2(n3418),
    .B1(n2954),
    .C1(n3021),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2979));
 sky130_fd_sc_hd__nor2_1 U3349 (.A(n2956),
    .B(n2955),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2957));
 sky130_fd_sc_hd__a22o_1 U3350 (.A1(n2959),
    .A2(n2958),
    .B1(n2957),
    .B2(n3434),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2976));
 sky130_fd_sc_hd__and3_1 U3351 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .B(n3019),
    .C(n3007),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2968));
 sky130_fd_sc_hd__a21o_1 U3352 (.A1(n3005),
    .A2(n3012),
    .B1(n2963),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2999));
 sky130_fd_sc_hd__a22o_1 U3353 (.A1(n3004),
    .A2(n3011),
    .B1(n3426),
    .B2(n2999),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2960));
 sky130_fd_sc_hd__a31o_1 U3354 (.A1(n3416),
    .A2(n3359),
    .A3(n3005),
    .B1(n2960),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2967));
 sky130_fd_sc_hd__nor2_1 U3355 (.A(n2962),
    .B(n2961),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2965));
 sky130_fd_sc_hd__a22o_1 U3356 (.A1(n3004),
    .A2(n2999),
    .B1(n3434),
    .B2(n2963),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2964));
 sky130_fd_sc_hd__a211o_1 U3357 (.A1(n3433),
    .A2(n3012),
    .B1(n2965),
    .C1(n2964),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2966));
 sky130_fd_sc_hd__o32a_1 U3358 (.A1(n2968),
    .A2(n2967),
    .A3(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .B1(n2966),
    .B2(n3368),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2975));
 sky130_fd_sc_hd__a22o_1 U3359 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[65] ),
    .B1(n2980),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2973));
 sky130_fd_sc_hd__a22o_1 U3360 (.A1(n2983),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[1] ),
    .B1(n2982),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2972));
 sky130_fd_sc_hd__a22o_1 U3361 (.A1(n2985),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[33] ),
    .B1(n2984),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2970));
 sky130_fd_sc_hd__a22o_1 U3362 (.A1(n2987),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[49] ),
    .B1(n2986),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2969));
 sky130_fd_sc_hd__a211o_1 U3363 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[57] ),
    .B1(n2970),
    .C1(n2969),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2971));
 sky130_fd_sc_hd__o31a_1 U3364 (.A1(n2973),
    .A2(n2972),
    .A3(n2971),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2974));
 sky130_fd_sc_hd__a221o_1 U3365 (.A1(n3023),
    .A2(n2976),
    .B1(n3023),
    .B2(n2975),
    .C1(n2974),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2978));
 sky130_fd_sc_hd__a22o_1 U3366 (.A1(net185),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .B1(n3028),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2977));
 sky130_fd_sc_hd__a221o_1 U3367 (.A1(n3032),
    .A2(n2979),
    .B1(n3032),
    .B2(n2978),
    .C1(n2977),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2186));
 sky130_fd_sc_hd__a22o_1 U3368 (.A1(n2981),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[64] ),
    .B1(n2980),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2993));
 sky130_fd_sc_hd__a22o_1 U3369 (.A1(n2983),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[0] ),
    .B1(n2982),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2992));
 sky130_fd_sc_hd__a22o_1 U3370 (.A1(n2985),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[32] ),
    .B1(n2984),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2989));
 sky130_fd_sc_hd__a22o_1 U3371 (.A1(n2987),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[48] ),
    .B1(n2986),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2988));
 sky130_fd_sc_hd__a211o_1 U3372 (.A1(n3103),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[56] ),
    .B1(n2989),
    .C1(n2988),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2991));
 sky130_fd_sc_hd__o31a_1 U3373 (.A1(n2993),
    .A2(n2992),
    .A3(n2991),
    .B1(n2990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2994));
 sky130_fd_sc_hd__a31o_1 U3374 (.A1(n2997),
    .A2(n2996),
    .A3(n2995),
    .B1(n2994),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3025));
 sky130_fd_sc_hd__and2_1 U3375 (.A(n3418),
    .B(n2998),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3001));
 sky130_fd_sc_hd__o221a_1 U3376 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .A2(n3012),
    .B1(n3010),
    .B2(n2999),
    .C1(n3019),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3000));
 sky130_fd_sc_hd__a211o_1 U3377 (.A1(n3011),
    .A2(n3002),
    .B1(n3001),
    .C1(n3000),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3018));
 sky130_fd_sc_hd__a31o_1 U3378 (.A1(n3440),
    .A2(n3361),
    .A3(n3011),
    .B1(n3003),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3006));
 sky130_fd_sc_hd__o221a_1 U3379 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .A2(n3006),
    .B1(n3005),
    .B2(n3004),
    .C1(n3359),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3017));
 sky130_fd_sc_hd__a32o_1 U3380 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .A2(n3368),
    .A3(n3008),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .B2(n3007),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3009));
 sky130_fd_sc_hd__or3_1 U3381 (.A(n3011),
    .B(n3010),
    .C(n3009),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3015));
 sky130_fd_sc_hd__a21o_1 U3382 (.A1(n3368),
    .A2(n3012),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3014));
 sky130_fd_sc_hd__a31o_1 U3383 (.A1(n3361),
    .A2(n3015),
    .A3(n3014),
    .B1(n3013),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3016));
 sky130_fd_sc_hd__a221o_1 U3384 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .A2(n3018),
    .B1(n3368),
    .B2(n3017),
    .C1(n3016),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3022));
 sky130_fd_sc_hd__a22o_1 U3385 (.A1(n3019),
    .A2(n3372),
    .B1(n3426),
    .B2(n3368),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3020));
 sky130_fd_sc_hd__a22o_1 U3386 (.A1(n3023),
    .A2(n3022),
    .B1(n3021),
    .B2(n3020),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3024));
 sky130_fd_sc_hd__a211o_1 U3387 (.A1(n3027),
    .A2(n3026),
    .B1(n3025),
    .C1(n3024),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3031));
 sky130_fd_sc_hd__a22o_1 U3388 (.A1(net185),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ),
    .B1(n3028),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3030));
 sky130_fd_sc_hd__a21o_1 U3389 (.A1(n3032),
    .A2(n3031),
    .B1(n3030),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2185));
 sky130_fd_sc_hd__or2_4 U3390 (.A(n3034),
    .B(n3033),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3035));
 sky130_fd_sc_hd__a22o_1 U3391 (.A1(\inst_to_wrap_u_usb_cdc_endp[3] ),
    .A2(n3035),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .B2(n3036),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2184));
 sky130_fd_sc_hd__a22o_1 U3392 (.A1(\inst_to_wrap_u_usb_cdc_endp[2] ),
    .A2(n3035),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .B2(n3036),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2183));
 sky130_fd_sc_hd__a22o_1 U3393 (.A1(\inst_to_wrap_u_usb_cdc_endp[1] ),
    .A2(n3035),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ),
    .B2(n3036),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2182));
 sky130_fd_sc_hd__a22o_1 U3394 (.A1(\inst_to_wrap_u_usb_cdc_endp[0] ),
    .A2(n3035),
    .B1(net214),
    .B2(n3036),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2181));
 sky130_fd_sc_hd__a22o_1 U3395 (.A1(net215),
    .A2(n3036),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[6] ),
    .B2(n3035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2180));
 sky130_fd_sc_hd__a22o_1 U3396 (.A1(net216),
    .A2(n3036),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[5] ),
    .B2(n3035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2179));
 sky130_fd_sc_hd__a22o_1 U3397 (.A1(net217),
    .A2(n3036),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[4] ),
    .B2(n3035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2178));
 sky130_fd_sc_hd__a22o_1 U3398 (.A1(net218),
    .A2(n3036),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[3] ),
    .B2(n3035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2177));
 sky130_fd_sc_hd__a22o_1 U3399 (.A1(\inst_to_wrap_u_usb_cdc_out_data[2] ),
    .A2(n3036),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[2] ),
    .B2(n3035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2176));
 sky130_fd_sc_hd__a22o_1 U3400 (.A1(net210),
    .A2(n3036),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[1] ),
    .B2(n3035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2175));
 sky130_fd_sc_hd__a22o_1 U3401 (.A1(net212),
    .A2(n3036),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[0] ),
    .B2(n3035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2174));
 sky130_fd_sc_hd__a21oi_1 U3402 (.A1(n3037),
    .A2(n3087),
    .B1(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3041));
 sky130_fd_sc_hd__a22o_1 U3403 (.A1(n3038),
    .A2(n3041),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ),
    .B2(n3042),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3039));
 sky130_fd_sc_hd__a21o_1 U3404 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[2] ),
    .A2(n3043),
    .B1(n3039),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2172));
 sky130_fd_sc_hd__a22o_1 U3405 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[1] ),
    .A2(n3043),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ),
    .B2(n3042),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3040));
 sky130_fd_sc_hd__or2_1 U3406 (.A(n3041),
    .B(n3040),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2171));
 sky130_fd_sc_hd__a22o_1 U3407 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[0] ),
    .A2(n3043),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ),
    .B2(n3042),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3044));
 sky130_fd_sc_hd__a31o_1 U3408 (.A1(n3047),
    .A2(n3046),
    .A3(n3045),
    .B1(n3044),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2170));
 sky130_fd_sc_hd__nor2_1 U3409 (.A(n3049),
    .B(n3048),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3062));
 sky130_fd_sc_hd__a31oi_1 U3410 (.A1(n3062),
    .A2(n3079),
    .A3(n3050),
    .B1(n3064),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3053));
 sky130_fd_sc_hd__o21ai_1 U3411 (.A1(n3053),
    .A2(n3052),
    .B1(n3051),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3054));
 sky130_fd_sc_hd__a31o_1 U3412 (.A1(n3069),
    .A2(n3087),
    .A3(n3054),
    .B1(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3055));
 sky130_fd_sc_hd__o21ai_1 U3413 (.A1(n3080),
    .A2(n3056),
    .B1(n3055),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2169));
 sky130_fd_sc_hd__a31o_1 U3414 (.A1(n3060),
    .A2(n3059),
    .A3(n3058),
    .B1(n3057),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3061));
 sky130_fd_sc_hd__and3_1 U3415 (.A(n3063),
    .B(n3062),
    .C(n3061),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3066));
 sky130_fd_sc_hd__a31o_1 U3416 (.A1(n3066),
    .A2(n3079),
    .A3(n3065),
    .B1(n3064),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3067));
 sky130_fd_sc_hd__o22a_1 U3417 (.A1(n3079),
    .A2(n3069),
    .B1(n3068),
    .B2(n3067),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3077));
 sky130_fd_sc_hd__o22a_1 U3418 (.A1(n3073),
    .A2(n3072),
    .B1(n3071),
    .B2(n3070),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3075));
 sky130_fd_sc_hd__a31o_1 U3419 (.A1(n3077),
    .A2(n3076),
    .A3(n3075),
    .B1(n3074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3078));
 sky130_fd_sc_hd__o21ai_1 U3420 (.A1(n3080),
    .A2(n3079),
    .B1(n3078),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2168));
 sky130_fd_sc_hd__o22a_1 U3421 (.A1(n3087),
    .A2(n3086),
    .B1(n3085),
    .B2(n3084),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3088));
 sky130_fd_sc_hd__nor2_1 U3422 (.A(n3089),
    .B(n3088),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3090));
 sky130_fd_sc_hd__a211o_1 U3423 (.A1(inst_to_wrap_u_usb_cdc_u_sie_out_eop_q),
    .A2(n3093),
    .B1(n3092),
    .C1(n3090),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2167));
 sky130_fd_sc_hd__or2_2 U3424 (.A(n3091),
    .B(n3094),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3569));
 sky130_fd_sc_hd__inv_2 U3425 (.A(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_state_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3097));
 sky130_fd_sc_hd__a32o_1 U3426 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_state_q),
    .A2(n3477),
    .A3(n3569),
    .B1(n3097),
    .B2(n3841),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2166));
 sky130_fd_sc_hd__a21o_1 U3427 (.A1(inst_to_wrap_u_usb_cdc_in_data_ack),
    .A2(n3093),
    .B1(n3092),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2165));
 sky130_fd_sc_hd__inv_2 U3428 (.A(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3106));
 sky130_fd_sc_hd__and2_1 U3429 (.A(n3106),
    .B(n3841),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3341));
 sky130_fd_sc_hd__or2_1 U3430 (.A(n3095),
    .B(n3094),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3099));
 sky130_fd_sc_hd__nor2_1 U3431 (.A(n3106),
    .B(n3099),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3112));
 sky130_fd_sc_hd__nor2_1 U3432 (.A(n3341),
    .B(n3112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3100));
 sky130_fd_sc_hd__and2_1 U3433 (.A(n3101),
    .B(n3112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3102));
 sky130_fd_sc_hd__a22o_1 U3434 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .A2(n3341),
    .B1(n3102),
    .B2(n3326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3096));
 sky130_fd_sc_hd__a21o_1 U3435 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .A2(n3100),
    .B1(n3096),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2164));
 sky130_fd_sc_hd__or2_1 U3436 (.A(n3097),
    .B(n3841),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3098));
 sky130_fd_sc_hd__or4_2 U3437 (.A(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q),
    .B(n3099),
    .C(n3344),
    .D(n3098),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3113));
 sky130_fd_sc_hd__inv_2 U3438 (.A(n3113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3114));
 sky130_fd_sc_hd__mux2_1 U3439 (.A0(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .S(n3114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2163));
 sky130_fd_sc_hd__a31o_1 U3440 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q),
    .A2(n3326),
    .A3(n3101),
    .B1(n3100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3110));
 sky130_fd_sc_hd__a31o_1 U3441 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q),
    .A2(n3330),
    .A3(n3101),
    .B1(n3110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3107));
 sky130_fd_sc_hd__a31o_1 U3442 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q),
    .A2(n3323),
    .A3(n3101),
    .B1(n3107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3104));
 sky130_fd_sc_hd__a22o_1 U3443 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ),
    .A2(n3104),
    .B1(n3103),
    .B2(n3102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3105));
 sky130_fd_sc_hd__a31o_1 U3444 (.A1(n3841),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ),
    .A3(n3106),
    .B1(n3105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2162));
 sky130_fd_sc_hd__a22o_1 U3445 (.A1(n3114),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ),
    .B1(n3113),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2161));
 sky130_fd_sc_hd__a22o_1 U3446 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .A2(n3107),
    .B1(n3341),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3108));
 sky130_fd_sc_hd__a31o_1 U3447 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .A2(n3112),
    .A3(n3109),
    .B1(n3108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2160));
 sky130_fd_sc_hd__a22o_1 U3448 (.A1(n3114),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .B1(n3113),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2159));
 sky130_fd_sc_hd__a22o_1 U3449 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ),
    .A2(n3110),
    .B1(n3341),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3111));
 sky130_fd_sc_hd__a31o_1 U3450 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .A2(n3112),
    .A3(n3330),
    .B1(n3111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2158));
 sky130_fd_sc_hd__a22o_1 U3451 (.A1(n3114),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ),
    .B1(n3113),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2157));
 sky130_fd_sc_hd__o21a_1 U3452 (.A1(n3325),
    .A2(n3121),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3115));
 sky130_fd_sc_hd__a31o_1 U3453 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .A2(n3123),
    .A3(n3331),
    .B1(n3115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2156));
 sky130_fd_sc_hd__a32o_1 U3454 (.A1(n3123),
    .A2(n3325),
    .A3(n3116),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .B2(n3121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2155));
 sky130_fd_sc_hd__a32o_1 U3455 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .A2(n3337),
    .A3(n3118),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .B2(n3117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2154));
 sky130_fd_sc_hd__and3_1 U3456 (.A(n3123),
    .B(n3333),
    .C(n3331),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3119));
 sky130_fd_sc_hd__and3_2 U3457 (.A(n3119),
    .B(n3337),
    .C(n3325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3306));
 sky130_fd_sc_hd__clkinv_2 U3458 (.A(n3306),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3305));
 sky130_fd_sc_hd__a22o_1 U3459 (.A1(n3306),
    .A2(net91),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2152));
 sky130_fd_sc_hd__and3_2 U3460 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .B(n3119),
    .C(n3337),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3308));
 sky130_fd_sc_hd__clkinv_2 U3461 (.A(n3308),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3307));
 sky130_fd_sc_hd__a22o_1 U3462 (.A1(n3308),
    .A2(net96),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2151));
 sky130_fd_sc_hd__and3_2 U3463 (.A(n3120),
    .B(n3337),
    .C(n3325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3310));
 sky130_fd_sc_hd__clkinv_2 U3464 (.A(n3310),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3309));
 sky130_fd_sc_hd__a22o_1 U3465 (.A1(n3310),
    .A2(net96),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2150));
 sky130_fd_sc_hd__and3_2 U3466 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .B(n3120),
    .C(n3337),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3312));
 sky130_fd_sc_hd__clkinv_2 U3467 (.A(n3312),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3311));
 sky130_fd_sc_hd__a22o_1 U3468 (.A1(n3312),
    .A2(net96),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2149));
 sky130_fd_sc_hd__and3_2 U3469 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .B(n3119),
    .C(n3325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3314));
 sky130_fd_sc_hd__clkinv_2 U3470 (.A(n3314),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3313));
 sky130_fd_sc_hd__a22o_1 U3471 (.A1(n3314),
    .A2(net96),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2148));
 sky130_fd_sc_hd__and3_2 U3472 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .C(n3119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3316));
 sky130_fd_sc_hd__clkinv_2 U3473 (.A(n3316),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3315));
 sky130_fd_sc_hd__a22o_1 U3474 (.A1(n3316),
    .A2(net96),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2147));
 sky130_fd_sc_hd__and3_2 U3475 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .B(n3120),
    .C(n3325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3318));
 sky130_fd_sc_hd__clkinv_2 U3476 (.A(n3318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3317));
 sky130_fd_sc_hd__a22o_1 U3477 (.A1(n3318),
    .A2(net96),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2146));
 sky130_fd_sc_hd__clkinv_2 U3478 (.A(n3320),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3319));
 sky130_fd_sc_hd__a22o_1 U3479 (.A1(n3320),
    .A2(net96),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2145));
 sky130_fd_sc_hd__mux2_1 U3480 (.A0(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[0] ),
    .A1(n3121),
    .S(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2144));
 sky130_fd_sc_hd__nand2_1 U3481 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[1] ),
    .B(n3121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3122));
 sky130_fd_sc_hd__nand2_1 U3482 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[0] ),
    .B(n3122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n2143));
 sky130_fd_sc_hd__nand2_1 U3483 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3124));
 sky130_fd_sc_hd__a221o_1 U3484 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_mask_q),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq[0] ),
    .B1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_mask_q),
    .B2(n3124),
    .C1(n3123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2142));
 sky130_fd_sc_hd__a21o_1 U3485 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_mask_q),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq[0] ),
    .B1(n3304),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2141));
 sky130_fd_sc_hd__a21o_1 U3486 (.A1(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A2(net209),
    .B1(n3300),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2140));
 sky130_fd_sc_hd__nand2_1 U3487 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .B(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3177));
 sky130_fd_sc_hd__o21a_1 U3488 (.A1(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .A2(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ),
    .B1(n3177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3152));
 sky130_fd_sc_hd__nand2_1 U3489 (.A(n3158),
    .B(n3152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3129));
 sky130_fd_sc_hd__nor2_1 U3490 (.A(n3190),
    .B(n3177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3125));
 sky130_fd_sc_hd__mux2_1 U3491 (.A0(\inst_to_wrap_tx_fifo_w_ptr_reg[3] ),
    .A1(n3193),
    .S(n3125),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3154));
 sky130_fd_sc_hd__a22oi_1 U3492 (.A1(n3127),
    .A2(n3154),
    .B1(n3157),
    .B2(n3153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3126));
 sky130_fd_sc_hd__o221a_1 U3493 (.A1(n3127),
    .A2(n3154),
    .B1(n3157),
    .B2(n3153),
    .C1(n3126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3128));
 sky130_fd_sc_hd__inv_2 U3494 (.A(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3159));
 sky130_fd_sc_hd__a22o_1 U3495 (.A1(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ),
    .A2(n3159),
    .B1(n3183),
    .B2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3163));
 sky130_fd_sc_hd__o2111a_1 U3496 (.A1(n3158),
    .A2(n3152),
    .B1(n3129),
    .C1(n3128),
    .D1(n3163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3130));
 sky130_fd_sc_hd__or2_1 U3497 (.A(n3304),
    .B(n3194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3134));
 sky130_fd_sc_hd__inv_2 U3498 (.A(n3134),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3138));
 sky130_fd_sc_hd__a22o_1 U3499 (.A1(n3130),
    .A2(n3138),
    .B1(n_TX_FULL_FLAG_FLAG_),
    .B2(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2139));
 sky130_fd_sc_hd__inv_1 U3500 (.A(\ICR_REG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3131));
 sky130_fd_sc_hd__a21o_1 U3501 (.A1(n3131),
    .A2(\RIS_REG[5] ),
    .B1(n_TX_FULL_FLAG_FLAG_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2138));
 sky130_fd_sc_hd__inv_2 U3502 (.A(n3194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3155));
 sky130_fd_sc_hd__or2_1 U3503 (.A(n3155),
    .B(net209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3133));
 sky130_fd_sc_hd__inv_2 U3504 (.A(n3133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3166));
 sky130_fd_sc_hd__o21a_1 U3505 (.A1(n3166),
    .A2(n3138),
    .B1(n3143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3132));
 sky130_fd_sc_hd__a31o_1 U3506 (.A1(n3133),
    .A2(n3134),
    .A3(\TXFIFOLEVEL_REG[0] ),
    .B1(n3132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2137));
 sky130_fd_sc_hd__inv_2 U3507 (.A(\TXFIFOLEVEL_REG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3142));
 sky130_fd_sc_hd__a22o_1 U3508 (.A1(\TXFIFOLEVEL_REG[0] ),
    .A2(n3134),
    .B1(n3143),
    .B2(n3133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3135));
 sky130_fd_sc_hd__mux2_1 U3509 (.A0(n3142),
    .A1(\TXFIFOLEVEL_REG[1] ),
    .S(n3135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2136));
 sky130_fd_sc_hd__and3_1 U3510 (.A(n3138),
    .B(\TXFIFOLEVEL_REG[0] ),
    .C(\TXFIFOLEVEL_REG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3136));
 sky130_fd_sc_hd__a31o_1 U3511 (.A1(n3166),
    .A2(n3143),
    .A3(n3142),
    .B1(\TXFIFOLEVEL_REG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3141));
 sky130_fd_sc_hd__inv_2 U3512 (.A(\TXFIFOLEVEL_REG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3146));
 sky130_fd_sc_hd__a221o_1 U3513 (.A1(\TXFIFOLEVEL_REG[1] ),
    .A2(n3166),
    .B1(n3142),
    .B2(n3138),
    .C1(n3135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3137));
 sky130_fd_sc_hd__o22a_1 U3514 (.A1(n3136),
    .A2(n3141),
    .B1(n3146),
    .B2(n3137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2135));
 sky130_fd_sc_hd__inv_2 U3515 (.A(\TXFIFOLEVEL_REG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3149));
 sky130_fd_sc_hd__a31o_1 U3516 (.A1(\TXFIFOLEVEL_REG[0] ),
    .A2(n3138),
    .A3(\TXFIFOLEVEL_REG[1] ),
    .B1(n3146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3140));
 sky130_fd_sc_hd__a221o_1 U3517 (.A1(\TXFIFOLEVEL_REG[2] ),
    .A2(n3166),
    .B1(n3146),
    .B2(n3138),
    .C1(n3137),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3139));
 sky130_fd_sc_hd__a32o_1 U3518 (.A1(n3149),
    .A2(n3141),
    .A3(n3140),
    .B1(\TXFIFOLEVEL_REG[3] ),
    .B2(n3139),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2134));
 sky130_fd_sc_hd__or2_1 U3519 (.A(n3149),
    .B(\tx_fifo_th[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3151));
 sky130_fd_sc_hd__or2_1 U3520 (.A(\tx_fifo_th[1] ),
    .B(n3142),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3144));
 sky130_fd_sc_hd__a32o_1 U3521 (.A1(n3144),
    .A2(n3143),
    .A3(\tx_fifo_th[0] ),
    .B1(n3142),
    .B2(\tx_fifo_th[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3147));
 sky130_fd_sc_hd__or2_1 U3522 (.A(n3147),
    .B(n3146),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3145));
 sky130_fd_sc_hd__a22o_1 U3523 (.A1(n3147),
    .A2(n3146),
    .B1(\tx_fifo_th[2] ),
    .B2(n3145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3150));
 sky130_fd_sc_hd__nor2b_1 U3524 (.A(\ICR_REG[1] ),
    .B_N(\RIS_REG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3148));
 sky130_fd_sc_hd__a221o_1 U3525 (.A1(n3151),
    .A2(n3150),
    .B1(\tx_fifo_th[3] ),
    .B2(n3149),
    .C1(n3148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2133));
 sky130_fd_sc_hd__a22o_1 U3526 (.A1(n3155),
    .A2(n3183),
    .B1(n3194),
    .B2(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2132));
 sky130_fd_sc_hd__a22o_1 U3527 (.A1(n3155),
    .A2(n3152),
    .B1(n3194),
    .B2(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2131));
 sky130_fd_sc_hd__a22o_1 U3528 (.A1(n3155),
    .A2(n3153),
    .B1(n3194),
    .B2(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2130));
 sky130_fd_sc_hd__a22o_1 U3529 (.A1(n3155),
    .A2(n3154),
    .B1(n3194),
    .B2(\inst_to_wrap_tx_fifo_w_ptr_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2129));
 sky130_fd_sc_hd__a22o_1 U3530 (.A1(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ),
    .B1(n3159),
    .B2(n3158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3168));
 sky130_fd_sc_hd__nor2_1 U3531 (.A(n3159),
    .B(n3158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3156));
 sky130_fd_sc_hd__mux2_1 U3532 (.A0(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ),
    .A1(n3157),
    .S(n3156),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3169));
 sky130_fd_sc_hd__or3_1 U3533 (.A(n3159),
    .B(n3158),
    .C(n3157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3160));
 sky130_fd_sc_hd__a22o_1 U3534 (.A1(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A2(n3289),
    .B1(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ),
    .B2(n3160),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3170));
 sky130_fd_sc_hd__a22oi_1 U3535 (.A1(n3193),
    .A2(n3170),
    .B1(n3190),
    .B2(n3169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3161));
 sky130_fd_sc_hd__o221a_1 U3536 (.A1(n3190),
    .A2(n3169),
    .B1(n3193),
    .B2(n3170),
    .C1(n3161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3164));
 sky130_fd_sc_hd__nand2_1 U3537 (.A(n3168),
    .B(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3162));
 sky130_fd_sc_hd__o2111a_1 U3538 (.A1(n3168),
    .A2(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .B1(n3164),
    .C1(n3163),
    .D1(n3162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3165));
 sky130_fd_sc_hd__a22o_1 U3539 (.A1(n_TX_EMPTY_FLAG_FLAG_),
    .A2(n3194),
    .B1(n3166),
    .B2(n3165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2128));
 sky130_fd_sc_hd__inv_1 U3540 (.A(\ICR_REG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3167));
 sky130_fd_sc_hd__a21o_1 U3541 (.A1(\RIS_REG[0] ),
    .A2(n3167),
    .B1(n_TX_EMPTY_FLAG_FLAG_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2127));
 sky130_fd_sc_hd__a22o_1 U3542 (.A1(n3304),
    .A2(n3169),
    .B1(net209),
    .B2(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2125));
 sky130_fd_sc_hd__a22o_1 U3543 (.A1(n3304),
    .A2(n3170),
    .B1(net209),
    .B2(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2124));
 sky130_fd_sc_hd__or2_1 U3544 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .B(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3197));
 sky130_fd_sc_hd__or3_1 U3545 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ),
    .B(\inst_to_wrap_tx_fifo_w_ptr_reg[3] ),
    .C(n3194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3186));
 sky130_fd_sc_hd__or2_4 U3546 (.A(n3197),
    .B(n3186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3171));
 sky130_fd_sc_hd__clkinv_2 U3547 (.A(n3171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3172));
 sky130_fd_sc_hd__a22o_1 U3548 (.A1(n3172),
    .A2(net237),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2123));
 sky130_fd_sc_hd__a22o_1 U3549 (.A1(n3172),
    .A2(net27),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2122));
 sky130_fd_sc_hd__a22o_1 U3550 (.A1(n3172),
    .A2(net26),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2121));
 sky130_fd_sc_hd__a22o_1 U3551 (.A1(n3172),
    .A2(net232),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2120));
 sky130_fd_sc_hd__a22o_1 U3552 (.A1(n3172),
    .A2(net233),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2119));
 sky130_fd_sc_hd__a22o_1 U3553 (.A1(n3172),
    .A2(net234),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2118));
 sky130_fd_sc_hd__a22o_1 U3554 (.A1(n3172),
    .A2(net235),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2117));
 sky130_fd_sc_hd__a22o_1 U3555 (.A1(n3172),
    .A2(net236),
    .B1(n3171),
    .B2(\inst_to_wrap_tx_fifo_array_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2116));
 sky130_fd_sc_hd__nor2_1 U3556 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[3] ),
    .B(n3194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3182));
 sky130_fd_sc_hd__or3b_4 U3557 (.A(n3183),
    .B(n3197),
    .C_N(n3182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3173));
 sky130_fd_sc_hd__clkinv_2 U3558 (.A(n3173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3174));
 sky130_fd_sc_hd__a22o_1 U3559 (.A1(n3174),
    .A2(net237),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2115));
 sky130_fd_sc_hd__a22o_1 U3560 (.A1(n3174),
    .A2(net27),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2114));
 sky130_fd_sc_hd__a22o_1 U3561 (.A1(n3174),
    .A2(net26),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2113));
 sky130_fd_sc_hd__a22o_1 U3562 (.A1(n3174),
    .A2(net25),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2112));
 sky130_fd_sc_hd__a22o_1 U3563 (.A1(n3174),
    .A2(net24),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2111));
 sky130_fd_sc_hd__a22o_1 U3564 (.A1(n3174),
    .A2(net234),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2110));
 sky130_fd_sc_hd__a22o_1 U3565 (.A1(n3174),
    .A2(net235),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2109));
 sky130_fd_sc_hd__a22o_1 U3566 (.A1(n3174),
    .A2(net21),
    .B1(n3173),
    .B2(\inst_to_wrap_tx_fifo_array_reg[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2108));
 sky130_fd_sc_hd__nand2_1 U3567 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .B(n3190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3202));
 sky130_fd_sc_hd__or2_4 U3568 (.A(n3186),
    .B(n3202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3175));
 sky130_fd_sc_hd__clkinv_2 U3569 (.A(n3175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3176));
 sky130_fd_sc_hd__a22o_1 U3570 (.A1(n3176),
    .A2(net237),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2107));
 sky130_fd_sc_hd__a22o_1 U3571 (.A1(n3176),
    .A2(net27),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2106));
 sky130_fd_sc_hd__a22o_1 U3572 (.A1(n3176),
    .A2(net26),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2105));
 sky130_fd_sc_hd__a22o_1 U3573 (.A1(n3176),
    .A2(net232),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2104));
 sky130_fd_sc_hd__a22o_1 U3574 (.A1(n3176),
    .A2(net233),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2103));
 sky130_fd_sc_hd__a22o_1 U3575 (.A1(n3176),
    .A2(net234),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2102));
 sky130_fd_sc_hd__a22o_1 U3576 (.A1(n3176),
    .A2(net235),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2101));
 sky130_fd_sc_hd__a22o_1 U3577 (.A1(n3176),
    .A2(net236),
    .B1(n3175),
    .B2(\inst_to_wrap_tx_fifo_array_reg[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2100));
 sky130_fd_sc_hd__or3_1 U3578 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[3] ),
    .B(n3194),
    .C(n3177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3189));
 sky130_fd_sc_hd__or2_4 U3579 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ),
    .B(n3189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3178));
 sky130_fd_sc_hd__clkinv_2 U3580 (.A(n3178),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3179));
 sky130_fd_sc_hd__a22o_1 U3581 (.A1(n3179),
    .A2(net20),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2099));
 sky130_fd_sc_hd__a22o_1 U3582 (.A1(n3179),
    .A2(net27),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2098));
 sky130_fd_sc_hd__a22o_1 U3583 (.A1(n3179),
    .A2(net26),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2097));
 sky130_fd_sc_hd__a22o_1 U3584 (.A1(n3179),
    .A2(net232),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2096));
 sky130_fd_sc_hd__a22o_1 U3585 (.A1(n3179),
    .A2(net233),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2095));
 sky130_fd_sc_hd__a22o_1 U3586 (.A1(n3179),
    .A2(net23),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2094));
 sky130_fd_sc_hd__a22o_1 U3587 (.A1(n3179),
    .A2(net22),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2093));
 sky130_fd_sc_hd__a22o_1 U3588 (.A1(n3179),
    .A2(net236),
    .B1(n3178),
    .B2(\inst_to_wrap_tx_fifo_array_reg[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2092));
 sky130_fd_sc_hd__or2_1 U3589 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .B(n3190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3207));
 sky130_fd_sc_hd__or2_4 U3590 (.A(n3186),
    .B(n3207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3180));
 sky130_fd_sc_hd__clkinv_2 U3591 (.A(n3180),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3181));
 sky130_fd_sc_hd__a22o_1 U3592 (.A1(n3181),
    .A2(net237),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2091));
 sky130_fd_sc_hd__a22o_1 U3593 (.A1(n3181),
    .A2(net27),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2090));
 sky130_fd_sc_hd__a22o_1 U3594 (.A1(n3181),
    .A2(net26),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2089));
 sky130_fd_sc_hd__a22o_1 U3595 (.A1(n3181),
    .A2(net232),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2088));
 sky130_fd_sc_hd__a22o_1 U3596 (.A1(n3181),
    .A2(net233),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2087));
 sky130_fd_sc_hd__a22o_1 U3597 (.A1(n3181),
    .A2(net234),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2086));
 sky130_fd_sc_hd__a22o_1 U3598 (.A1(n3181),
    .A2(net235),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2085));
 sky130_fd_sc_hd__a22o_1 U3599 (.A1(n3181),
    .A2(net236),
    .B1(n3180),
    .B2(\inst_to_wrap_tx_fifo_array_reg[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2084));
 sky130_fd_sc_hd__or3b_4 U3600 (.A(n3183),
    .B(n3207),
    .C_N(n3182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3184));
 sky130_fd_sc_hd__clkinv_2 U3601 (.A(n3184),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3185));
 sky130_fd_sc_hd__a22o_1 U3602 (.A1(n3185),
    .A2(net237),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2083));
 sky130_fd_sc_hd__a22o_1 U3603 (.A1(n3185),
    .A2(net27),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2082));
 sky130_fd_sc_hd__a22o_1 U3604 (.A1(n3185),
    .A2(net26),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2081));
 sky130_fd_sc_hd__a22o_1 U3605 (.A1(n3185),
    .A2(net25),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2080));
 sky130_fd_sc_hd__a22o_1 U3606 (.A1(n3185),
    .A2(net24),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2079));
 sky130_fd_sc_hd__a22o_1 U3607 (.A1(n3185),
    .A2(net234),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2078));
 sky130_fd_sc_hd__a22o_1 U3608 (.A1(n3185),
    .A2(net235),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2077));
 sky130_fd_sc_hd__a22o_1 U3609 (.A1(n3185),
    .A2(net21),
    .B1(n3184),
    .B2(\inst_to_wrap_tx_fifo_array_reg[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2076));
 sky130_fd_sc_hd__nand2_1 U3610 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ),
    .B(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3212));
 sky130_fd_sc_hd__or2_4 U3611 (.A(n3212),
    .B(n3186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3187));
 sky130_fd_sc_hd__clkinv_2 U3612 (.A(n3187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3188));
 sky130_fd_sc_hd__a22o_1 U3613 (.A1(n3188),
    .A2(net237),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2075));
 sky130_fd_sc_hd__a22o_1 U3614 (.A1(n3188),
    .A2(net27),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2074));
 sky130_fd_sc_hd__a22o_1 U3615 (.A1(n3188),
    .A2(net26),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2073));
 sky130_fd_sc_hd__a22o_1 U3616 (.A1(n3188),
    .A2(net232),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2072));
 sky130_fd_sc_hd__a22o_1 U3617 (.A1(n3188),
    .A2(net233),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2071));
 sky130_fd_sc_hd__a22o_1 U3618 (.A1(n3188),
    .A2(net234),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2070));
 sky130_fd_sc_hd__a22o_1 U3619 (.A1(n3188),
    .A2(net235),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2069));
 sky130_fd_sc_hd__a22o_1 U3620 (.A1(n3188),
    .A2(net236),
    .B1(n3187),
    .B2(\inst_to_wrap_tx_fifo_array_reg[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2068));
 sky130_fd_sc_hd__or2_4 U3621 (.A(n3190),
    .B(n3189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3191));
 sky130_fd_sc_hd__clkinv_2 U3622 (.A(n3191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3192));
 sky130_fd_sc_hd__a22o_1 U3623 (.A1(n3192),
    .A2(net20),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2067));
 sky130_fd_sc_hd__a22o_1 U3624 (.A1(n3192),
    .A2(net27),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2066));
 sky130_fd_sc_hd__a22o_1 U3625 (.A1(n3192),
    .A2(net26),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2065));
 sky130_fd_sc_hd__a22o_1 U3626 (.A1(n3192),
    .A2(net232),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2064));
 sky130_fd_sc_hd__a22o_1 U3627 (.A1(n3192),
    .A2(net233),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2063));
 sky130_fd_sc_hd__a22o_1 U3628 (.A1(n3192),
    .A2(net23),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2062));
 sky130_fd_sc_hd__a22o_1 U3629 (.A1(n3192),
    .A2(net22),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2061));
 sky130_fd_sc_hd__a22o_1 U3630 (.A1(n3192),
    .A2(net236),
    .B1(n3191),
    .B2(\inst_to_wrap_tx_fifo_array_reg[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2060));
 sky130_fd_sc_hd__or3_2 U3631 (.A(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ),
    .B(n3194),
    .C(n3193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3211));
 sky130_fd_sc_hd__or2_4 U3632 (.A(n3197),
    .B(n3211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3195));
 sky130_fd_sc_hd__clkinv_2 U3633 (.A(n3195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3196));
 sky130_fd_sc_hd__a22o_1 U3634 (.A1(n3196),
    .A2(net237),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2059));
 sky130_fd_sc_hd__a22o_1 U3635 (.A1(n3196),
    .A2(net27),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2058));
 sky130_fd_sc_hd__a22o_1 U3636 (.A1(n3196),
    .A2(net26),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2057));
 sky130_fd_sc_hd__a22o_1 U3637 (.A1(n3196),
    .A2(net232),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2056));
 sky130_fd_sc_hd__a22o_1 U3638 (.A1(n3196),
    .A2(net233),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2055));
 sky130_fd_sc_hd__a22o_1 U3639 (.A1(n3196),
    .A2(net234),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2054));
 sky130_fd_sc_hd__a22o_1 U3640 (.A1(n3196),
    .A2(net235),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2053));
 sky130_fd_sc_hd__a22o_1 U3641 (.A1(n3196),
    .A2(net236),
    .B1(n3195),
    .B2(\inst_to_wrap_tx_fifo_array_reg[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2052));
 sky130_fd_sc_hd__or2_4 U3642 (.A(n3208),
    .B(n3197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3198));
 sky130_fd_sc_hd__clkinv_2 U3643 (.A(n3198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3199));
 sky130_fd_sc_hd__a22o_1 U3644 (.A1(n3199),
    .A2(net237),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2051));
 sky130_fd_sc_hd__a22o_1 U3645 (.A1(n3199),
    .A2(net27),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2050));
 sky130_fd_sc_hd__a22o_1 U3646 (.A1(n3199),
    .A2(net26),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2049));
 sky130_fd_sc_hd__a22o_1 U3647 (.A1(n3199),
    .A2(net232),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2048));
 sky130_fd_sc_hd__a22o_1 U3648 (.A1(n3199),
    .A2(net233),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2047));
 sky130_fd_sc_hd__a22o_1 U3649 (.A1(n3199),
    .A2(net234),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2046));
 sky130_fd_sc_hd__a22o_1 U3650 (.A1(n3199),
    .A2(net235),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2045));
 sky130_fd_sc_hd__a22o_1 U3651 (.A1(n3199),
    .A2(net236),
    .B1(n3198),
    .B2(\inst_to_wrap_tx_fifo_array_reg[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2044));
 sky130_fd_sc_hd__or2_4 U3652 (.A(n3202),
    .B(n3211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3200));
 sky130_fd_sc_hd__clkinv_2 U3653 (.A(n3200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3201));
 sky130_fd_sc_hd__a22o_1 U3654 (.A1(n3201),
    .A2(net237),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2043));
 sky130_fd_sc_hd__a22o_1 U3655 (.A1(n3201),
    .A2(net27),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2042));
 sky130_fd_sc_hd__a22o_1 U3656 (.A1(n3201),
    .A2(net26),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2041));
 sky130_fd_sc_hd__a22o_1 U3657 (.A1(n3201),
    .A2(net232),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2040));
 sky130_fd_sc_hd__a22o_1 U3658 (.A1(n3201),
    .A2(net233),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2039));
 sky130_fd_sc_hd__a22o_1 U3659 (.A1(n3201),
    .A2(net234),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2038));
 sky130_fd_sc_hd__a22o_1 U3660 (.A1(n3201),
    .A2(net235),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2037));
 sky130_fd_sc_hd__a22o_1 U3661 (.A1(n3201),
    .A2(net236),
    .B1(n3200),
    .B2(\inst_to_wrap_tx_fifo_array_reg[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2036));
 sky130_fd_sc_hd__or2_4 U3662 (.A(n3208),
    .B(n3202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3203));
 sky130_fd_sc_hd__clkinv_2 U3663 (.A(n3203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3204));
 sky130_fd_sc_hd__a22o_1 U3664 (.A1(n3204),
    .A2(net237),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2035));
 sky130_fd_sc_hd__a22o_1 U3665 (.A1(n3204),
    .A2(net27),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2034));
 sky130_fd_sc_hd__a22o_1 U3666 (.A1(n3204),
    .A2(net26),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2033));
 sky130_fd_sc_hd__a22o_1 U3667 (.A1(n3204),
    .A2(net232),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2032));
 sky130_fd_sc_hd__a22o_1 U3668 (.A1(n3204),
    .A2(net233),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2031));
 sky130_fd_sc_hd__a22o_1 U3669 (.A1(n3204),
    .A2(net234),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2030));
 sky130_fd_sc_hd__a22o_1 U3670 (.A1(n3204),
    .A2(net235),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2029));
 sky130_fd_sc_hd__a22o_1 U3671 (.A1(n3204),
    .A2(net236),
    .B1(n3203),
    .B2(\inst_to_wrap_tx_fifo_array_reg[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2028));
 sky130_fd_sc_hd__or2_4 U3672 (.A(n3207),
    .B(n3211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3205));
 sky130_fd_sc_hd__clkinv_2 U3673 (.A(n3205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3206));
 sky130_fd_sc_hd__a22o_1 U3674 (.A1(n3206),
    .A2(net237),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2027));
 sky130_fd_sc_hd__a22o_1 U3675 (.A1(n3206),
    .A2(net27),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2026));
 sky130_fd_sc_hd__a22o_1 U3676 (.A1(n3206),
    .A2(net26),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2025));
 sky130_fd_sc_hd__a22o_1 U3677 (.A1(n3206),
    .A2(net232),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2024));
 sky130_fd_sc_hd__a22o_1 U3678 (.A1(n3206),
    .A2(net233),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2023));
 sky130_fd_sc_hd__a22o_1 U3679 (.A1(n3206),
    .A2(net234),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2022));
 sky130_fd_sc_hd__a22o_1 U3680 (.A1(n3206),
    .A2(net235),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2021));
 sky130_fd_sc_hd__a22o_1 U3681 (.A1(n3206),
    .A2(net236),
    .B1(n3205),
    .B2(\inst_to_wrap_tx_fifo_array_reg[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2020));
 sky130_fd_sc_hd__or2_4 U3682 (.A(n3208),
    .B(n3207),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3209));
 sky130_fd_sc_hd__clkinv_2 U3683 (.A(n3209),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3210));
 sky130_fd_sc_hd__a22o_1 U3684 (.A1(n3210),
    .A2(net237),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2019));
 sky130_fd_sc_hd__a22o_1 U3685 (.A1(n3210),
    .A2(net27),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2018));
 sky130_fd_sc_hd__a22o_1 U3686 (.A1(n3210),
    .A2(net26),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2017));
 sky130_fd_sc_hd__a22o_1 U3687 (.A1(n3210),
    .A2(net232),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2016));
 sky130_fd_sc_hd__a22o_1 U3688 (.A1(n3210),
    .A2(net233),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2015));
 sky130_fd_sc_hd__a22o_1 U3689 (.A1(n3210),
    .A2(net234),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2014));
 sky130_fd_sc_hd__a22o_1 U3690 (.A1(n3210),
    .A2(net235),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2013));
 sky130_fd_sc_hd__a22o_1 U3691 (.A1(n3210),
    .A2(net236),
    .B1(n3209),
    .B2(\inst_to_wrap_tx_fifo_array_reg[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2012));
 sky130_fd_sc_hd__or2_4 U3692 (.A(n3212),
    .B(n3211),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3213));
 sky130_fd_sc_hd__clkinv_2 U3693 (.A(n3213),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3214));
 sky130_fd_sc_hd__a22o_1 U3694 (.A1(n3214),
    .A2(net237),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2011));
 sky130_fd_sc_hd__a22o_1 U3695 (.A1(n3214),
    .A2(net27),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2010));
 sky130_fd_sc_hd__a22o_1 U3696 (.A1(n3214),
    .A2(net26),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2009));
 sky130_fd_sc_hd__a22o_1 U3697 (.A1(n3214),
    .A2(net232),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2008));
 sky130_fd_sc_hd__a22o_1 U3698 (.A1(n3214),
    .A2(net233),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2007));
 sky130_fd_sc_hd__a22o_1 U3699 (.A1(n3214),
    .A2(net234),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2006));
 sky130_fd_sc_hd__a22o_1 U3700 (.A1(n3214),
    .A2(net235),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2005));
 sky130_fd_sc_hd__a22o_1 U3701 (.A1(n3214),
    .A2(net236),
    .B1(n3213),
    .B2(\inst_to_wrap_tx_fifo_array_reg[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2004));
 sky130_fd_sc_hd__a22o_1 U3702 (.A1(n3216),
    .A2(net237),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2003));
 sky130_fd_sc_hd__a22o_1 U3703 (.A1(n3216),
    .A2(net26),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2002));
 sky130_fd_sc_hd__a22o_1 U3704 (.A1(n3216),
    .A2(net232),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2001));
 sky130_fd_sc_hd__a22o_1 U3705 (.A1(n3216),
    .A2(net233),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n2000));
 sky130_fd_sc_hd__a22o_1 U3706 (.A1(n3216),
    .A2(net234),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1999));
 sky130_fd_sc_hd__a22o_1 U3707 (.A1(n3216),
    .A2(net235),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1998));
 sky130_fd_sc_hd__a22o_1 U3708 (.A1(n3216),
    .A2(net236),
    .B1(n3215),
    .B2(\inst_to_wrap_tx_fifo_array_reg[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1997));
 sky130_fd_sc_hd__a22o_1 U3709 (.A1(\inst_to_wrap_tx_fifo_array_reg[14] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[46] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3220));
 sky130_fd_sc_hd__a22o_1 U3710 (.A1(\inst_to_wrap_tx_fifo_array_reg[30] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[62] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3219));
 sky130_fd_sc_hd__a22o_1 U3711 (.A1(\inst_to_wrap_tx_fifo_array_reg[78] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[110] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3218));
 sky130_fd_sc_hd__a22o_1 U3712 (.A1(\inst_to_wrap_tx_fifo_array_reg[94] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[126] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3217));
 sky130_fd_sc_hd__or4_1 U3713 (.A(n3220),
    .B(n3219),
    .C(n3218),
    .D(n3217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3227));
 sky130_fd_sc_hd__a22o_1 U3714 (.A1(\inst_to_wrap_tx_fifo_array_reg[6] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[38] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3224));
 sky130_fd_sc_hd__a22o_1 U3715 (.A1(\inst_to_wrap_tx_fifo_array_reg[22] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[54] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3223));
 sky130_fd_sc_hd__a22o_1 U3716 (.A1(\inst_to_wrap_tx_fifo_array_reg[70] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[102] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3222));
 sky130_fd_sc_hd__a22o_1 U3717 (.A1(\inst_to_wrap_tx_fifo_array_reg[86] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[118] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3221));
 sky130_fd_sc_hd__or4_1 U3718 (.A(n3224),
    .B(n3223),
    .C(n3222),
    .D(n3221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3225));
 sky130_fd_sc_hd__a22o_1 U3719 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[6] ),
    .A2(net209),
    .B1(n3300),
    .B2(n3225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3226));
 sky130_fd_sc_hd__a31o_1 U3720 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n3227),
    .B1(n3226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1996));
 sky130_fd_sc_hd__a22o_1 U3721 (.A1(n3306),
    .A2(net120),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1995));
 sky130_fd_sc_hd__a22o_1 U3722 (.A1(n3308),
    .A2(net120),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1994));
 sky130_fd_sc_hd__a22o_1 U3723 (.A1(n3310),
    .A2(net120),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1993));
 sky130_fd_sc_hd__a22o_1 U3724 (.A1(n3312),
    .A2(net120),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1992));
 sky130_fd_sc_hd__a22o_1 U3725 (.A1(n3314),
    .A2(net111),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1991));
 sky130_fd_sc_hd__a22o_1 U3726 (.A1(n3316),
    .A2(net111),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1990));
 sky130_fd_sc_hd__a22o_1 U3727 (.A1(n3318),
    .A2(net120),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1989));
 sky130_fd_sc_hd__a22o_1 U3728 (.A1(n3320),
    .A2(net120),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1988));
 sky130_fd_sc_hd__a22o_1 U3729 (.A1(n3322),
    .A2(net120),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1987));
 sky130_fd_sc_hd__a22o_1 U3730 (.A1(\inst_to_wrap_tx_fifo_array_reg[13] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[45] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3231));
 sky130_fd_sc_hd__a22o_1 U3731 (.A1(\inst_to_wrap_tx_fifo_array_reg[29] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[61] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3230));
 sky130_fd_sc_hd__a22o_1 U3732 (.A1(\inst_to_wrap_tx_fifo_array_reg[77] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[109] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3229));
 sky130_fd_sc_hd__a22o_1 U3733 (.A1(\inst_to_wrap_tx_fifo_array_reg[93] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[125] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3228));
 sky130_fd_sc_hd__or4_1 U3734 (.A(n3231),
    .B(n3230),
    .C(n3229),
    .D(n3228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3238));
 sky130_fd_sc_hd__a22o_1 U3735 (.A1(\inst_to_wrap_tx_fifo_array_reg[5] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[37] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3235));
 sky130_fd_sc_hd__a22o_1 U3736 (.A1(\inst_to_wrap_tx_fifo_array_reg[21] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[53] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3234));
 sky130_fd_sc_hd__a22o_1 U3737 (.A1(\inst_to_wrap_tx_fifo_array_reg[69] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[101] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3233));
 sky130_fd_sc_hd__a22o_1 U3738 (.A1(\inst_to_wrap_tx_fifo_array_reg[85] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[117] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3232));
 sky130_fd_sc_hd__or4_1 U3739 (.A(n3235),
    .B(n3234),
    .C(n3233),
    .D(n3232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3236));
 sky130_fd_sc_hd__a22o_1 U3740 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[5] ),
    .A2(net209),
    .B1(n3300),
    .B2(n3236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3237));
 sky130_fd_sc_hd__a31o_1 U3741 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n3238),
    .B1(n3237),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1986));
 sky130_fd_sc_hd__a22o_1 U3742 (.A1(n3306),
    .A2(net100),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1985));
 sky130_fd_sc_hd__a22o_1 U3743 (.A1(n3308),
    .A2(net106),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1984));
 sky130_fd_sc_hd__a22o_1 U3744 (.A1(n3310),
    .A2(net106),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1983));
 sky130_fd_sc_hd__a22o_1 U3745 (.A1(n3312),
    .A2(net100),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1982));
 sky130_fd_sc_hd__a22o_1 U3746 (.A1(n3314),
    .A2(net106),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1981));
 sky130_fd_sc_hd__a22o_1 U3747 (.A1(n3316),
    .A2(net106),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1980));
 sky130_fd_sc_hd__a22o_1 U3748 (.A1(n3318),
    .A2(net106),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1979));
 sky130_fd_sc_hd__a22o_1 U3749 (.A1(n3320),
    .A2(net106),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1978));
 sky130_fd_sc_hd__a22o_1 U3750 (.A1(n3322),
    .A2(net106),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1977));
 sky130_fd_sc_hd__a22o_1 U3751 (.A1(\inst_to_wrap_tx_fifo_array_reg[12] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[44] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3242));
 sky130_fd_sc_hd__a22o_1 U3752 (.A1(\inst_to_wrap_tx_fifo_array_reg[28] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[60] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3241));
 sky130_fd_sc_hd__a22o_1 U3753 (.A1(\inst_to_wrap_tx_fifo_array_reg[76] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[108] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3240));
 sky130_fd_sc_hd__a22o_1 U3754 (.A1(\inst_to_wrap_tx_fifo_array_reg[92] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[124] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3239));
 sky130_fd_sc_hd__or4_1 U3755 (.A(n3242),
    .B(n3241),
    .C(n3240),
    .D(n3239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3249));
 sky130_fd_sc_hd__a22o_1 U3756 (.A1(\inst_to_wrap_tx_fifo_array_reg[4] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[36] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3246));
 sky130_fd_sc_hd__a22o_1 U3757 (.A1(\inst_to_wrap_tx_fifo_array_reg[20] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[52] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3245));
 sky130_fd_sc_hd__a22o_1 U3758 (.A1(\inst_to_wrap_tx_fifo_array_reg[68] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[100] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3244));
 sky130_fd_sc_hd__a22o_1 U3759 (.A1(\inst_to_wrap_tx_fifo_array_reg[84] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[116] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3243));
 sky130_fd_sc_hd__or4_1 U3760 (.A(n3246),
    .B(n3245),
    .C(n3244),
    .D(n3243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3247));
 sky130_fd_sc_hd__a22o_1 U3761 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[4] ),
    .A2(net209),
    .B1(n3300),
    .B2(n3247),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3248));
 sky130_fd_sc_hd__a31o_1 U3762 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n3249),
    .B1(n3248),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1976));
 sky130_fd_sc_hd__a22o_1 U3763 (.A1(n3306),
    .A2(net79),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1975));
 sky130_fd_sc_hd__a22o_1 U3764 (.A1(n3308),
    .A2(net84),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1974));
 sky130_fd_sc_hd__a22o_1 U3765 (.A1(n3310),
    .A2(net84),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1973));
 sky130_fd_sc_hd__a22o_1 U3766 (.A1(n3312),
    .A2(net84),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1972));
 sky130_fd_sc_hd__a22o_1 U3767 (.A1(n3314),
    .A2(net84),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1971));
 sky130_fd_sc_hd__a22o_1 U3768 (.A1(n3316),
    .A2(net84),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1970));
 sky130_fd_sc_hd__a22o_1 U3769 (.A1(n3318),
    .A2(net79),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1969));
 sky130_fd_sc_hd__a22o_1 U3770 (.A1(n3320),
    .A2(net84),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1968));
 sky130_fd_sc_hd__a22o_1 U3771 (.A1(n3322),
    .A2(net84),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1967));
 sky130_fd_sc_hd__a22o_1 U3772 (.A1(\inst_to_wrap_tx_fifo_array_reg[11] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[43] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3253));
 sky130_fd_sc_hd__a22o_1 U3773 (.A1(\inst_to_wrap_tx_fifo_array_reg[27] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[59] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3252));
 sky130_fd_sc_hd__a22o_1 U3774 (.A1(\inst_to_wrap_tx_fifo_array_reg[75] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[107] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3251));
 sky130_fd_sc_hd__a22o_1 U3775 (.A1(\inst_to_wrap_tx_fifo_array_reg[91] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[123] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3250));
 sky130_fd_sc_hd__or4_1 U3776 (.A(n3253),
    .B(n3252),
    .C(n3251),
    .D(n3250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3260));
 sky130_fd_sc_hd__a22o_1 U3777 (.A1(\inst_to_wrap_tx_fifo_array_reg[3] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[35] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3257));
 sky130_fd_sc_hd__a22o_1 U3778 (.A1(\inst_to_wrap_tx_fifo_array_reg[19] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[51] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3256));
 sky130_fd_sc_hd__a22o_1 U3779 (.A1(\inst_to_wrap_tx_fifo_array_reg[67] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[99] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3255));
 sky130_fd_sc_hd__a22o_1 U3780 (.A1(\inst_to_wrap_tx_fifo_array_reg[83] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[115] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3254));
 sky130_fd_sc_hd__or4_1 U3781 (.A(n3257),
    .B(n3256),
    .C(n3255),
    .D(n3254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3258));
 sky130_fd_sc_hd__a22o_1 U3782 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[3] ),
    .A2(net209),
    .B1(n3300),
    .B2(n3258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3259));
 sky130_fd_sc_hd__a31o_1 U3783 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n3260),
    .B1(n3259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1966));
 sky130_fd_sc_hd__a22o_1 U3784 (.A1(n3306),
    .A2(net108),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1965));
 sky130_fd_sc_hd__a22o_1 U3785 (.A1(n3308),
    .A2(net116),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1964));
 sky130_fd_sc_hd__a22o_1 U3786 (.A1(n3310),
    .A2(net116),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1963));
 sky130_fd_sc_hd__a22o_1 U3787 (.A1(n3312),
    .A2(net116),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1962));
 sky130_fd_sc_hd__a22o_1 U3788 (.A1(n3314),
    .A2(net116),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1961));
 sky130_fd_sc_hd__a22o_1 U3789 (.A1(n3316),
    .A2(net116),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1960));
 sky130_fd_sc_hd__a22o_1 U3790 (.A1(n3318),
    .A2(net116),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1959));
 sky130_fd_sc_hd__a22o_1 U3791 (.A1(n3320),
    .A2(net108),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1958));
 sky130_fd_sc_hd__a22o_1 U3792 (.A1(n3322),
    .A2(net116),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1957));
 sky130_fd_sc_hd__a22o_1 U3793 (.A1(\inst_to_wrap_tx_fifo_array_reg[10] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[42] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3264));
 sky130_fd_sc_hd__a22o_1 U3794 (.A1(\inst_to_wrap_tx_fifo_array_reg[26] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[58] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3263));
 sky130_fd_sc_hd__a22o_1 U3795 (.A1(\inst_to_wrap_tx_fifo_array_reg[74] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[106] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3262));
 sky130_fd_sc_hd__a22o_1 U3796 (.A1(\inst_to_wrap_tx_fifo_array_reg[90] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[122] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3261));
 sky130_fd_sc_hd__or4_1 U3797 (.A(n3264),
    .B(n3263),
    .C(n3262),
    .D(n3261),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3271));
 sky130_fd_sc_hd__a22o_1 U3798 (.A1(\inst_to_wrap_tx_fifo_array_reg[2] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[34] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3268));
 sky130_fd_sc_hd__a22o_1 U3799 (.A1(\inst_to_wrap_tx_fifo_array_reg[18] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[50] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3267));
 sky130_fd_sc_hd__a22o_1 U3800 (.A1(\inst_to_wrap_tx_fifo_array_reg[66] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[98] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3266));
 sky130_fd_sc_hd__a22o_1 U3801 (.A1(\inst_to_wrap_tx_fifo_array_reg[82] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[114] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3265));
 sky130_fd_sc_hd__or4_1 U3802 (.A(n3268),
    .B(n3267),
    .C(n3266),
    .D(n3265),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3269));
 sky130_fd_sc_hd__a22o_1 U3803 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[2] ),
    .A2(net209),
    .B1(n3300),
    .B2(n3269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3270));
 sky130_fd_sc_hd__a31o_1 U3804 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n3271),
    .B1(n3270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1956));
 sky130_fd_sc_hd__a22o_1 U3805 (.A1(n3306),
    .A2(net136),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1955));
 sky130_fd_sc_hd__a22o_1 U3806 (.A1(n3308),
    .A2(net146),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1954));
 sky130_fd_sc_hd__a22o_1 U3807 (.A1(n3310),
    .A2(net146),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1953));
 sky130_fd_sc_hd__a22o_1 U3808 (.A1(n3312),
    .A2(net146),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1952));
 sky130_fd_sc_hd__a22o_1 U3809 (.A1(n3314),
    .A2(net146),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1951));
 sky130_fd_sc_hd__a22o_1 U3810 (.A1(n3316),
    .A2(net146),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1950));
 sky130_fd_sc_hd__a22o_1 U3811 (.A1(n3318),
    .A2(net146),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1949));
 sky130_fd_sc_hd__a22o_1 U3812 (.A1(n3320),
    .A2(net146),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1948));
 sky130_fd_sc_hd__a22o_1 U3813 (.A1(n3322),
    .A2(net136),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1947));
 sky130_fd_sc_hd__a22o_1 U3814 (.A1(\inst_to_wrap_tx_fifo_array_reg[9] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[41] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3275));
 sky130_fd_sc_hd__a22o_1 U3815 (.A1(\inst_to_wrap_tx_fifo_array_reg[25] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[57] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3274));
 sky130_fd_sc_hd__a22o_1 U3816 (.A1(\inst_to_wrap_tx_fifo_array_reg[73] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[105] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3273));
 sky130_fd_sc_hd__a22o_1 U3817 (.A1(\inst_to_wrap_tx_fifo_array_reg[89] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[121] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3272));
 sky130_fd_sc_hd__or4_1 U3818 (.A(n3275),
    .B(n3274),
    .C(n3273),
    .D(n3272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3282));
 sky130_fd_sc_hd__a22o_1 U3819 (.A1(\inst_to_wrap_tx_fifo_array_reg[1] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[33] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3279));
 sky130_fd_sc_hd__a22o_1 U3820 (.A1(\inst_to_wrap_tx_fifo_array_reg[17] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[49] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3278));
 sky130_fd_sc_hd__a22o_1 U3821 (.A1(\inst_to_wrap_tx_fifo_array_reg[65] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[97] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3277));
 sky130_fd_sc_hd__a22o_1 U3822 (.A1(\inst_to_wrap_tx_fifo_array_reg[81] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[113] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3276));
 sky130_fd_sc_hd__or4_1 U3823 (.A(n3279),
    .B(n3278),
    .C(n3277),
    .D(n3276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3280));
 sky130_fd_sc_hd__a22o_1 U3824 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[1] ),
    .A2(net209),
    .B1(n3300),
    .B2(n3280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3281));
 sky130_fd_sc_hd__a31o_1 U3825 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n3282),
    .B1(n3281),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1946));
 sky130_fd_sc_hd__a22o_1 U3826 (.A1(n3306),
    .A2(net134),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1945));
 sky130_fd_sc_hd__a22o_1 U3827 (.A1(n3308),
    .A2(net134),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1944));
 sky130_fd_sc_hd__a22o_1 U3828 (.A1(n3310),
    .A2(net134),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1943));
 sky130_fd_sc_hd__a22o_1 U3829 (.A1(n3312),
    .A2(net127),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1942));
 sky130_fd_sc_hd__a22o_1 U3830 (.A1(n3314),
    .A2(net134),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1941));
 sky130_fd_sc_hd__a22o_1 U3831 (.A1(n3316),
    .A2(net134),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1940));
 sky130_fd_sc_hd__a22o_1 U3832 (.A1(n3318),
    .A2(net134),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1939));
 sky130_fd_sc_hd__a22o_1 U3833 (.A1(n3320),
    .A2(net134),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1938));
 sky130_fd_sc_hd__a22o_1 U3834 (.A1(n3322),
    .A2(net127),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1937));
 sky130_fd_sc_hd__a22o_1 U3835 (.A1(\inst_to_wrap_tx_fifo_array_reg[8] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[40] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3286));
 sky130_fd_sc_hd__a22o_1 U3836 (.A1(\inst_to_wrap_tx_fifo_array_reg[24] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[56] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3285));
 sky130_fd_sc_hd__a22o_1 U3837 (.A1(\inst_to_wrap_tx_fifo_array_reg[72] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[104] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3284));
 sky130_fd_sc_hd__a22o_1 U3838 (.A1(\inst_to_wrap_tx_fifo_array_reg[88] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[120] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3283));
 sky130_fd_sc_hd__or4_1 U3839 (.A(n3286),
    .B(n3285),
    .C(n3284),
    .D(n3283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3303));
 sky130_fd_sc_hd__a22o_1 U3840 (.A1(\inst_to_wrap_tx_fifo_array_reg[0] ),
    .A2(n3288),
    .B1(\inst_to_wrap_tx_fifo_array_reg[32] ),
    .B2(n3287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3298));
 sky130_fd_sc_hd__a22o_1 U3841 (.A1(\inst_to_wrap_tx_fifo_array_reg[16] ),
    .A2(n3290),
    .B1(\inst_to_wrap_tx_fifo_array_reg[48] ),
    .B2(net206),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3297));
 sky130_fd_sc_hd__a22o_1 U3842 (.A1(\inst_to_wrap_tx_fifo_array_reg[64] ),
    .A2(n3292),
    .B1(\inst_to_wrap_tx_fifo_array_reg[96] ),
    .B2(n3291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3296));
 sky130_fd_sc_hd__a22o_1 U3843 (.A1(\inst_to_wrap_tx_fifo_array_reg[80] ),
    .A2(n3294),
    .B1(\inst_to_wrap_tx_fifo_array_reg[112] ),
    .B2(n3293),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3295));
 sky130_fd_sc_hd__or4_1 U3844 (.A(n3298),
    .B(n3297),
    .C(n3296),
    .D(n3295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3299));
 sky130_fd_sc_hd__a22o_1 U3845 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[0] ),
    .A2(net209),
    .B1(n3300),
    .B2(n3299),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3302));
 sky130_fd_sc_hd__a31o_1 U3846 (.A1(n3304),
    .A2(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ),
    .A3(n3303),
    .B1(n3302),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1936));
 sky130_fd_sc_hd__a22o_1 U3847 (.A1(n3306),
    .A2(net150),
    .B1(n3305),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1935));
 sky130_fd_sc_hd__a22o_1 U3848 (.A1(n3308),
    .A2(net150),
    .B1(n3307),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1934));
 sky130_fd_sc_hd__a22o_1 U3849 (.A1(n3310),
    .A2(net141),
    .B1(n3309),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1933));
 sky130_fd_sc_hd__a22o_1 U3850 (.A1(n3312),
    .A2(net150),
    .B1(n3311),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1932));
 sky130_fd_sc_hd__a22o_1 U3851 (.A1(n3314),
    .A2(net150),
    .B1(n3313),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1931));
 sky130_fd_sc_hd__a22o_1 U3852 (.A1(n3316),
    .A2(net150),
    .B1(n3315),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1930));
 sky130_fd_sc_hd__a22o_1 U3853 (.A1(n3318),
    .A2(net150),
    .B1(n3317),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1929));
 sky130_fd_sc_hd__a22o_1 U3854 (.A1(n3320),
    .A2(net150),
    .B1(n3319),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1928));
 sky130_fd_sc_hd__a22o_1 U3855 (.A1(n3322),
    .A2(net141),
    .B1(n3321),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1927));
 sky130_fd_sc_hd__a22o_1 U3856 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ),
    .A2(n3337),
    .B1(n3323),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3324));
 sky130_fd_sc_hd__a221o_1 U3857 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .A2(n3326),
    .B1(n3325),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ),
    .C1(n3324),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3327));
 sky130_fd_sc_hd__a221o_1 U3858 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ),
    .A2(n3333),
    .B1(n3328),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[3] ),
    .C1(n3327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3329));
 sky130_fd_sc_hd__a221o_1 U3859 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ),
    .A2(n3331),
    .B1(n3330),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ),
    .C1(n3329),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3343));
 sky130_fd_sc_hd__or2_1 U3860 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3340));
 sky130_fd_sc_hd__nand2_1 U3861 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3339));
 sky130_fd_sc_hd__inv_1 U3862 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3334));
 sky130_fd_sc_hd__a221o_1 U3863 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[3] ),
    .A2(n3334),
    .B1(n3333),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ),
    .C1(n3332),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3335));
 sky130_fd_sc_hd__a221o_1 U3864 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[2] ),
    .A2(n3337),
    .B1(n3336),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ),
    .C1(n3335),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3338));
 sky130_fd_sc_hd__a32o_1 U3865 (.A1(n3341),
    .A2(n3340),
    .A3(n3339),
    .B1(n3341),
    .B2(n3338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3342));
 sky130_fd_sc_hd__a31o_1 U3866 (.A1(inst_to_wrap_u_usb_cdc_bulk_in_valid),
    .A2(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q),
    .A3(n3343),
    .B1(n3342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1926));
 sky130_fd_sc_hd__nor2_1 U3867 (.A(n3345),
    .B(n3344),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3346));
 sky130_fd_sc_hd__o31a_1 U3868 (.A1(n3499),
    .A2(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q),
    .A3(n3346),
    .B1(n3467),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3347));
 sky130_fd_sc_hd__a31o_1 U3869 (.A1(n3349),
    .A2(n3351),
    .A3(n3348),
    .B1(n3347),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3354));
 sky130_fd_sc_hd__nand2_1 U3870 (.A(n3351),
    .B(n3350),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3352));
 sky130_fd_sc_hd__nand2_1 U3871 (.A(n3355),
    .B(n3352),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3353));
 sky130_fd_sc_hd__a22o_1 U3872 (.A1(n3355),
    .A2(n3354),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ),
    .B2(n3353),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1925));
 sky130_fd_sc_hd__or2_2 U3873 (.A(n3356),
    .B(n3442),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3375));
 sky130_fd_sc_hd__inv_2 U3874 (.A(n3375),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3376));
 sky130_fd_sc_hd__a22o_1 U3875 (.A1(n3376),
    .A2(net214),
    .B1(n3375),
    .B2(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1924));
 sky130_fd_sc_hd__clkinv_2 U3876 (.A(n3365),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3370));
 sky130_fd_sc_hd__nand2_1 U3877 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ),
    .B(n3357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3358));
 sky130_fd_sc_hd__mux2_1 U3878 (.A0(n3359),
    .A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ),
    .S(n3358),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3360));
 sky130_fd_sc_hd__a22o_1 U3879 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ),
    .A2(n3367),
    .B1(n3370),
    .B2(n3360),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1923));
 sky130_fd_sc_hd__a22o_1 U3880 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[0] ),
    .A2(n3367),
    .B1(n3361),
    .B2(n3370),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1922));
 sky130_fd_sc_hd__a22o_1 U3881 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ),
    .A2(n3367),
    .B1(n3370),
    .B2(n3362),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1921));
 sky130_fd_sc_hd__a21o_1 U3882 (.A1(n3370),
    .A2(n3363),
    .B1(n3367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3364));
 sky130_fd_sc_hd__a22o_1 U3883 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .A2(n3364),
    .B1(n3418),
    .B2(n3370),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1920));
 sky130_fd_sc_hd__a21o_1 U3884 (.A1(n3370),
    .A2(n3369),
    .B1(n3367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3366));
 sky130_fd_sc_hd__nor2_1 U3885 (.A(n3369),
    .B(n3365),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3371));
 sky130_fd_sc_hd__a22o_1 U3886 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ),
    .A2(n3366),
    .B1(n3368),
    .B2(n3371),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1919));
 sky130_fd_sc_hd__a221o_1 U3887 (.A1(n3370),
    .A2(n3369),
    .B1(n3370),
    .B2(n3368),
    .C1(n3367),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3373));
 sky130_fd_sc_hd__a22o_1 U3888 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ),
    .A2(n3373),
    .B1(n3372),
    .B2(n3371),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1918));
 sky130_fd_sc_hd__nor2_1 U3889 (.A(n3442),
    .B(n3395),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3374));
 sky130_fd_sc_hd__mux2_1 U3890 (.A0(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_endp_q),
    .A1(net214),
    .S(n3374),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1916));
 sky130_fd_sc_hd__a22o_1 U3891 (.A1(n3376),
    .A2(net216),
    .B1(n3375),
    .B2(inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1915));
 sky130_fd_sc_hd__a22o_1 U3892 (.A1(n3376),
    .A2(net210),
    .B1(n3375),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1914));
 sky130_fd_sc_hd__a22o_1 U3893 (.A1(n3376),
    .A2(net212),
    .B1(n3375),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1913));
 sky130_fd_sc_hd__inv_2 U3894 (.A(inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3412));
 sky130_fd_sc_hd__or4_1 U3895 (.A(net219),
    .B(n3379),
    .C(n3378),
    .D(n3377),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3382));
 sky130_fd_sc_hd__inv_1 U3896 (.A(n3426),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3381));
 sky130_fd_sc_hd__a211o_1 U3897 (.A1(n3382),
    .A2(n3393),
    .B1(n3381),
    .C1(n3380),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3383));
 sky130_fd_sc_hd__and4b_1 U3898 (.A_N(n3383),
    .B(n3384),
    .C(n3428),
    .D(n3412),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3385));
 sky130_fd_sc_hd__a31o_1 U3899 (.A1(n3418),
    .A2(n3387),
    .A3(n3386),
    .B1(n3385),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3401));
 sky130_fd_sc_hd__o22a_1 U3900 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .A2(n3417),
    .B1(n2283),
    .B2(n3388),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3398));
 sky130_fd_sc_hd__o21ai_1 U3901 (.A1(n3391),
    .A2(n3390),
    .B1(n3389),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3392));
 sky130_fd_sc_hd__o31a_1 U3902 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .A2(n3394),
    .A3(n3393),
    .B1(n3392),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3396));
 sky130_fd_sc_hd__o22a_1 U3903 (.A1(n3398),
    .A2(n3397),
    .B1(n3396),
    .B2(n3395),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3399));
 sky130_fd_sc_hd__nand2_1 U3904 (.A(n3438),
    .B(n3399),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3400));
 sky130_fd_sc_hd__a22o_1 U3905 (.A1(n3438),
    .A2(n3401),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[2] ),
    .B2(n3400),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1912));
 sky130_fd_sc_hd__nand2_1 U3906 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3403));
 sky130_fd_sc_hd__or4_1 U3907 (.A(net214),
    .B(n3404),
    .C(n3403),
    .D(n3402),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3413));
 sky130_fd_sc_hd__o31a_1 U3908 (.A1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .A2(n3405),
    .A3(n3425),
    .B1(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3408));
 sky130_fd_sc_hd__or4_1 U3909 (.A(n3409),
    .B(n3408),
    .C(n3407),
    .D(n3406),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3411));
 sky130_fd_sc_hd__a221o_1 U3910 (.A1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q),
    .A2(n3413),
    .B1(n3412),
    .B2(n3411),
    .C1(n3410),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3421));
 sky130_fd_sc_hd__inv_1 U3911 (.A(n3414),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3420));
 sky130_fd_sc_hd__a211o_1 U3912 (.A1(n3418),
    .A2(n3417),
    .B1(n3416),
    .C1(n3415),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3419));
 sky130_fd_sc_hd__a211o_1 U3913 (.A1(n3426),
    .A2(n3421),
    .B1(n3420),
    .C1(n3419),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3423));
 sky130_fd_sc_hd__or2_1 U3914 (.A(n3435),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3422));
 sky130_fd_sc_hd__a22o_1 U3915 (.A1(n3438),
    .A2(n3423),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B2(n3422),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1911));
 sky130_fd_sc_hd__o21a_1 U3916 (.A1(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q),
    .A2(n3425),
    .B1(n3424),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3429));
 sky130_fd_sc_hd__o31a_1 U3917 (.A1(n3429),
    .A2(n3428),
    .A3(n3427),
    .B1(n3426),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3431));
 sky130_fd_sc_hd__or4_1 U3918 (.A(n3433),
    .B(n3432),
    .C(n3431),
    .D(n3430),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3437));
 sky130_fd_sc_hd__or2_1 U3919 (.A(n3435),
    .B(n3434),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3436));
 sky130_fd_sc_hd__a22o_1 U3920 (.A1(n3438),
    .A2(n3437),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[1] ),
    .B2(n3436),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1910));
 sky130_fd_sc_hd__or4_1 U3921 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[0] ),
    .C(n3440),
    .D(n3439),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3441));
 sky130_fd_sc_hd__or2_1 U3922 (.A(n3442),
    .B(n3441),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3448));
 sky130_fd_sc_hd__nor2_1 U3923 (.A(n3443),
    .B(n3448),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3447));
 sky130_fd_sc_hd__nand2_1 U3924 (.A(n3447),
    .B(n3446),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3444));
 sky130_fd_sc_hd__a22o_1 U3925 (.A1(n3447),
    .A2(n3445),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[0] ),
    .B2(n3444),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1909));
 sky130_fd_sc_hd__a21o_1 U3926 (.A1(n3447),
    .A2(n3446),
    .B1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1908));
 sky130_fd_sc_hd__or3_4 U3927 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(n3448),
    .C(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3449));
 sky130_fd_sc_hd__inv_2 U3928 (.A(n3449),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3450));
 sky130_fd_sc_hd__a22o_1 U3929 (.A1(n3450),
    .A2(\inst_to_wrap_u_usb_cdc_out_data[2] ),
    .B1(n3449),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1907));
 sky130_fd_sc_hd__a22o_1 U3930 (.A1(n3450),
    .A2(net210),
    .B1(n3449),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1906));
 sky130_fd_sc_hd__a22o_1 U3931 (.A1(n3450),
    .A2(net212),
    .B1(n3449),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1905));
 sky130_fd_sc_hd__a22o_1 U3932 (.A1(n3450),
    .A2(\inst_to_wrap_u_usb_cdc_out_data[6] ),
    .B1(n3449),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1904));
 sky130_fd_sc_hd__a22o_1 U3933 (.A1(n3450),
    .A2(\inst_to_wrap_u_usb_cdc_out_data[5] ),
    .B1(n3449),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1903));
 sky130_fd_sc_hd__a22o_1 U3934 (.A1(n3450),
    .A2(\inst_to_wrap_u_usb_cdc_out_data[4] ),
    .B1(n3449),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1902));
 sky130_fd_sc_hd__a22o_1 U3935 (.A1(n3450),
    .A2(\inst_to_wrap_u_usb_cdc_out_data[3] ),
    .B1(n3449),
    .B2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1901));
 sky130_fd_sc_hd__o22a_1 U3936 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[4] ),
    .A2(n3452),
    .B1(net217),
    .B2(n3451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1900));
 sky130_fd_sc_hd__o22a_1 U3937 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[5] ),
    .A2(n3452),
    .B1(net216),
    .B2(n3451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1899));
 sky130_fd_sc_hd__o22a_1 U3938 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[6] ),
    .A2(n3452),
    .B1(net215),
    .B2(n3451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1898));
 sky130_fd_sc_hd__o22a_1 U3939 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[2] ),
    .A2(n3452),
    .B1(net219),
    .B2(n3451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1897));
 sky130_fd_sc_hd__o22a_1 U3940 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[1] ),
    .A2(n3452),
    .B1(net210),
    .B2(n3451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1896));
 sky130_fd_sc_hd__o22a_1 U3941 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[0] ),
    .A2(n3452),
    .B1(net212),
    .B2(n3451),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1895));
 sky130_fd_sc_hd__a21oi_1 U3942 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[0] ),
    .A2(n3454),
    .B1(n3453),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1894));
 sky130_fd_sc_hd__or2_1 U3943 (.A(n3457),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3455));
 sky130_fd_sc_hd__a31o_1 U3944 (.A1(n3456),
    .A2(n3462),
    .A3(n3455),
    .B1(n3460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1893));
 sky130_fd_sc_hd__inv_1 U3945 (.A(n3457),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3459));
 sky130_fd_sc_hd__nand2_1 U3946 (.A(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3463));
 sky130_fd_sc_hd__nand2b_1 U3947 (.A_N(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[2] ),
    .B(n3463),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3458));
 sky130_fd_sc_hd__a31o_1 U3948 (.A1(n3459),
    .A2(n3462),
    .A3(n3458),
    .B1(n3460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1892));
 sky130_fd_sc_hd__or2_1 U3949 (.A(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[0] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3461));
 sky130_fd_sc_hd__a31o_1 U3950 (.A1(n3463),
    .A2(n3462),
    .A3(n3461),
    .B1(n3460),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1891));
 sky130_fd_sc_hd__nor2_2 U3951 (.A(n3470),
    .B(n3468),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3472));
 sky130_fd_sc_hd__or3_2 U3952 (.A(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ),
    .B(n3470),
    .C(n3469),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3471));
 sky130_fd_sc_hd__a22o_1 U3953 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[0] ),
    .A2(n3472),
    .B1(\inst_to_wrap_u_usb_cdc_addr[0] ),
    .B2(n3471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1890));
 sky130_fd_sc_hd__a22o_1 U3954 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[1] ),
    .A2(n3472),
    .B1(\inst_to_wrap_u_usb_cdc_addr[1] ),
    .B2(n3471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1889));
 sky130_fd_sc_hd__a22o_1 U3955 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[2] ),
    .A2(n3472),
    .B1(\inst_to_wrap_u_usb_cdc_addr[2] ),
    .B2(n3471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1888));
 sky130_fd_sc_hd__a22o_1 U3956 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[3] ),
    .A2(n3472),
    .B1(\inst_to_wrap_u_usb_cdc_addr[3] ),
    .B2(n3471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1887));
 sky130_fd_sc_hd__a22o_1 U3957 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[4] ),
    .A2(n3472),
    .B1(\inst_to_wrap_u_usb_cdc_addr[4] ),
    .B2(n3471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1886));
 sky130_fd_sc_hd__a22o_1 U3958 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[5] ),
    .A2(n3472),
    .B1(\inst_to_wrap_u_usb_cdc_addr[5] ),
    .B2(n3471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1885));
 sky130_fd_sc_hd__a22o_1 U3959 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[6] ),
    .A2(n3472),
    .B1(\inst_to_wrap_u_usb_cdc_addr[6] ),
    .B2(n3471),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1884));
 sky130_fd_sc_hd__inv_2 U3960 (.A(n3569),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3496));
 sky130_fd_sc_hd__inv_1 U3961 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3473));
 sky130_fd_sc_hd__a21oi_1 U3962 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[1] ),
    .A2(n3473),
    .B1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_full_o),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3474));
 sky130_fd_sc_hd__and3_1 U3963 (.A(n3475),
    .B(n3499),
    .C(n3474),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3568));
 sky130_fd_sc_hd__a22o_1 U3964 (.A1(n3496),
    .A2(n3568),
    .B1(n3569),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1883));
 sky130_fd_sc_hd__or3_1 U3965 (.A(inst_to_wrap_u_usb_cdc_out_err),
    .B(n3474),
    .C(n3477),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3498));
 sky130_fd_sc_hd__nand2_1 U3966 (.A(n3496),
    .B(n3498),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3476));
 sky130_fd_sc_hd__o21a_1 U3967 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[1] ),
    .A2(n3496),
    .B1(n3476),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1882));
 sky130_fd_sc_hd__a31o_1 U3968 (.A1(n3477),
    .A2(n3475),
    .A3(n3495),
    .B1(n3476),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3483));
 sky130_fd_sc_hd__inv_2 U3969 (.A(n3476),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3478));
 sky130_fd_sc_hd__a32o_1 U3970 (.A1(n3478),
    .A2(inst_to_wrap_u_usb_cdc_bulk_out_nak),
    .A3(n3477),
    .B1(n3478),
    .B2(inst_to_wrap_u_usb_cdc_out_err),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3488));
 sky130_fd_sc_hd__inv_2 U3971 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3810));
 sky130_fd_sc_hd__or3_1 U3972 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3577));
 sky130_fd_sc_hd__nor2_1 U3973 (.A(n3810),
    .B(n3577),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3492));
 sky130_fd_sc_hd__nor2b_1 U3974 (.A(n3492),
    .B_N(n3568),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3487));
 sky130_fd_sc_hd__and2_1 U3975 (.A(n3487),
    .B(n3478),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3480));
 sky130_fd_sc_hd__inv_2 U3976 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3813));
 sky130_fd_sc_hd__a22o_1 U3977 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[0] ),
    .A2(n3488),
    .B1(n3480),
    .B2(n3813),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3479));
 sky130_fd_sc_hd__a21o_1 U3978 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .A2(n3483),
    .B1(n3479),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1881));
 sky130_fd_sc_hd__nand2_1 U3979 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .B(n3480),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3484));
 sky130_fd_sc_hd__nor2_1 U3980 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .B(n3484),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3482));
 sky130_fd_sc_hd__a32o_1 U3981 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .A2(n3487),
    .A3(n3813),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .B2(n3483),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3481));
 sky130_fd_sc_hd__a211o_1 U3982 (.A1(n3488),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[1] ),
    .B1(n3482),
    .C1(n3481),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1880));
 sky130_fd_sc_hd__clkinv_2 U3983 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3804));
 sky130_fd_sc_hd__a221o_1 U3984 (.A1(n3487),
    .A2(n3813),
    .B1(n3487),
    .B2(n3804),
    .C1(n3483),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3486));
 sky130_fd_sc_hd__nor2_1 U3985 (.A(n3804),
    .B(n3484),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3491));
 sky130_fd_sc_hd__inv_2 U3986 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3806));
 sky130_fd_sc_hd__a22o_1 U3987 (.A1(n3488),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[2] ),
    .B1(n3491),
    .B2(n3806),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3485));
 sky130_fd_sc_hd__a21o_1 U3988 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ),
    .A2(n3486),
    .B1(n3485),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1879));
 sky130_fd_sc_hd__a21o_1 U3989 (.A1(n3487),
    .A2(n3806),
    .B1(n3486),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3489));
 sky130_fd_sc_hd__a22o_1 U3990 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[3] ),
    .A2(n3489),
    .B1(n3488),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3490));
 sky130_fd_sc_hd__a31o_1 U3991 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ),
    .A2(n3491),
    .A3(n3810),
    .B1(n3490),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1878));
 sky130_fd_sc_hd__and3_2 U3992 (.A(n3568),
    .B(n3492),
    .C(n3496),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3494));
 sky130_fd_sc_hd__clkinv_2 U3993 (.A(n3494),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3493));
 sky130_fd_sc_hd__a22o_1 U3994 (.A1(n3494),
    .A2(net214),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1877));
 sky130_fd_sc_hd__a22o_1 U3995 (.A1(n3494),
    .A2(net215),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1876));
 sky130_fd_sc_hd__a22o_1 U3996 (.A1(n3494),
    .A2(net216),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1875));
 sky130_fd_sc_hd__a22o_1 U3997 (.A1(n3494),
    .A2(net217),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1874));
 sky130_fd_sc_hd__a22o_1 U3998 (.A1(n3494),
    .A2(net218),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1873));
 sky130_fd_sc_hd__a22o_1 U3999 (.A1(n3494),
    .A2(net219),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1872));
 sky130_fd_sc_hd__a22o_1 U4000 (.A1(n3494),
    .A2(net210),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1871));
 sky130_fd_sc_hd__a22o_1 U4001 (.A1(n3494),
    .A2(net212),
    .B1(n3493),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1870));
 sky130_fd_sc_hd__a221o_1 U4002 (.A1(n3496),
    .A2(n3499),
    .B1(n3496),
    .B2(inst_to_wrap_u_usb_cdc_out_err),
    .C1(n3495),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3497));
 sky130_fd_sc_hd__o21ai_1 U4003 (.A1(n3498),
    .A2(n3569),
    .B1(n3497),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1869));
 sky130_fd_sc_hd__or4_2 U4004 (.A(n3499),
    .B(inst_to_wrap_u_usb_cdc_out_err),
    .C(inst_to_wrap_u_usb_cdc_bulk_out_nak),
    .D(n3569),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3500));
 sky130_fd_sc_hd__inv_2 U4005 (.A(n3500),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3501));
 sky130_fd_sc_hd__mux2_1 U4006 (.A0(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[0] ),
    .A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .S(n3501),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1868));
 sky130_fd_sc_hd__a22o_1 U4007 (.A1(n3501),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .B1(n3500),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1867));
 sky130_fd_sc_hd__a22o_1 U4008 (.A1(n3501),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ),
    .B1(n3500),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1866));
 sky130_fd_sc_hd__a22o_1 U4009 (.A1(n3501),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[3] ),
    .B1(n3500),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1865));
 sky130_fd_sc_hd__inv_2 U4010 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3797));
 sky130_fd_sc_hd__nor2_1 U4011 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3798));
 sky130_fd_sc_hd__inv_2 U4012 (.A(n3798),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3796));
 sky130_fd_sc_hd__inv_2 U4013 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3505));
 sky130_fd_sc_hd__or3_2 U4014 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .C(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3795));
 sky130_fd_sc_hd__or2_2 U4015 (.A(n3505),
    .B(n3795),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3596));
 sky130_fd_sc_hd__inv_2 U4016 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3799));
 sky130_fd_sc_hd__clkinv_2 U4017 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3592));
 sky130_fd_sc_hd__inv_1 U4018 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3507));
 sky130_fd_sc_hd__inv_1 U4019 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3504));
 sky130_fd_sc_hd__o22ai_1 U4020 (.A1(n3592),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[0] ),
    .B1(n3799),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3502));
 sky130_fd_sc_hd__a221o_1 U4021 (.A1(n3592),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[0] ),
    .B1(n3799),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[1] ),
    .C1(n3502),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3503));
 sky130_fd_sc_hd__a221o_1 U4022 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[3] ),
    .A2(n3505),
    .B1(n3504),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .C1(n3503),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3506));
 sky130_fd_sc_hd__a221o_1 U4023 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[2] ),
    .A2(n3797),
    .B1(n3507),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ),
    .C1(n3506),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3508));
 sky130_fd_sc_hd__and3_4 U4024 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[0] ),
    .C(n3567),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3666));
 sky130_fd_sc_hd__inv_2 U4025 (.A(n3666),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3664));
 sky130_fd_sc_hd__a221o_1 U4026 (.A1(n3596),
    .A2(n3799),
    .B1(n3596),
    .B2(n3592),
    .C1(n3664),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3511));
 sky130_fd_sc_hd__or2_1 U4027 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .B(n3797),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3595));
 sky130_fd_sc_hd__inv_2 U4028 (.A(n3595),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3591));
 sky130_fd_sc_hd__and3_2 U4029 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .C(n3591),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3655));
 sky130_fd_sc_hd__a22o_1 U4030 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .A2(n3511),
    .B1(n3666),
    .B2(n3655),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3509));
 sky130_fd_sc_hd__a31o_1 U4031 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .A2(n3797),
    .A3(n3796),
    .B1(n3509),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1864));
 sky130_fd_sc_hd__a21o_1 U4032 (.A1(n3592),
    .A2(n3596),
    .B1(n3664),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3510));
 sky130_fd_sc_hd__o21a_1 U4033 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .A2(n3666),
    .B1(n3510),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1863));
 sky130_fd_sc_hd__nor2_1 U4034 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .B(n3592),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3593));
 sky130_fd_sc_hd__a22o_1 U4035 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .A2(n3510),
    .B1(n3666),
    .B2(n3593),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1862));
 sky130_fd_sc_hd__nor2_1 U4036 (.A(n3799),
    .B(n3592),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3512));
 sky130_fd_sc_hd__a32o_1 U4037 (.A1(n3666),
    .A2(n3797),
    .A3(n3512),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ),
    .B2(n3511),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1861));
 sky130_fd_sc_hd__nand2_1 U4038 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3814));
 sky130_fd_sc_hd__a221o_1 U4039 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_mask_q),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq[0] ),
    .B1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_mask_q),
    .B2(n3814),
    .C1(n3666),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1860));
 sky130_fd_sc_hd__o21a_1 U4040 (.A1(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_mask_q),
    .A2(n3513),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1859));
 sky130_fd_sc_hd__nand2_2 U4041 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[0] ),
    .B(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3610));
 sky130_fd_sc_hd__a22o_1 U4042 (.A1(n3524),
    .A2(n3546),
    .B1(n3609),
    .B2(\inst_to_wrap_rx_fifo_w_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1858));
 sky130_fd_sc_hd__inv_2 U4043 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3603));
 sky130_fd_sc_hd__a22o_1 U4044 (.A1(n3524),
    .A2(n3603),
    .B1(n3609),
    .B2(\inst_to_wrap_rx_fifo_w_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1857));
 sky130_fd_sc_hd__or2_2 U4045 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[0] ),
    .B(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3614));
 sky130_fd_sc_hd__a32o_1 U4046 (.A1(n3524),
    .A2(n3610),
    .A3(n3614),
    .B1(n3609),
    .B2(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1856));
 sky130_fd_sc_hd__inv_2 U4047 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3605));
 sky130_fd_sc_hd__inv_2 U4048 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3607));
 sky130_fd_sc_hd__nor2_1 U4049 (.A(n3607),
    .B(n3610),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3514));
 sky130_fd_sc_hd__mux2_1 U4050 (.A0(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ),
    .A1(n3605),
    .S(n3514),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3548));
 sky130_fd_sc_hd__a22o_1 U4051 (.A1(n3524),
    .A2(n3548),
    .B1(n3609),
    .B2(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1855));
 sky130_fd_sc_hd__nor2_1 U4052 (.A(n3524),
    .B(n3520),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3527));
 sky130_fd_sc_hd__a22o_1 U4053 (.A1(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .A2(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .B1(n3560),
    .B2(n3559),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3561));
 sky130_fd_sc_hd__nand2_1 U4054 (.A(n3561),
    .B(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3519));
 sky130_fd_sc_hd__nor2_1 U4055 (.A(n3560),
    .B(n3559),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3515));
 sky130_fd_sc_hd__mux2_1 U4056 (.A0(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .A1(n3547),
    .S(n3515),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3564));
 sky130_fd_sc_hd__a22oi_1 U4057 (.A1(n3607),
    .A2(n3564),
    .B1(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ),
    .B2(n3517),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3516));
 sky130_fd_sc_hd__o221a_1 U4058 (.A1(n3607),
    .A2(n3564),
    .B1(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ),
    .B2(n3517),
    .C1(n3516),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3518));
 sky130_fd_sc_hd__a22o_1 U4059 (.A1(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .A2(n3603),
    .B1(n3559),
    .B2(\inst_to_wrap_rx_fifo_w_ptr_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3551));
 sky130_fd_sc_hd__o2111a_1 U4060 (.A1(n3561),
    .A2(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ),
    .B1(n3519),
    .C1(n3518),
    .D1(n3551),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3521));
 sky130_fd_sc_hd__inv_2 U4061 (.A(n3520),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3523));
 sky130_fd_sc_hd__o21ai_2 U4062 (.A1(n3524),
    .A2(n_RX_EMPTY_FLAG_FLAG_),
    .B1(n3523),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3530));
 sky130_fd_sc_hd__o21ai_1 U4063 (.A1(n3524),
    .A2(n3523),
    .B1(n3530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3556));
 sky130_fd_sc_hd__a22o_1 U4064 (.A1(n3527),
    .A2(n3521),
    .B1(n_RX_EMPTY_FLAG_FLAG_),
    .B2(n3556),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1854));
 sky130_fd_sc_hd__inv_2 U4065 (.A(\RXFIFOLEVEL_REG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3535));
 sky130_fd_sc_hd__nor2_1 U4066 (.A(n3523),
    .B(n3609),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3555));
 sky130_fd_sc_hd__or2_1 U4067 (.A(n3527),
    .B(n3555),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3522));
 sky130_fd_sc_hd__a32o_1 U4068 (.A1(n3535),
    .A2(n3530),
    .A3(n3522),
    .B1(\RXFIFOLEVEL_REG[0] ),
    .B2(n3556),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1853));
 sky130_fd_sc_hd__o221ai_2 U4069 (.A1(n3535),
    .A2(n3524),
    .B1(\RXFIFOLEVEL_REG[0] ),
    .B2(n3523),
    .C1(n3530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3526));
 sky130_fd_sc_hd__inv_2 U4070 (.A(\RXFIFOLEVEL_REG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3536));
 sky130_fd_sc_hd__o221a_1 U4071 (.A1(\RXFIFOLEVEL_REG[0] ),
    .A2(n3527),
    .B1(n3535),
    .B2(n3555),
    .C1(n3530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3525));
 sky130_fd_sc_hd__a22o_1 U4072 (.A1(\RXFIFOLEVEL_REG[1] ),
    .A2(n3526),
    .B1(n3536),
    .B2(n3525),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1852));
 sky130_fd_sc_hd__inv_2 U4073 (.A(\RXFIFOLEVEL_REG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3537));
 sky130_fd_sc_hd__and3_1 U4074 (.A(n3555),
    .B(\RXFIFOLEVEL_REG[1] ),
    .C(\RXFIFOLEVEL_REG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3531));
 sky130_fd_sc_hd__and3_1 U4075 (.A(n3527),
    .B(n3536),
    .C(n3535),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3532));
 sky130_fd_sc_hd__or2_1 U4076 (.A(n3531),
    .B(n3532),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3529));
 sky130_fd_sc_hd__a221o_1 U4077 (.A1(\RXFIFOLEVEL_REG[1] ),
    .A2(n3527),
    .B1(n3536),
    .B2(n3555),
    .C1(n3526),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3528));
 sky130_fd_sc_hd__a32o_1 U4078 (.A1(n3537),
    .A2(n3530),
    .A3(n3529),
    .B1(\RXFIFOLEVEL_REG[2] ),
    .B2(n3528),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1851));
 sky130_fd_sc_hd__o221a_1 U4079 (.A1(\RXFIFOLEVEL_REG[2] ),
    .A2(n3532),
    .B1(n3537),
    .B2(n3531),
    .C1(n3530),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3533));
 sky130_fd_sc_hd__inv_2 U4081 (.A(\RXFIFOLEVEL_REG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3541));
 sky130_fd_sc_hd__inv_1 U4083 (.A(\RIS_REG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3544));
 sky130_fd_sc_hd__o22a_1 U4084 (.A1(\rx_fifo_th[1] ),
    .A2(n3536),
    .B1(\rx_fifo_th[2] ),
    .B2(n3537),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3539));
 sky130_fd_sc_hd__a211o_1 U4085 (.A1(\rx_fifo_th[1] ),
    .A2(n3536),
    .B1(\rx_fifo_th[0] ),
    .C1(n3535),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3538));
 sky130_fd_sc_hd__a22o_1 U4086 (.A1(n3539),
    .A2(n3538),
    .B1(\rx_fifo_th[2] ),
    .B2(n3537),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3542));
 sky130_fd_sc_hd__or2_1 U4087 (.A(n3542),
    .B(n3541),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3540));
 sky130_fd_sc_hd__a22o_1 U4088 (.A1(n3542),
    .A2(n3541),
    .B1(\rx_fifo_th[3] ),
    .B2(n3540),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3543));
 sky130_fd_sc_hd__o21ai_1 U4089 (.A1(\ICR_REG[3] ),
    .A2(n3544),
    .B1(n3543),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1849));
 sky130_fd_sc_hd__nand2_1 U4090 (.A(n3610),
    .B(n3614),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3553));
 sky130_fd_sc_hd__a22oi_1 U4091 (.A1(n3549),
    .A2(n3548),
    .B1(n3547),
    .B2(n3546),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3545));
 sky130_fd_sc_hd__o221a_1 U4092 (.A1(n3549),
    .A2(n3548),
    .B1(n3547),
    .B2(n3546),
    .C1(n3545),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3552));
 sky130_fd_sc_hd__nand2_1 U4093 (.A(n3553),
    .B(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3550));
 sky130_fd_sc_hd__o2111a_1 U4094 (.A1(n3553),
    .A2(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ),
    .B1(n3552),
    .C1(n3551),
    .D1(n3550),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3554));
 sky130_fd_sc_hd__a22o_1 U4095 (.A1(n_RX_FULL_FLAG_FLAG_),
    .A2(n3556),
    .B1(n3555),
    .B2(n3554),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1848));
 sky130_fd_sc_hd__inv_1 U4096 (.A(\ICR_REG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3557));
 sky130_fd_sc_hd__a21o_1 U4097 (.A1(n3557),
    .A2(\RIS_REG[2] ),
    .B1(n_RX_FULL_FLAG_FLAG_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1847));
 sky130_fd_sc_hd__inv_1 U4098 (.A(\ICR_REG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3558));
 sky130_fd_sc_hd__a21o_1 U4099 (.A1(\RIS_REG[4] ),
    .A2(n3558),
    .B1(n_RX_EMPTY_FLAG_FLAG_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1846));
 sky130_fd_sc_hd__inv_2 U4100 (.A(n3563),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3565));
 sky130_fd_sc_hd__a22o_1 U4101 (.A1(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ),
    .A2(n3563),
    .B1(n3559),
    .B2(n3565),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1845));
 sky130_fd_sc_hd__mux2_1 U4102 (.A0(n3561),
    .A1(n3560),
    .S(n3563),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3562));
 sky130_fd_sc_hd__inv_1 U4103 (.A(n3562),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1844));
 sky130_fd_sc_hd__a22o_1 U4104 (.A1(n3565),
    .A2(n3564),
    .B1(n3563),
    .B2(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1843));
 sky130_fd_sc_hd__inv_1 U4105 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3566));
 sky130_fd_sc_hd__o21ai_1 U4106 (.A1(n3567),
    .A2(n3566),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n1841));
 sky130_fd_sc_hd__a22o_1 U4107 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[1] ),
    .A2(n3664),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[0] ),
    .B2(n3814),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1840));
 sky130_fd_sc_hd__or3b_2 U4108 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[3] ),
    .B(n3569),
    .C_N(n3568),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3582));
 sky130_fd_sc_hd__or3_1 U4109 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ),
    .B(n3813),
    .C(n3582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3574));
 sky130_fd_sc_hd__or2_4 U4110 (.A(n3804),
    .B(n3574),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3570));
 sky130_fd_sc_hd__clkinv_2 U4111 (.A(n3570),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3571));
 sky130_fd_sc_hd__a22o_1 U4112 (.A1(n3571),
    .A2(net214),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1839));
 sky130_fd_sc_hd__a22o_1 U4113 (.A1(n3571),
    .A2(net215),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1838));
 sky130_fd_sc_hd__a22o_1 U4114 (.A1(n3571),
    .A2(net216),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1837));
 sky130_fd_sc_hd__a22o_1 U4115 (.A1(n3571),
    .A2(net217),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1836));
 sky130_fd_sc_hd__a22o_1 U4116 (.A1(n3571),
    .A2(net218),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1835));
 sky130_fd_sc_hd__a22o_1 U4117 (.A1(n3571),
    .A2(net219),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1834));
 sky130_fd_sc_hd__a22o_1 U4118 (.A1(n3571),
    .A2(net210),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1833));
 sky130_fd_sc_hd__a22o_1 U4119 (.A1(n3571),
    .A2(net212),
    .B1(n3570),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1832));
 sky130_fd_sc_hd__or4_4 U4120 (.A(n3804),
    .B(n3582),
    .C(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ),
    .D(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3572));
 sky130_fd_sc_hd__clkinv_2 U4121 (.A(n3572),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3573));
 sky130_fd_sc_hd__a22o_1 U4122 (.A1(n3573),
    .A2(net214),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1831));
 sky130_fd_sc_hd__a22o_1 U4123 (.A1(n3573),
    .A2(net215),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1830));
 sky130_fd_sc_hd__a22o_1 U4124 (.A1(n3573),
    .A2(net216),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1829));
 sky130_fd_sc_hd__a22o_1 U4125 (.A1(n3573),
    .A2(net217),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1828));
 sky130_fd_sc_hd__a22o_1 U4126 (.A1(n3573),
    .A2(net218),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1827));
 sky130_fd_sc_hd__a22o_1 U4127 (.A1(n3573),
    .A2(net219),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1826));
 sky130_fd_sc_hd__a22o_1 U4128 (.A1(n3573),
    .A2(net210),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1825));
 sky130_fd_sc_hd__a22o_1 U4129 (.A1(n3573),
    .A2(net212),
    .B1(n3572),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1824));
 sky130_fd_sc_hd__or2_4 U4130 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .B(n3574),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3575));
 sky130_fd_sc_hd__clkinv_2 U4131 (.A(n3575),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3576));
 sky130_fd_sc_hd__a22o_1 U4132 (.A1(n3576),
    .A2(net214),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1823));
 sky130_fd_sc_hd__a22o_1 U4133 (.A1(n3576),
    .A2(net215),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1822));
 sky130_fd_sc_hd__a22o_1 U4134 (.A1(n3576),
    .A2(net216),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1821));
 sky130_fd_sc_hd__a22o_1 U4135 (.A1(n3576),
    .A2(net217),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1820));
 sky130_fd_sc_hd__a22o_1 U4136 (.A1(n3576),
    .A2(net218),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1819));
 sky130_fd_sc_hd__a22o_1 U4137 (.A1(n3576),
    .A2(net219),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1818));
 sky130_fd_sc_hd__a22o_1 U4138 (.A1(n3576),
    .A2(net210),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1817));
 sky130_fd_sc_hd__a22o_1 U4139 (.A1(n3576),
    .A2(net212),
    .B1(n3575),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1816));
 sky130_fd_sc_hd__or2_4 U4140 (.A(n3577),
    .B(n3582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3578));
 sky130_fd_sc_hd__clkinv_2 U4141 (.A(n3578),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3579));
 sky130_fd_sc_hd__a22o_1 U4142 (.A1(n3579),
    .A2(net214),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1815));
 sky130_fd_sc_hd__a22o_1 U4143 (.A1(n3579),
    .A2(net215),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1814));
 sky130_fd_sc_hd__a22o_1 U4144 (.A1(n3579),
    .A2(net216),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1813));
 sky130_fd_sc_hd__a22o_1 U4145 (.A1(n3579),
    .A2(net217),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1812));
 sky130_fd_sc_hd__a22o_1 U4146 (.A1(n3579),
    .A2(net218),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1811));
 sky130_fd_sc_hd__a22o_1 U4147 (.A1(n3579),
    .A2(net219),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1810));
 sky130_fd_sc_hd__a22o_1 U4148 (.A1(n3579),
    .A2(net210),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1809));
 sky130_fd_sc_hd__a22o_1 U4149 (.A1(n3579),
    .A2(net212),
    .B1(n3578),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1808));
 sky130_fd_sc_hd__or3_1 U4150 (.A(n3806),
    .B(n3813),
    .C(n3582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3585));
 sky130_fd_sc_hd__or2_4 U4151 (.A(n3804),
    .B(n3585),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3580));
 sky130_fd_sc_hd__clkinv_2 U4152 (.A(n3580),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3581));
 sky130_fd_sc_hd__a22o_1 U4153 (.A1(n3581),
    .A2(net214),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1807));
 sky130_fd_sc_hd__a22o_1 U4154 (.A1(n3581),
    .A2(net215),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1806));
 sky130_fd_sc_hd__a22o_1 U4155 (.A1(n3581),
    .A2(net216),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1805));
 sky130_fd_sc_hd__a22o_1 U4156 (.A1(n3581),
    .A2(net217),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1804));
 sky130_fd_sc_hd__a22o_1 U4157 (.A1(n3581),
    .A2(net218),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1803));
 sky130_fd_sc_hd__a22o_1 U4158 (.A1(n3581),
    .A2(net219),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1802));
 sky130_fd_sc_hd__a22o_1 U4159 (.A1(n3581),
    .A2(net210),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1801));
 sky130_fd_sc_hd__a22o_1 U4160 (.A1(n3581),
    .A2(net212),
    .B1(n3580),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1800));
 sky130_fd_sc_hd__or3_1 U4161 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .B(n3806),
    .C(n3582),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3588));
 sky130_fd_sc_hd__or2_4 U4162 (.A(n3804),
    .B(n3588),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3583));
 sky130_fd_sc_hd__clkinv_2 U4163 (.A(n3583),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3584));
 sky130_fd_sc_hd__a22o_1 U4164 (.A1(n3584),
    .A2(net214),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1799));
 sky130_fd_sc_hd__a22o_1 U4165 (.A1(n3584),
    .A2(net215),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1798));
 sky130_fd_sc_hd__a22o_1 U4166 (.A1(n3584),
    .A2(net216),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1797));
 sky130_fd_sc_hd__a22o_1 U4167 (.A1(n3584),
    .A2(net217),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1796));
 sky130_fd_sc_hd__a22o_1 U4168 (.A1(n3584),
    .A2(net218),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1795));
 sky130_fd_sc_hd__a22o_1 U4169 (.A1(n3584),
    .A2(net219),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1794));
 sky130_fd_sc_hd__a22o_1 U4170 (.A1(n3584),
    .A2(net210),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1793));
 sky130_fd_sc_hd__a22o_1 U4171 (.A1(n3584),
    .A2(net212),
    .B1(n3583),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1792));
 sky130_fd_sc_hd__or2_2 U4172 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .B(n3585),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3586));
 sky130_fd_sc_hd__clkinv_2 U4173 (.A(n3586),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3587));
 sky130_fd_sc_hd__a22o_1 U4174 (.A1(n3587),
    .A2(net214),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1791));
 sky130_fd_sc_hd__a22o_1 U4175 (.A1(n3587),
    .A2(net215),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1790));
 sky130_fd_sc_hd__a22o_1 U4176 (.A1(n3587),
    .A2(net216),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1789));
 sky130_fd_sc_hd__a22o_1 U4177 (.A1(n3587),
    .A2(net217),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1788));
 sky130_fd_sc_hd__a22o_1 U4178 (.A1(n3587),
    .A2(net218),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1787));
 sky130_fd_sc_hd__a22o_1 U4179 (.A1(n3587),
    .A2(net219),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1786));
 sky130_fd_sc_hd__a22o_1 U4180 (.A1(n3587),
    .A2(net210),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1785));
 sky130_fd_sc_hd__a22o_1 U4181 (.A1(n3587),
    .A2(net212),
    .B1(n3586),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1784));
 sky130_fd_sc_hd__or2_4 U4182 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ),
    .B(n3588),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3589));
 sky130_fd_sc_hd__clkinv_2 U4183 (.A(n3589),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3590));
 sky130_fd_sc_hd__a22o_1 U4184 (.A1(n3590),
    .A2(net214),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1783));
 sky130_fd_sc_hd__a22o_1 U4185 (.A1(n3590),
    .A2(\inst_to_wrap_u_usb_cdc_out_data[6] ),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1782));
 sky130_fd_sc_hd__a22o_1 U4186 (.A1(n3590),
    .A2(net216),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1781));
 sky130_fd_sc_hd__a22o_1 U4187 (.A1(n3590),
    .A2(net217),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1780));
 sky130_fd_sc_hd__a22o_1 U4188 (.A1(n3590),
    .A2(net218),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1779));
 sky130_fd_sc_hd__a22o_1 U4189 (.A1(n3590),
    .A2(\inst_to_wrap_u_usb_cdc_out_data[2] ),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1778));
 sky130_fd_sc_hd__a22o_1 U4190 (.A1(n3590),
    .A2(net210),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1777));
 sky130_fd_sc_hd__a22o_1 U4191 (.A1(n3590),
    .A2(net212),
    .B1(n3589),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1776));
 sky130_fd_sc_hd__nor2_1 U4192 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3594));
 sky130_fd_sc_hd__and3_2 U4193 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .C(n3594),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3652));
 sky130_fd_sc_hd__and3_2 U4194 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .B(n3591),
    .C(n3592),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3651));
 sky130_fd_sc_hd__a22o_1 U4195 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[24] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[48] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3601));
 sky130_fd_sc_hd__inv_2 U4196 (.A(n3593),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3800));
 sky130_fd_sc_hd__nor2_2 U4197 (.A(n3595),
    .B(n3800),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3654));
 sky130_fd_sc_hd__and3_2 U4198 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ),
    .B(n3594),
    .C(n3592),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3653));
 sky130_fd_sc_hd__a22o_1 U4199 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[40] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[16] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3600));
 sky130_fd_sc_hd__and2_2 U4200 (.A(n3594),
    .B(n3593),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3660));
 sky130_fd_sc_hd__nor2_4 U4201 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .B(n3795),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3811));
 sky130_fd_sc_hd__a22o_1 U4202 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[56] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[0] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3598));
 sky130_fd_sc_hd__nor2_2 U4203 (.A(n3595),
    .B(n3796),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3657));
 sky130_fd_sc_hd__clkinv_2 U4204 (.A(n3596),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3656));
 sky130_fd_sc_hd__a22o_1 U4205 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[32] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[64] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3597));
 sky130_fd_sc_hd__a211o_1 U4206 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[8] ),
    .A2(n3660),
    .B1(n3598),
    .C1(n3597),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3599));
 sky130_fd_sc_hd__or3_1 U4207 (.A(n3601),
    .B(n3600),
    .C(n3599),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3602));
 sky130_fd_sc_hd__mux2_1 U4208 (.A0(n3602),
    .A1(net227),
    .S(n3664),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1775));
 sky130_fd_sc_hd__or3_2 U4209 (.A(n3609),
    .B(n3607),
    .C(n3605),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3604));
 sky130_fd_sc_hd__or2_2 U4210 (.A(n3610),
    .B(n3604),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3667));
 sky130_fd_sc_hd__clkinv_2 U4211 (.A(n3667),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3668));
 sky130_fd_sc_hd__a22o_1 U4212 (.A1(n3668),
    .A2(net252),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[120] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1774));
 sky130_fd_sc_hd__nand2_1 U4213 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ),
    .B(n3603),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3611));
 sky130_fd_sc_hd__or2_4 U4214 (.A(n3604),
    .B(n3611),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3669));
 sky130_fd_sc_hd__clkinv_2 U4215 (.A(n3669),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3670));
 sky130_fd_sc_hd__a22o_1 U4216 (.A1(n3670),
    .A2(net253),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[112] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1773));
 sky130_fd_sc_hd__or2_1 U4217 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ),
    .B(n3603),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3612));
 sky130_fd_sc_hd__or2_4 U4218 (.A(n3604),
    .B(n3612),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3671));
 sky130_fd_sc_hd__clkinv_2 U4219 (.A(n3671),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3672));
 sky130_fd_sc_hd__a22o_1 U4220 (.A1(n3672),
    .A2(net253),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[104] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1772));
 sky130_fd_sc_hd__or2_2 U4221 (.A(n3614),
    .B(n3604),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3673));
 sky130_fd_sc_hd__clkinv_2 U4222 (.A(n3673),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3674));
 sky130_fd_sc_hd__a22o_1 U4223 (.A1(n3674),
    .A2(net253),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[96] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1771));
 sky130_fd_sc_hd__or3_1 U4224 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[2] ),
    .B(n3609),
    .C(n3605),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3606));
 sky130_fd_sc_hd__or2_4 U4225 (.A(n3610),
    .B(n3606),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3675));
 sky130_fd_sc_hd__clkinv_2 U4226 (.A(n3675),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3676));
 sky130_fd_sc_hd__a22o_1 U4227 (.A1(n3676),
    .A2(net253),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[88] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1770));
 sky130_fd_sc_hd__or2_2 U4228 (.A(n3611),
    .B(n3606),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3677));
 sky130_fd_sc_hd__clkinv_2 U4229 (.A(n3677),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3678));
 sky130_fd_sc_hd__a22o_1 U4230 (.A1(n3678),
    .A2(net253),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[80] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1769));
 sky130_fd_sc_hd__or2_2 U4231 (.A(n3612),
    .B(n3606),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3679));
 sky130_fd_sc_hd__clkinv_2 U4232 (.A(n3679),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3680));
 sky130_fd_sc_hd__a22o_1 U4233 (.A1(n3680),
    .A2(net253),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[72] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1768));
 sky130_fd_sc_hd__or2_4 U4234 (.A(n3614),
    .B(n3606),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3681));
 sky130_fd_sc_hd__clkinv_2 U4235 (.A(n3681),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3682));
 sky130_fd_sc_hd__a22o_1 U4236 (.A1(n3682),
    .A2(net253),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[64] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1767));
 sky130_fd_sc_hd__or3_2 U4237 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ),
    .B(n3607),
    .C(n3609),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3608));
 sky130_fd_sc_hd__or2_4 U4238 (.A(n3610),
    .B(n3608),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3683));
 sky130_fd_sc_hd__clkinv_2 U4239 (.A(n3683),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3684));
 sky130_fd_sc_hd__a22o_1 U4240 (.A1(n3684),
    .A2(net253),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[56] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1766));
 sky130_fd_sc_hd__or2_4 U4241 (.A(n3611),
    .B(n3608),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3685));
 sky130_fd_sc_hd__clkinv_2 U4242 (.A(n3685),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3686));
 sky130_fd_sc_hd__a22o_1 U4243 (.A1(n3686),
    .A2(net253),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[48] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1765));
 sky130_fd_sc_hd__or2_4 U4244 (.A(n3612),
    .B(n3608),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3687));
 sky130_fd_sc_hd__clkinv_2 U4245 (.A(n3687),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3688));
 sky130_fd_sc_hd__a22o_1 U4246 (.A1(n3688),
    .A2(net253),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[40] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1764));
 sky130_fd_sc_hd__or2_4 U4247 (.A(n3614),
    .B(n3608),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3689));
 sky130_fd_sc_hd__clkinv_2 U4248 (.A(n3689),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3690));
 sky130_fd_sc_hd__a22o_1 U4249 (.A1(n3690),
    .A2(net253),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[32] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1763));
 sky130_fd_sc_hd__or3_2 U4250 (.A(\inst_to_wrap_rx_fifo_w_ptr_reg[2] ),
    .B(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ),
    .C(n3609),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3613));
 sky130_fd_sc_hd__or2_2 U4251 (.A(n3610),
    .B(n3613),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3691));
 sky130_fd_sc_hd__clkinv_2 U4252 (.A(n3691),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3692));
 sky130_fd_sc_hd__a22o_1 U4253 (.A1(n3692),
    .A2(net253),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[24] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1762));
 sky130_fd_sc_hd__or2_4 U4254 (.A(n3611),
    .B(n3613),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3693));
 sky130_fd_sc_hd__clkinv_2 U4255 (.A(n3693),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3694));
 sky130_fd_sc_hd__a22o_1 U4256 (.A1(n3694),
    .A2(net253),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[16] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1761));
 sky130_fd_sc_hd__or2_4 U4257 (.A(n3612),
    .B(n3613),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3695));
 sky130_fd_sc_hd__clkinv_2 U4258 (.A(n3695),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3696));
 sky130_fd_sc_hd__a22o_1 U4259 (.A1(n3696),
    .A2(net253),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1760));
 sky130_fd_sc_hd__or2_4 U4260 (.A(n3614),
    .B(n3613),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3697));
 sky130_fd_sc_hd__clkinv_2 U4261 (.A(n3697),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3698));
 sky130_fd_sc_hd__a22o_1 U4262 (.A1(n3698),
    .A2(net253),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1759));
 sky130_fd_sc_hd__a22o_1 U4263 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[25] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[49] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3619));
 sky130_fd_sc_hd__a22o_1 U4264 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[41] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[17] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3618));
 sky130_fd_sc_hd__a22o_1 U4265 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[57] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[1] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3616));
 sky130_fd_sc_hd__a22o_1 U4266 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[33] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[65] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3615));
 sky130_fd_sc_hd__a211o_1 U4267 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[9] ),
    .A2(n3660),
    .B1(n3616),
    .C1(n3615),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3617));
 sky130_fd_sc_hd__or3_1 U4268 (.A(n3619),
    .B(n3618),
    .C(n3617),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3620));
 sky130_fd_sc_hd__a22o_1 U4269 (.A1(n3666),
    .A2(n3620),
    .B1(n3664),
    .B2(net226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1758));
 sky130_fd_sc_hd__a22o_1 U4270 (.A1(n3668),
    .A2(net270),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[121] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1757));
 sky130_fd_sc_hd__a22o_1 U4271 (.A1(n3670),
    .A2(net271),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[113] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1756));
 sky130_fd_sc_hd__a22o_1 U4272 (.A1(n3672),
    .A2(net271),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[105] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1755));
 sky130_fd_sc_hd__a22o_1 U4273 (.A1(n3674),
    .A2(net271),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[97] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1754));
 sky130_fd_sc_hd__a22o_1 U4274 (.A1(n3676),
    .A2(net271),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[89] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1753));
 sky130_fd_sc_hd__a22o_1 U4275 (.A1(n3678),
    .A2(net271),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[81] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1752));
 sky130_fd_sc_hd__a22o_1 U4276 (.A1(n3680),
    .A2(net271),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[73] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1751));
 sky130_fd_sc_hd__a22o_1 U4277 (.A1(n3682),
    .A2(net271),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[65] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1750));
 sky130_fd_sc_hd__a22o_1 U4278 (.A1(n3684),
    .A2(net271),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[57] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1749));
 sky130_fd_sc_hd__a22o_1 U4279 (.A1(n3686),
    .A2(net271),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[49] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1748));
 sky130_fd_sc_hd__a22o_1 U4280 (.A1(n3688),
    .A2(net271),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[41] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1747));
 sky130_fd_sc_hd__a22o_1 U4281 (.A1(n3690),
    .A2(net271),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[33] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1746));
 sky130_fd_sc_hd__a22o_1 U4282 (.A1(n3692),
    .A2(net271),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[25] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1745));
 sky130_fd_sc_hd__a22o_1 U4283 (.A1(n3694),
    .A2(net271),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[17] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1744));
 sky130_fd_sc_hd__a22o_1 U4284 (.A1(n3696),
    .A2(net271),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1743));
 sky130_fd_sc_hd__a22o_1 U4285 (.A1(n3698),
    .A2(net271),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1742));
 sky130_fd_sc_hd__a22o_1 U4286 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[26] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[50] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3625));
 sky130_fd_sc_hd__a22o_1 U4287 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[42] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[18] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3624));
 sky130_fd_sc_hd__a22o_1 U4288 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[58] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[2] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3622));
 sky130_fd_sc_hd__a22o_1 U4289 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[34] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[66] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3621));
 sky130_fd_sc_hd__a211o_1 U4290 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[10] ),
    .A2(n3660),
    .B1(n3622),
    .C1(n3621),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3623));
 sky130_fd_sc_hd__or3_1 U4291 (.A(n3625),
    .B(n3624),
    .C(n3623),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3626));
 sky130_fd_sc_hd__a22o_1 U4292 (.A1(n3666),
    .A2(n3626),
    .B1(n3664),
    .B2(net225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1741));
 sky130_fd_sc_hd__a22o_1 U4293 (.A1(n3668),
    .A2(net260),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[122] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1740));
 sky130_fd_sc_hd__a22o_1 U4294 (.A1(n3670),
    .A2(net261),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[114] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1739));
 sky130_fd_sc_hd__a22o_1 U4295 (.A1(n3672),
    .A2(net261),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[106] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1738));
 sky130_fd_sc_hd__a22o_1 U4296 (.A1(n3674),
    .A2(net261),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[98] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1737));
 sky130_fd_sc_hd__a22o_1 U4297 (.A1(n3676),
    .A2(net261),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[90] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1736));
 sky130_fd_sc_hd__a22o_1 U4298 (.A1(n3678),
    .A2(net261),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[82] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1735));
 sky130_fd_sc_hd__a22o_1 U4299 (.A1(n3680),
    .A2(net261),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[74] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1734));
 sky130_fd_sc_hd__a22o_1 U4300 (.A1(n3682),
    .A2(net261),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[66] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1733));
 sky130_fd_sc_hd__a22o_1 U4301 (.A1(n3684),
    .A2(net261),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[58] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1732));
 sky130_fd_sc_hd__a22o_1 U4302 (.A1(n3686),
    .A2(net261),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[50] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1731));
 sky130_fd_sc_hd__a22o_1 U4303 (.A1(n3688),
    .A2(net261),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[42] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1730));
 sky130_fd_sc_hd__a22o_1 U4304 (.A1(n3690),
    .A2(net261),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[34] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1729));
 sky130_fd_sc_hd__a22o_1 U4305 (.A1(n3692),
    .A2(net261),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[26] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1728));
 sky130_fd_sc_hd__a22o_1 U4306 (.A1(n3694),
    .A2(net261),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[18] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1727));
 sky130_fd_sc_hd__a22o_1 U4307 (.A1(n3696),
    .A2(net261),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1726));
 sky130_fd_sc_hd__a22o_1 U4308 (.A1(n3698),
    .A2(net261),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1725));
 sky130_fd_sc_hd__a22o_1 U4309 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[27] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[51] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3631));
 sky130_fd_sc_hd__a22o_1 U4310 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[43] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[19] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3630));
 sky130_fd_sc_hd__a22o_1 U4311 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[59] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[3] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3628));
 sky130_fd_sc_hd__a22o_1 U4312 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[35] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[67] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3627));
 sky130_fd_sc_hd__a211o_1 U4313 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[11] ),
    .A2(n3660),
    .B1(n3628),
    .C1(n3627),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3629));
 sky130_fd_sc_hd__or3_1 U4314 (.A(n3631),
    .B(n3630),
    .C(n3629),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3632));
 sky130_fd_sc_hd__a22o_1 U4315 (.A1(n3666),
    .A2(n3632),
    .B1(n3664),
    .B2(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1724));
 sky130_fd_sc_hd__a22o_1 U4316 (.A1(n3668),
    .A2(net287),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[123] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1723));
 sky130_fd_sc_hd__a22o_1 U4317 (.A1(n3670),
    .A2(net288),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[115] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1722));
 sky130_fd_sc_hd__a22o_1 U4318 (.A1(n3672),
    .A2(net288),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[107] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1721));
 sky130_fd_sc_hd__a22o_1 U4319 (.A1(n3674),
    .A2(net288),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[99] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1720));
 sky130_fd_sc_hd__a22o_1 U4320 (.A1(n3676),
    .A2(net288),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[91] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1719));
 sky130_fd_sc_hd__a22o_1 U4321 (.A1(n3678),
    .A2(net288),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[83] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1718));
 sky130_fd_sc_hd__a22o_1 U4322 (.A1(n3680),
    .A2(net288),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[75] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1717));
 sky130_fd_sc_hd__a22o_1 U4323 (.A1(n3682),
    .A2(net288),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[67] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1716));
 sky130_fd_sc_hd__a22o_1 U4324 (.A1(n3684),
    .A2(net288),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[59] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1715));
 sky130_fd_sc_hd__a22o_1 U4325 (.A1(n3686),
    .A2(net288),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[51] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1714));
 sky130_fd_sc_hd__a22o_1 U4326 (.A1(n3688),
    .A2(net288),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[43] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1713));
 sky130_fd_sc_hd__a22o_1 U4327 (.A1(n3690),
    .A2(net288),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[35] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1712));
 sky130_fd_sc_hd__a22o_1 U4328 (.A1(n3692),
    .A2(net288),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[27] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1711));
 sky130_fd_sc_hd__a22o_1 U4329 (.A1(n3694),
    .A2(net288),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[19] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1710));
 sky130_fd_sc_hd__a22o_1 U4330 (.A1(n3696),
    .A2(net288),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1709));
 sky130_fd_sc_hd__a22o_1 U4331 (.A1(n3698),
    .A2(net288),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1708));
 sky130_fd_sc_hd__a22o_1 U4332 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[28] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[52] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3637));
 sky130_fd_sc_hd__a22o_1 U4333 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[44] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[20] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3636));
 sky130_fd_sc_hd__a22o_1 U4334 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[60] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[4] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3634));
 sky130_fd_sc_hd__a22o_1 U4335 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[36] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[68] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3633));
 sky130_fd_sc_hd__a211o_1 U4336 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[12] ),
    .A2(n3660),
    .B1(n3634),
    .C1(n3633),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3635));
 sky130_fd_sc_hd__or3_1 U4337 (.A(n3637),
    .B(n3636),
    .C(n3635),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3638));
 sky130_fd_sc_hd__a22o_1 U4338 (.A1(n3666),
    .A2(n3638),
    .B1(n3664),
    .B2(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1707));
 sky130_fd_sc_hd__a22o_1 U4339 (.A1(n3668),
    .A2(net256),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[124] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1706));
 sky130_fd_sc_hd__a22o_1 U4340 (.A1(n3670),
    .A2(net257),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[116] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1705));
 sky130_fd_sc_hd__a22o_1 U4341 (.A1(n3672),
    .A2(net257),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[108] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1704));
 sky130_fd_sc_hd__a22o_1 U4342 (.A1(n3674),
    .A2(net257),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[100] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1703));
 sky130_fd_sc_hd__a22o_1 U4343 (.A1(n3676),
    .A2(net257),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[92] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1702));
 sky130_fd_sc_hd__a22o_1 U4344 (.A1(n3678),
    .A2(net257),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[84] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1701));
 sky130_fd_sc_hd__a22o_1 U4345 (.A1(n3680),
    .A2(net257),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[76] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1700));
 sky130_fd_sc_hd__a22o_1 U4346 (.A1(n3682),
    .A2(net257),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[68] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1699));
 sky130_fd_sc_hd__a22o_1 U4347 (.A1(n3684),
    .A2(net257),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[60] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1698));
 sky130_fd_sc_hd__a22o_1 U4348 (.A1(n3686),
    .A2(net257),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[52] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1697));
 sky130_fd_sc_hd__a22o_1 U4349 (.A1(n3688),
    .A2(net257),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[44] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1696));
 sky130_fd_sc_hd__a22o_1 U4350 (.A1(n3690),
    .A2(net257),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[36] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1695));
 sky130_fd_sc_hd__a22o_1 U4351 (.A1(n3692),
    .A2(net257),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[28] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1694));
 sky130_fd_sc_hd__a22o_1 U4352 (.A1(n3694),
    .A2(net257),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[20] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1693));
 sky130_fd_sc_hd__a22o_1 U4353 (.A1(n3696),
    .A2(net257),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1692));
 sky130_fd_sc_hd__a22o_1 U4354 (.A1(n3698),
    .A2(net257),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1691));
 sky130_fd_sc_hd__a22o_1 U4355 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[29] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[53] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3643));
 sky130_fd_sc_hd__a22o_1 U4356 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[45] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[21] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3642));
 sky130_fd_sc_hd__a22o_1 U4357 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[61] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[5] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3640));
 sky130_fd_sc_hd__a22o_1 U4358 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[37] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[69] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3639));
 sky130_fd_sc_hd__a211o_1 U4359 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[13] ),
    .A2(n3660),
    .B1(n3640),
    .C1(n3639),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3641));
 sky130_fd_sc_hd__or3_1 U4360 (.A(n3643),
    .B(n3642),
    .C(n3641),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3644));
 sky130_fd_sc_hd__a22o_1 U4361 (.A1(n3666),
    .A2(n3644),
    .B1(n3664),
    .B2(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1690));
 sky130_fd_sc_hd__a22o_1 U4362 (.A1(n3668),
    .A2(net274),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[125] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1689));
 sky130_fd_sc_hd__a22o_1 U4363 (.A1(n3670),
    .A2(net275),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[117] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1688));
 sky130_fd_sc_hd__a22o_1 U4364 (.A1(n3672),
    .A2(net275),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[109] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1687));
 sky130_fd_sc_hd__a22o_1 U4365 (.A1(n3674),
    .A2(net275),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[101] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1686));
 sky130_fd_sc_hd__a22o_1 U4366 (.A1(n3676),
    .A2(net275),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[93] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1685));
 sky130_fd_sc_hd__a22o_1 U4367 (.A1(n3678),
    .A2(net275),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[85] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1684));
 sky130_fd_sc_hd__a22o_1 U4368 (.A1(n3680),
    .A2(net275),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[77] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1683));
 sky130_fd_sc_hd__a22o_1 U4369 (.A1(n3682),
    .A2(net275),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[69] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1682));
 sky130_fd_sc_hd__a22o_1 U4370 (.A1(n3684),
    .A2(net275),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[61] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1681));
 sky130_fd_sc_hd__a22o_1 U4371 (.A1(n3686),
    .A2(net275),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[53] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1680));
 sky130_fd_sc_hd__a22o_1 U4372 (.A1(n3688),
    .A2(net275),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[45] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1679));
 sky130_fd_sc_hd__a22o_1 U4373 (.A1(n3690),
    .A2(net275),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[37] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1678));
 sky130_fd_sc_hd__a22o_1 U4374 (.A1(n3692),
    .A2(net275),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[29] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1677));
 sky130_fd_sc_hd__a22o_1 U4375 (.A1(n3694),
    .A2(net275),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[21] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1676));
 sky130_fd_sc_hd__a22o_1 U4376 (.A1(n3696),
    .A2(net275),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1675));
 sky130_fd_sc_hd__a22o_1 U4377 (.A1(n3698),
    .A2(net275),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1674));
 sky130_fd_sc_hd__a22o_1 U4378 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[30] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[54] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3649));
 sky130_fd_sc_hd__a22o_1 U4379 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[46] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[22] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3648));
 sky130_fd_sc_hd__a22o_1 U4380 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[62] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[6] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3646));
 sky130_fd_sc_hd__a22o_1 U4381 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[38] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[70] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3645));
 sky130_fd_sc_hd__a211o_1 U4382 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[14] ),
    .A2(n3660),
    .B1(n3646),
    .C1(n3645),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3647));
 sky130_fd_sc_hd__or3_1 U4383 (.A(n3649),
    .B(n3648),
    .C(n3647),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3650));
 sky130_fd_sc_hd__a22o_1 U4384 (.A1(n3666),
    .A2(n3650),
    .B1(n3664),
    .B2(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1673));
 sky130_fd_sc_hd__a22o_1 U4385 (.A1(n3668),
    .A2(net177),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[126] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1672));
 sky130_fd_sc_hd__a22o_1 U4386 (.A1(n3670),
    .A2(net178),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[118] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1671));
 sky130_fd_sc_hd__a22o_1 U4387 (.A1(n3672),
    .A2(net178),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[110] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1670));
 sky130_fd_sc_hd__a22o_1 U4388 (.A1(n3674),
    .A2(net178),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[102] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1669));
 sky130_fd_sc_hd__a22o_1 U4389 (.A1(n3676),
    .A2(net178),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[94] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1668));
 sky130_fd_sc_hd__a22o_1 U4390 (.A1(n3678),
    .A2(net178),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[86] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1667));
 sky130_fd_sc_hd__a22o_1 U4391 (.A1(n3680),
    .A2(net178),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[78] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1666));
 sky130_fd_sc_hd__a22o_1 U4392 (.A1(n3682),
    .A2(net178),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[70] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1665));
 sky130_fd_sc_hd__a22o_1 U4393 (.A1(n3684),
    .A2(net178),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[62] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1664));
 sky130_fd_sc_hd__a22o_1 U4394 (.A1(n3686),
    .A2(net178),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[54] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1663));
 sky130_fd_sc_hd__a22o_1 U4395 (.A1(n3688),
    .A2(net178),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[46] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1662));
 sky130_fd_sc_hd__a22o_1 U4396 (.A1(n3690),
    .A2(net178),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[38] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1661));
 sky130_fd_sc_hd__a22o_1 U4397 (.A1(n3692),
    .A2(net178),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[30] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1660));
 sky130_fd_sc_hd__a22o_1 U4398 (.A1(n3694),
    .A2(net178),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[22] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1659));
 sky130_fd_sc_hd__a22o_1 U4399 (.A1(n3696),
    .A2(net178),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1658));
 sky130_fd_sc_hd__a22o_1 U4400 (.A1(n3698),
    .A2(net178),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1657));
 sky130_fd_sc_hd__a22o_1 U4401 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[31] ),
    .A2(n3652),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[55] ),
    .B2(n3651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3663));
 sky130_fd_sc_hd__a22o_1 U4402 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[47] ),
    .A2(n3654),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[23] ),
    .B2(n3653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3662));
 sky130_fd_sc_hd__a22o_1 U4403 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[63] ),
    .A2(n3655),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[7] ),
    .B2(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3659));
 sky130_fd_sc_hd__a22o_1 U4404 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[39] ),
    .A2(n3657),
    .B1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[71] ),
    .B2(n3656),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3658));
 sky130_fd_sc_hd__a211o_1 U4405 (.A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[15] ),
    .A2(n3660),
    .B1(n3659),
    .C1(n3658),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3661));
 sky130_fd_sc_hd__or3_1 U4406 (.A(n3663),
    .B(n3662),
    .C(n3661),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3665));
 sky130_fd_sc_hd__a22o_1 U4407 (.A1(n3666),
    .A2(n3665),
    .B1(n3664),
    .B2(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1656));
 sky130_fd_sc_hd__a22o_1 U4408 (.A1(n3668),
    .A2(net245),
    .B1(n3667),
    .B2(\inst_to_wrap_rx_fifo_array_reg[127] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1655));
 sky130_fd_sc_hd__a22o_1 U4409 (.A1(n3670),
    .A2(net246),
    .B1(n3669),
    .B2(\inst_to_wrap_rx_fifo_array_reg[119] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1654));
 sky130_fd_sc_hd__a22o_1 U4410 (.A1(n3672),
    .A2(net246),
    .B1(n3671),
    .B2(\inst_to_wrap_rx_fifo_array_reg[111] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1653));
 sky130_fd_sc_hd__a22o_1 U4411 (.A1(n3674),
    .A2(net246),
    .B1(n3673),
    .B2(\inst_to_wrap_rx_fifo_array_reg[103] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1652));
 sky130_fd_sc_hd__a22o_1 U4412 (.A1(n3676),
    .A2(net246),
    .B1(n3675),
    .B2(\inst_to_wrap_rx_fifo_array_reg[95] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1651));
 sky130_fd_sc_hd__a22o_1 U4413 (.A1(n3678),
    .A2(net246),
    .B1(n3677),
    .B2(\inst_to_wrap_rx_fifo_array_reg[87] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1650));
 sky130_fd_sc_hd__a22o_1 U4414 (.A1(n3680),
    .A2(net246),
    .B1(n3679),
    .B2(\inst_to_wrap_rx_fifo_array_reg[79] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1649));
 sky130_fd_sc_hd__a22o_1 U4415 (.A1(n3682),
    .A2(net246),
    .B1(n3681),
    .B2(\inst_to_wrap_rx_fifo_array_reg[71] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1648));
 sky130_fd_sc_hd__a22o_1 U4416 (.A1(n3684),
    .A2(net246),
    .B1(n3683),
    .B2(\inst_to_wrap_rx_fifo_array_reg[63] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1647));
 sky130_fd_sc_hd__a22o_1 U4417 (.A1(n3686),
    .A2(net246),
    .B1(n3685),
    .B2(\inst_to_wrap_rx_fifo_array_reg[55] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1646));
 sky130_fd_sc_hd__a22o_1 U4418 (.A1(n3688),
    .A2(net246),
    .B1(n3687),
    .B2(\inst_to_wrap_rx_fifo_array_reg[47] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1645));
 sky130_fd_sc_hd__a22o_1 U4419 (.A1(n3690),
    .A2(net246),
    .B1(n3689),
    .B2(\inst_to_wrap_rx_fifo_array_reg[39] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1644));
 sky130_fd_sc_hd__a22o_1 U4420 (.A1(n3692),
    .A2(net246),
    .B1(n3691),
    .B2(\inst_to_wrap_rx_fifo_array_reg[31] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1643));
 sky130_fd_sc_hd__a22o_1 U4421 (.A1(n3694),
    .A2(net246),
    .B1(n3693),
    .B2(\inst_to_wrap_rx_fifo_array_reg[23] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1642));
 sky130_fd_sc_hd__a22o_1 U4422 (.A1(n3696),
    .A2(net246),
    .B1(n3695),
    .B2(\inst_to_wrap_rx_fifo_array_reg[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1641));
 sky130_fd_sc_hd__a22o_1 U4423 (.A1(n3698),
    .A2(net246),
    .B1(n3697),
    .B2(\inst_to_wrap_rx_fifo_array_reg[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1640));
 sky130_fd_sc_hd__inv_2 U4424 (.A(net244),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3699));
 sky130_fd_sc_hd__a22o_1 U4425 (.A1(net17),
    .A2(net7),
    .B1(n3699),
    .B2(\last_HADDR[15] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1639));
 sky130_fd_sc_hd__a22o_1 U4426 (.A1(net244),
    .A2(net6),
    .B1(n3699),
    .B2(\last_HADDR[14] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1638));
 sky130_fd_sc_hd__a22o_1 U4427 (.A1(net244),
    .A2(net5),
    .B1(n3699),
    .B2(\last_HADDR[13] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1637));
 sky130_fd_sc_hd__a22o_1 U4428 (.A1(net244),
    .A2(net4),
    .B1(net231),
    .B2(\last_HADDR[12] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1636));
 sky130_fd_sc_hd__a22o_1 U4429 (.A1(net244),
    .A2(net3),
    .B1(net231),
    .B2(\last_HADDR[11] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1635));
 sky130_fd_sc_hd__a22o_1 U4430 (.A1(net244),
    .A2(net2),
    .B1(net231),
    .B2(\last_HADDR[10] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1634));
 sky130_fd_sc_hd__a22o_1 U4431 (.A1(net244),
    .A2(net16),
    .B1(net231),
    .B2(\last_HADDR[9] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1633));
 sky130_fd_sc_hd__a22o_1 U4432 (.A1(net244),
    .A2(net15),
    .B1(net231),
    .B2(\last_HADDR[8] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1632));
 sky130_fd_sc_hd__a22o_1 U4433 (.A1(net17),
    .A2(net14),
    .B1(net231),
    .B2(\last_HADDR[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1631));
 sky130_fd_sc_hd__a22o_1 U4434 (.A1(net244),
    .A2(net13),
    .B1(net231),
    .B2(\last_HADDR[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1630));
 sky130_fd_sc_hd__a22o_1 U4435 (.A1(net244),
    .A2(net12),
    .B1(net231),
    .B2(\last_HADDR[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1629));
 sky130_fd_sc_hd__a22o_1 U4436 (.A1(net17),
    .A2(net11),
    .B1(net231),
    .B2(\last_HADDR[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1628));
 sky130_fd_sc_hd__a22o_1 U4437 (.A1(net17),
    .A2(net10),
    .B1(net231),
    .B2(\last_HADDR[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1627));
 sky130_fd_sc_hd__a22o_1 U4438 (.A1(net244),
    .A2(net9),
    .B1(net231),
    .B2(\last_HADDR[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1626));
 sky130_fd_sc_hd__a22o_1 U4439 (.A1(net244),
    .A2(net8),
    .B1(net231),
    .B2(\last_HADDR[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1625));
 sky130_fd_sc_hd__a22o_1 U4440 (.A1(net244),
    .A2(net1),
    .B1(net231),
    .B2(\last_HADDR[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1624));
 sky130_fd_sc_hd__a22o_1 U4441 (.A1(net244),
    .A2(net28),
    .B1(net231),
    .B2(last_HWRITE),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1623));
 sky130_fd_sc_hd__a22o_1 U4442 (.A1(net244),
    .A2(net19),
    .B1(net231),
    .B2(last_HTRANS_1_),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1622));
 sky130_fd_sc_hd__a22o_1 U4443 (.A1(net244),
    .A2(net18),
    .B1(net231),
    .B2(last_HSEL),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1621));
 sky130_fd_sc_hd__nand2_1 U4444 (.A(n3713),
    .B(n3700),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3701));
 sky130_fd_sc_hd__inv_2 U4445 (.A(n3701),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3702));
 sky130_fd_sc_hd__a22o_1 U4446 (.A1(n3702),
    .A2(net23),
    .B1(n3701),
    .B2(\tx_fifo_th[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1620));
 sky130_fd_sc_hd__a22o_1 U4447 (.A1(n3702),
    .A2(net22),
    .B1(n3701),
    .B2(\tx_fifo_th[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1619));
 sky130_fd_sc_hd__a22o_1 U4448 (.A1(n3702),
    .A2(net21),
    .B1(n3701),
    .B2(\tx_fifo_th[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1618));
 sky130_fd_sc_hd__a22o_1 U4449 (.A1(n3702),
    .A2(net237),
    .B1(n3701),
    .B2(\tx_fifo_th[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1617));
 sky130_fd_sc_hd__nand2_2 U4450 (.A(n3713),
    .B(n3703),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3704));
 sky130_fd_sc_hd__inv_2 U4451 (.A(n3704),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3705));
 sky130_fd_sc_hd__a22o_1 U4452 (.A1(n3705),
    .A2(net234),
    .B1(n3704),
    .B2(\rx_fifo_th[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1616));
 sky130_fd_sc_hd__a22o_1 U4453 (.A1(n3705),
    .A2(net235),
    .B1(n3704),
    .B2(\rx_fifo_th[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1615));
 sky130_fd_sc_hd__a22o_1 U4454 (.A1(n3705),
    .A2(net236),
    .B1(n3704),
    .B2(\rx_fifo_th[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1614));
 sky130_fd_sc_hd__a22o_1 U4455 (.A1(n3705),
    .A2(net20),
    .B1(n3704),
    .B2(\rx_fifo_th[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1613));
 sky130_fd_sc_hd__and3_1 U4456 (.A(\last_HADDR[4] ),
    .B(\last_HADDR[3] ),
    .C(n3706),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3707));
 sky130_fd_sc_hd__mux2_1 U4457 (.A0(CONTROL_REG_0_),
    .A1(net20),
    .S(n3707),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1612));
 sky130_fd_sc_hd__and3_2 U4458 (.A(n3713),
    .B(n3709),
    .C(n3708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3711));
 sky130_fd_sc_hd__inv_2 U4459 (.A(n3711),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3710));
 sky130_fd_sc_hd__a22o_1 U4460 (.A1(n3711),
    .A2(net232),
    .B1(n3710),
    .B2(\IM_REG[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1611));
 sky130_fd_sc_hd__a22o_1 U4461 (.A1(n3711),
    .A2(net233),
    .B1(n3710),
    .B2(\IM_REG[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1610));
 sky130_fd_sc_hd__a22o_1 U4462 (.A1(n3711),
    .A2(net234),
    .B1(n3710),
    .B2(\IM_REG[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1609));
 sky130_fd_sc_hd__a22o_1 U4463 (.A1(n3711),
    .A2(net235),
    .B1(n3710),
    .B2(\IM_REG[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1608));
 sky130_fd_sc_hd__a22o_1 U4464 (.A1(n3711),
    .A2(net236),
    .B1(n3710),
    .B2(\IM_REG[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1607));
 sky130_fd_sc_hd__a22o_1 U4465 (.A1(n3711),
    .A2(net20),
    .B1(n3710),
    .B2(\IM_REG[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1606));
 sky130_fd_sc_hd__nand2_1 U4466 (.A(n3713),
    .B(n3712),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3714));
 sky130_fd_sc_hd__mux2_1 U4467 (.A0(net20),
    .A1(CG_REG_0_),
    .S(n3714),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1605));
 sky130_fd_sc_hd__a22o_1 U4468 (.A1(n3825),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[0] ),
    .B1(n3826),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1604));
 sky130_fd_sc_hd__a22o_1 U4469 (.A1(n3825),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[0] ),
    .B1(n3826),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1603));
 sky130_fd_sc_hd__a22o_1 U4470 (.A1(n3825),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ),
    .B1(n3826),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1602));
 sky130_fd_sc_hd__a22o_1 U4471 (.A1(n3825),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[2] ),
    .B1(n3826),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1601));
 sky130_fd_sc_hd__and2_1 U4472 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[1] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3721));
 sky130_fd_sc_hd__inv_1 U4473 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3720));
 sky130_fd_sc_hd__a31o_1 U4474 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[1] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[2] ),
    .A3(n3792),
    .B1(n3715),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3828));
 sky130_fd_sc_hd__a221o_1 U4475 (.A1(n3718),
    .A2(n3717),
    .B1(n3718),
    .B2(n3716),
    .C1(n3828),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3719));
 sky130_fd_sc_hd__nor2_1 U4476 (.A(n3793),
    .B(n3719),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3791));
 sky130_fd_sc_hd__inv_2 U4477 (.A(n3793),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3829));
 sky130_fd_sc_hd__o21ai_1 U4478 (.A1(n3721),
    .A2(n3719),
    .B1(n3829),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3794));
 sky130_fd_sc_hd__a32o_1 U4479 (.A1(n3721),
    .A2(n3720),
    .A3(n3791),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[2] ),
    .B2(n3794),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1600));
 sky130_fd_sc_hd__o31a_1 U4480 (.A1(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ),
    .A2(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[0] ),
    .A3(inst_to_wrap_u_usb_cdc_u_ctrl_endp_usb_reset_q),
    .B1(n3722),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3723));
 sky130_fd_sc_hd__and3_1 U4481 (.A(n3825),
    .B(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q),
    .C(n3723),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3763));
 sky130_fd_sc_hd__inv_2 U4482 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3759));
 sky130_fd_sc_hd__inv_2 U4483 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3725));
 sky130_fd_sc_hd__a22o_1 U4484 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[2] ),
    .A2(n3725),
    .B1(n3752),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3724));
 sky130_fd_sc_hd__a221o_1 U4485 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ),
    .A2(n3759),
    .B1(n3746),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[1] ),
    .C1(n3724),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3750));
 sky130_fd_sc_hd__o21ai_1 U4486 (.A1(n3752),
    .A2(n3746),
    .B1(n3756),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3821));
 sky130_fd_sc_hd__a21o_1 U4487 (.A1(n3759),
    .A2(n3725),
    .B1(n3821),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3819));
 sky130_fd_sc_hd__nor2_1 U4488 (.A(n3734),
    .B(n3819),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3820));
 sky130_fd_sc_hd__inv_2 U4489 (.A(n3820),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3739));
 sky130_fd_sc_hd__or2_1 U4490 (.A(n3746),
    .B(n3752),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3729));
 sky130_fd_sc_hd__inv_2 U4491 (.A(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3737));
 sky130_fd_sc_hd__or4_1 U4492 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_0_),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[0] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[1] ),
    .D(n3737),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3726));
 sky130_fd_sc_hd__or4_1 U4493 (.A(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[5] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[4] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[3] ),
    .D(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3745));
 sky130_fd_sc_hd__or3b_1 U4494 (.A(n3726),
    .B(n3745),
    .C_N(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3757));
 sky130_fd_sc_hd__a21o_1 U4495 (.A1(n3776),
    .A2(n3757),
    .B1(n3756),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3748));
 sky130_fd_sc_hd__inv_1 U4496 (.A(n3748),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3727));
 sky130_fd_sc_hd__a221o_1 U4497 (.A1(n3756),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[1] ),
    .B1(n3756),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[0] ),
    .C1(n3727),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3728));
 sky130_fd_sc_hd__o211a_1 U4498 (.A1(n3750),
    .A2(n3739),
    .B1(n3729),
    .C1(n3728),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3733));
 sky130_fd_sc_hd__or2_1 U4499 (.A(n3736),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3818));
 sky130_fd_sc_hd__inv_2 U4500 (.A(n3784),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3753));
 sky130_fd_sc_hd__or2_1 U4501 (.A(n3779),
    .B(n3736),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3730));
 sky130_fd_sc_hd__o22a_1 U4502 (.A1(n3753),
    .A2(n3760),
    .B1(n3731),
    .B2(n3730),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3732));
 sky130_fd_sc_hd__o21ai_1 U4503 (.A1(n3733),
    .A2(n3818),
    .B1(n3732),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3785));
 sky130_fd_sc_hd__a22o_1 U4504 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .A2(n3826),
    .B1(n3763),
    .B2(n3785),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1599));
 sky130_fd_sc_hd__nor2_1 U4505 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_0_),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3735));
 sky130_fd_sc_hd__nand2b_1 U4506 (.A_N(n3819),
    .B(n3734),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3747));
 sky130_fd_sc_hd__o22a_1 U4507 (.A1(n3735),
    .A2(n3747),
    .B1(n3776),
    .B2(n3756),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3738));
 sky130_fd_sc_hd__or3_2 U4508 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[0] ),
    .C(n3736),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3755));
 sky130_fd_sc_hd__inv_2 U4509 (.A(n3750),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3822));
 sky130_fd_sc_hd__or2_1 U4510 (.A(n3779),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3823));
 sky130_fd_sc_hd__or4_1 U4511 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .B(n3822),
    .C(n3823),
    .D(n3821),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3754));
 sky130_fd_sc_hd__o22a_1 U4512 (.A1(n3738),
    .A2(n3755),
    .B1(n3737),
    .B2(n3754),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3740));
 sky130_fd_sc_hd__or2_1 U4513 (.A(n3739),
    .B(n3822),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3749));
 sky130_fd_sc_hd__o21ai_4 U4514 (.A1(n3749),
    .A2(n3755),
    .B1(n3825),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3743));
 sky130_fd_sc_hd__or2_1 U4515 (.A(n3747),
    .B(n3755),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3767));
 sky130_fd_sc_hd__o21a_1 U4516 (.A1(n3767),
    .A2(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_0_),
    .B1(n3754),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3741));
 sky130_fd_sc_hd__nor2_2 U4517 (.A(n3826),
    .B(n3741),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3742));
 sky130_fd_sc_hd__a22o_1 U4518 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[6] ),
    .A2(n3742),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[5] ),
    .B2(n3743),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1597));
 sky130_fd_sc_hd__a22o_1 U4519 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[5] ),
    .A2(n3742),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[4] ),
    .B2(n3743),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1596));
 sky130_fd_sc_hd__a22o_1 U4520 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[4] ),
    .A2(n3742),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[3] ),
    .B2(n3743),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1595));
 sky130_fd_sc_hd__a22o_1 U4521 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[3] ),
    .A2(n3742),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[2] ),
    .B2(n3743),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1594));
 sky130_fd_sc_hd__a22o_1 U4522 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[2] ),
    .A2(n3742),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[1] ),
    .B2(n3743),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1593));
 sky130_fd_sc_hd__a22o_1 U4523 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[0] ),
    .A2(n3743),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[1] ),
    .B2(n3742),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1592));
 sky130_fd_sc_hd__a22o_1 U4524 (.A1(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_0_),
    .A2(n3743),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[0] ),
    .B2(n3742),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1591));
 sky130_fd_sc_hd__or4_1 U4525 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .B(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[6] ),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ),
    .D(n3823),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3744));
 sky130_fd_sc_hd__or4_1 U4526 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[2] ),
    .B(n3746),
    .C(n3745),
    .D(n3744),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3768));
 sky130_fd_sc_hd__a31o_1 U4527 (.A1(n3749),
    .A2(n3748),
    .A3(n3747),
    .B1(n3755),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3783));
 sky130_fd_sc_hd__o21ai_1 U4528 (.A1(n3750),
    .A2(n3768),
    .B1(n3783),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3751));
 sky130_fd_sc_hd__a22o_1 U4529 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[1] ),
    .A2(n3826),
    .B1(n3763),
    .B2(n3751),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1590));
 sky130_fd_sc_hd__and4_1 U4530 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ),
    .B(n3753),
    .C(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[0] ),
    .D(n3752),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3761));
 sky130_fd_sc_hd__o31ai_1 U4531 (.A1(n3757),
    .A2(n3756),
    .A3(n3755),
    .B1(n3754),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3758));
 sky130_fd_sc_hd__a31o_1 U4532 (.A1(n3761),
    .A2(n3760),
    .A3(n3759),
    .B1(n3758),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3762));
 sky130_fd_sc_hd__a22o_1 U4533 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[0] ),
    .A2(n3826),
    .B1(n3763),
    .B2(n3762),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1589));
 sky130_fd_sc_hd__nand2_1 U4534 (.A(n3825),
    .B(n3822),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3766));
 sky130_fd_sc_hd__nor2_1 U4535 (.A(n3768),
    .B(n3766),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3764));
 sky130_fd_sc_hd__mux2_1 U4536 (.A0(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq),
    .A1(n3765),
    .S(n3764),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1588));
 sky130_fd_sc_hd__inv_2 U4537 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3770));
 sky130_fd_sc_hd__a21oi_1 U4538 (.A1(n3768),
    .A2(n3767),
    .B1(n3766),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3773));
 sky130_fd_sc_hd__a22o_1 U4539 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[0] ),
    .A2(n3826),
    .B1(n3770),
    .B2(n3773),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1587));
 sky130_fd_sc_hd__o21ai_1 U4540 (.A1(n3771),
    .A2(n3770),
    .B1(n3773),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3769));
 sky130_fd_sc_hd__nand2_1 U4541 (.A(n3825),
    .B(n3769),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3772));
 sky130_fd_sc_hd__a32o_1 U4542 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[0] ),
    .A2(n3771),
    .A3(n3773),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[1] ),
    .B2(n3772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1586));
 sky130_fd_sc_hd__nor2_1 U4543 (.A(n3771),
    .B(n3770),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3775));
 sky130_fd_sc_hd__a32o_1 U4544 (.A1(n3775),
    .A2(n3774),
    .A3(n3773),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[2] ),
    .B2(n3772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1585));
 sky130_fd_sc_hd__a211o_1 U4545 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[1] ),
    .A2(n3780),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .C1(n3779),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3782));
 sky130_fd_sc_hd__a31o_1 U4546 (.A1(n3784),
    .A2(n3783),
    .A3(n3782),
    .B1(n3781),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3787));
 sky130_fd_sc_hd__o21ai_1 U4547 (.A1(n3785),
    .A2(n3788),
    .B1(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3786));
 sky130_fd_sc_hd__o21ai_1 U4548 (.A1(n3788),
    .A2(n3787),
    .B1(n3786),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3789));
 sky130_fd_sc_hd__a22o_1 U4549 (.A1(n3825),
    .A2(n3789),
    .B1(n3826),
    .B2(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_fq),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1584));
 sky130_fd_sc_hd__a22o_1 U4550 (.A1(n3829),
    .A2(n3790),
    .B1(n3793),
    .B2(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1583));
 sky130_fd_sc_hd__a22o_1 U4551 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[0] ),
    .A2(n3793),
    .B1(n3792),
    .B2(n3791),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1582));
 sky130_fd_sc_hd__a32o_1 U4552 (.A1(n3794),
    .A2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[0] ),
    .A3(n3829),
    .B1(n3794),
    .B2(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1581));
 sky130_fd_sc_hd__and2_1 U4553 (.A(n3795),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3809));
 sky130_fd_sc_hd__o21ai_1 U4554 (.A1(n3811),
    .A2(n3809),
    .B1(n3810),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3808));
 sky130_fd_sc_hd__a32o_1 U4555 (.A1(n3798),
    .A2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ),
    .A3(n3797),
    .B1(n3796),
    .B2(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3805));
 sky130_fd_sc_hd__or2_1 U4556 (.A(n3799),
    .B(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3801));
 sky130_fd_sc_hd__a22oi_1 U4557 (.A1(n3806),
    .A2(n3805),
    .B1(n3804),
    .B2(n3803),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3802));
 sky130_fd_sc_hd__o221a_1 U4558 (.A1(n3806),
    .A2(n3805),
    .B1(n3804),
    .B2(n3803),
    .C1(n3802),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3807));
 sky130_fd_sc_hd__o311a_1 U4559 (.A1(n3810),
    .A2(n3811),
    .A3(n3809),
    .B1(n3808),
    .C1(n3807),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3817));
 sky130_fd_sc_hd__inv_1 U4560 (.A(n3814),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3816));
 sky130_fd_sc_hd__nor2_1 U4561 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ),
    .B(n3811),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3812));
 sky130_fd_sc_hd__mux2_1 U4562 (.A0(n3813),
    .A1(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ),
    .S(n3812),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3815));
 sky130_fd_sc_hd__a32o_1 U4563 (.A1(n3817),
    .A2(n3816),
    .A3(n3815),
    .B1(n3814),
    .B2(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_full_o),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1580));
 sky130_fd_sc_hd__a211o_1 U4564 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ),
    .A2(n3820),
    .B1(n3819),
    .C1(n3818),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3824));
 sky130_fd_sc_hd__a211o_1 U4565 (.A1(n3824),
    .A2(n3823),
    .B1(n3822),
    .C1(n3821),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3827));
 sky130_fd_sc_hd__o32a_1 U4566 (.A1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ),
    .A2(n3827),
    .A3(n3826),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ),
    .B2(n3825),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1578));
 sky130_fd_sc_hd__nand2_1 U4567 (.A(n3829),
    .B(n3828),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3833));
 sky130_fd_sc_hd__nor2_1 U4568 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q),
    .B(n3830),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3832));
 sky130_fd_sc_hd__nor2_1 U4569 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q),
    .B(n3833),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Y(n3831));
 sky130_fd_sc_hd__a221o_1 U4570 (.A1(n3833),
    .A2(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q),
    .B1(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ),
    .B2(n3832),
    .C1(n3831),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n3834));
 sky130_fd_sc_hd__a211o_1 U4571 (.A1(n3837),
    .A2(n3836),
    .B1(n3835),
    .C1(n3834),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(n1577));
 sky130_fd_sc_hd__buf_6 eco_cell (.A(eco_net),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net31));
 sky130_fd_sc_hd__buf_6 eco_cell_0 (.A(eco_net_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net40));
 sky130_fd_sc_hd__buf_1 eco_cell_10_0 (.A(eco_net_10_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net33));
 sky130_fd_sc_hd__buf_1 eco_cell_11_0 (.A(eco_net_11_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net34));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_12_0 (.A(eco_net_12_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net35));
 sky130_fd_sc_hd__buf_12 eco_cell_13_0 (.A(eco_net_13_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[14]));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_14_0 (.A(eco_net_14_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_15_0 (.A(eco_net_15_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net37));
 sky130_fd_sc_hd__buf_12 eco_cell_16_0 (.A(eco_net_16_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[17]));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_17_0 (.A(eco_net_17_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_18_0 (.A(eco_net_18_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net39));
 sky130_fd_sc_hd__buf_12 eco_cell_19_0 (.A(eco_net_19_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[20]));
 sky130_fd_sc_hd__buf_6 eco_cell_1_0 (.A(eco_net_1_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_20_0 (.A(eco_net_20_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net41));
 sky130_fd_sc_hd__buf_12 eco_cell_21_0 (.A(eco_net_21_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[22]));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_22_0 (.A(eco_net_22_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net42));
 sky130_fd_sc_hd__buf_12 eco_cell_23_0 (.A(eco_net_23_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[24]));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_24_0 (.A(eco_net_24_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_25_0 (.A(eco_net_25_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_26_0 (.A(eco_net_26_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_27_0 (.A(eco_net_27_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net46));
 sky130_fd_sc_hd__buf_12 eco_cell_28_0 (.A(eco_net_28_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[29]));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_29_0 (.A(eco_net_29_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net48));
 sky130_fd_sc_hd__buf_6 eco_cell_2_0 (.A(eco_net_2_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 eco_cell_30_0 (.A(eco_net_30_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_2 eco_cell_3_0 (.A(eco_net_3_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 eco_cell_4_0 (.A(eco_net_4_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_2 eco_cell_5_0 (.A(eco_net_5_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net53));
 sky130_fd_sc_hd__buf_6 eco_cell_6_0 (.A(eco_net_6_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net54));
 sky130_fd_sc_hd__buf_12 eco_cell_7_0 (.A(eco_net_7_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[8]));
 sky130_fd_sc_hd__buf_1 eco_cell_8_0 (.A(eco_net_8_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net55));
 sky130_fd_sc_hd__buf_6 eco_cell_9_0 (.A(eco_net_9_0),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net32));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__0_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1759),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__1_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1742),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__2_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1725),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__3_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1708),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__4_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1691),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__5_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1674),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__6_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1657),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_0__7_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1640),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__0_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1769),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[80] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__1_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1752),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[81] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__2_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1735),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[82] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__3_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1718),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[83] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__4_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1701),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[84] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__5_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1684),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[85] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__6_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1667),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[86] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_10__7_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1650),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[87] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__0_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1770),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[88] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__1_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1753),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[89] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__2_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1736),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[90] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__3_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1719),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[91] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__4_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1702),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[92] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__5_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1685),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[93] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__6_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1668),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[94] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_11__7_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1651),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[95] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__0_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1771),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[96] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__1_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1754),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[97] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__2_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1737),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[98] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__3_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1720),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[99] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__4_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1703),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[100] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__5_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1686),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[101] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__6_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1669),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[102] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_12__7_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1652),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[103] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__0_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1772),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[104] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__1_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1755),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[105] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__2_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1738),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[106] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__3_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1721),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[107] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__4_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1704),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[108] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__5_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1687),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[109] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__6_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1670),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[110] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_13__7_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1653),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[111] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__0_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1773),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[112] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__1_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1756),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[113] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__2_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1739),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[114] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__3_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1722),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[115] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__4_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1705),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[116] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__5_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1688),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[117] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__6_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1671),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[118] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_14__7_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1654),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[119] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__0_ (.CLK(clknet_leaf_4_HCLK),
    .D(net173),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[120] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__1_ (.CLK(clknet_leaf_5_HCLK),
    .D(net161),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[121] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__2_ (.CLK(clknet_leaf_4_HCLK),
    .D(net163),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[122] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__3_ (.CLK(clknet_leaf_5_HCLK),
    .D(net159),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[123] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__4_ (.CLK(clknet_leaf_4_HCLK),
    .D(net167),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[124] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__5_ (.CLK(clknet_leaf_4_HCLK),
    .D(net171),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[125] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__6_ (.CLK(clknet_leaf_4_HCLK),
    .D(net175),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[126] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_15__7_ (.CLK(clknet_leaf_4_HCLK),
    .D(net169),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[127] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__0_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1760),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__1_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1743),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__2_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1726),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__3_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1709),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__4_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1692),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__5_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1675),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__6_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1658),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_1__7_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1641),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__0_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1761),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__1_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1744),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__2_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1727),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__3_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1710),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[19] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__4_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1693),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[20] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__5_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1676),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[21] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__6_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1659),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[22] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_2__7_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1642),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[23] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__0_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1762),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[24] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__1_ (.CLK(clknet_leaf_3_HCLK),
    .D(net272),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[25] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__2_ (.CLK(clknet_leaf_3_HCLK),
    .D(net262),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[26] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__3_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1711),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[27] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__4_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1694),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[28] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__5_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1677),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[29] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__6_ (.CLK(clknet_leaf_3_HCLK),
    .D(net179),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[30] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_3__7_ (.CLK(clknet_leaf_3_HCLK),
    .D(net247),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[31] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__0_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1763),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[32] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__1_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1746),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[33] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__2_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1729),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[34] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__3_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1712),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[35] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__4_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1695),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[36] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__5_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1678),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[37] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__6_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1661),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[38] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_4__7_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1644),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[39] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__0_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1764),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[40] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__1_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1747),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[41] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__2_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1730),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[42] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__3_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1713),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[43] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__4_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1696),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[44] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__5_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1679),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[45] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__6_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1662),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[46] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_5__7_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1645),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[47] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__0_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1765),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[48] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__1_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1748),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[49] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__2_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1731),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[50] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__3_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1714),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[51] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__4_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1697),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[52] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__5_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1680),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[53] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__6_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1663),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[54] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_6__7_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1646),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[55] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__0_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1766),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[56] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__1_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1749),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[57] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__2_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1732),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[58] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__3_ (.CLK(clknet_leaf_4_HCLK),
    .D(n1715),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[59] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__4_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1698),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[60] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__5_ (.CLK(clknet_leaf_3_HCLK),
    .D(net276),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[61] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__6_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1664),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[62] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_7__7_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1647),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[63] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__0_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1767),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[64] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__1_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1750),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[65] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__2_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1733),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[66] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__3_ (.CLK(clknet_leaf_3_HCLK),
    .D(net289),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[67] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__4_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1699),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[68] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__5_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1682),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[69] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__6_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1665),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[70] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_8__7_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1648),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[71] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__0_ (.CLK(clknet_leaf_3_HCLK),
    .D(net254),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[72] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__1_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1751),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[73] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__2_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1734),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[74] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__3_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1717),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[75] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__4_ (.CLK(clknet_leaf_3_HCLK),
    .D(net258),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[76] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__5_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1683),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[77] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__6_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1666),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[78] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_rx_fifo_array_reg_reg_9__7_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1649),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_array_reg[79] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_rx_fifo_empty_reg_reg (.CLK(clknet_leaf_3_HCLK),
    .D(n1854),
    .SET_B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(n_RX_EMPTY_FLAG_FLAG_));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_rx_fifo_full_reg_reg (.CLK(clknet_leaf_3_HCLK),
    .D(n1848),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(n_RX_FULL_FLAG_FLAG_));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_rx_fifo_level_reg_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1853),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RXFIFOLEVEL_REG[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_rx_fifo_level_reg_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1852),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RXFIFOLEVEL_REG[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_rx_fifo_level_reg_reg_2_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1851),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RXFIFOLEVEL_REG[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_rx_fifo_level_reg_reg_3_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1850),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\RXFIFOLEVEL_REG[3] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_rx_fifo_r_ptr_reg_reg_0_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1845),
    .RESET_B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_r_ptr_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_rx_fifo_r_ptr_reg_reg_1_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1844),
    .RESET_B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_r_ptr_reg[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_rx_fifo_r_ptr_reg_reg_2_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1843),
    .RESET_B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_r_ptr_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_rx_fifo_r_ptr_reg_reg_3_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1842),
    .RESET_B(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_r_ptr_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_rx_fifo_w_ptr_reg_reg_0_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1857),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_w_ptr_reg[0] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_rx_fifo_w_ptr_reg_reg_1_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1856),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_w_ptr_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_rx_fifo_w_ptr_reg_reg_2_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1858),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_w_ptr_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_rx_fifo_w_ptr_reg_reg_3_ (.CLK(clknet_leaf_3_HCLK),
    .D(n1855),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_rx_fifo_w_ptr_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__0_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[0] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__1_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2116),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[1] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__2_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[2] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[3] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__4_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[4] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__5_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2120),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[5] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__6_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[6] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_0__7_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[7] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__0_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2043),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[80] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2036),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[81] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2037),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[82] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2038),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[83] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__4_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2039),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[84] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__5_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2040),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[85] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__6_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2041),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[86] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_10__7_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2042),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[87] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__0_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2035),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[88] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__1_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2028),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[89] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__2_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2029),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[90] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__3_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2030),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[91] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__4_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2031),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[92] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__5_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2032),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[93] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__6_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2033),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[94] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_11__7_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2034),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[95] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__0_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2027),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[96] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__1_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2020),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[97] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__2_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2021),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[98] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__3_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2022),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[99] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__4_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2023),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[100] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__5_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2024),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[101] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__6_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2025),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[102] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_12__7_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2026),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[103] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__0_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2019),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[104] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__1_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2012),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[105] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2013),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[106] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__3_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2014),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[107] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2015),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[108] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2016),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[109] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__6_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2017),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[110] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_13__7_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2018),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[111] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__0_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2011),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[112] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2004),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[113] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2005),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[114] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2006),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[115] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__4_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2007),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[116] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__5_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2008),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[117] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__6_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2009),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[118] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_14__7_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2010),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[119] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__0_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2003),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[120] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__1_ (.CLK(clknet_leaf_0_HCLK),
    .D(n1997),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[121] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__2_ (.CLK(clknet_leaf_8_HCLK),
    .D(n1998),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[122] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__3_ (.CLK(clknet_leaf_8_HCLK),
    .D(n1999),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[123] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2000),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[124] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2001),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[125] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__6_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2002),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[126] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_15__7_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[127] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[8] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[9] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2109),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[10] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__3_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[11] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[12] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2112),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[13] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__6_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[14] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_1__7_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[15] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[16] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[17] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2101),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[18] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[19] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__4_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[20] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__5_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[21] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__6_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[22] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_2__7_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2106),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[23] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__0_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2099),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[24] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__1_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2092),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[25] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__2_ (.CLK(clknet_leaf_1_HCLK),
    .D(n2093),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[26] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__3_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2094),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[27] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2095),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[28] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2096),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[29] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__6_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2097),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[30] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_3__7_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2098),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[31] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__0_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2091),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[32] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__1_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2084),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[33] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__2_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2085),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[34] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2086),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[35] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__4_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2087),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[36] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__5_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2088),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[37] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__6_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2089),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[38] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_4__7_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2090),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[39] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2083),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[40] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2076),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[41] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2077),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[42] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__3_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2078),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[43] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2079),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[44] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2080),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[45] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__6_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2081),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[46] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_5__7_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2082),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[47] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2075),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[48] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2068),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[49] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2069),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[50] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2070),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[51] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__4_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2071),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[52] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__5_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2072),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[53] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__6_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2073),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[54] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_6__7_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2074),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[55] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__0_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2067),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[56] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__1_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2060),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[57] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2061),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[58] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__3_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2062),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[59] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2063),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[60] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2064),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[61] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__6_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2065),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[62] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_7__7_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2066),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[63] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2059),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[64] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__1_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2052),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[65] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__2_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2053),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[66] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2054),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[67] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__4_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2055),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[68] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__5_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2056),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[69] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__6_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2057),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[70] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_8__7_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2058),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[71] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__0_ (.CLK(clknet_leaf_8_HCLK),
    .D(n2051),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[72] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__1_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2044),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[73] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2045),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[74] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__3_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2046),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[75] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__4_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2047),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[76] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__5_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2048),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[77] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__6_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2049),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[78] ));
 sky130_fd_sc_hd__dfxtp_1 inst_to_wrap_tx_fifo_array_reg_reg_9__7_ (.CLK(clknet_leaf_0_HCLK),
    .D(n2050),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_array_reg[79] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_tx_fifo_empty_reg_reg (.CLK(clknet_leaf_5_HCLK),
    .D(n2128),
    .SET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(n_TX_EMPTY_FLAG_FLAG_));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_tx_fifo_full_reg_reg (.CLK(clknet_leaf_7_HCLK),
    .D(n2139),
    .RESET_B(net238),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(n_TX_FULL_FLAG_FLAG_));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_tx_fifo_level_reg_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2137),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\TXFIFOLEVEL_REG[0] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_tx_fifo_level_reg_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2136),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\TXFIFOLEVEL_REG[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_tx_fifo_level_reg_reg_2_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2135),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\TXFIFOLEVEL_REG[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_tx_fifo_level_reg_reg_3_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2134),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\TXFIFOLEVEL_REG[3] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_tx_fifo_r_ptr_reg_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2140),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_r_ptr_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_tx_fifo_r_ptr_reg_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2126),
    .RESET_B(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_r_ptr_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_tx_fifo_r_ptr_reg_reg_2_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2125),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_r_ptr_reg[2] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_tx_fifo_r_ptr_reg_reg_3_ (.CLK(clknet_leaf_5_HCLK),
    .D(n2124),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_r_ptr_reg[3] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_tx_fifo_w_ptr_reg_reg_0_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2132),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_w_ptr_reg[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_tx_fifo_w_ptr_reg_reg_1_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2131),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_w_ptr_reg[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_tx_fifo_w_ptr_reg_reg_2_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2130),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_w_ptr_reg[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_tx_fifo_w_ptr_reg_reg_3_ (.CLK(clknet_leaf_7_HCLK),
    .D(n2129),
    .RESET_B(net242),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_tx_fifo_w_ptr_reg[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_rstn_sq_reg_0_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(net329),
    .RESET_B(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_rstn_sq[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_rstn_sq_reg_1_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(net69),
    .RESET_B(net155),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_rstn_sq[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(net331),
    .RESET_B(net298),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(net70),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2143),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q_reg_1_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2144),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1935),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_10_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1954),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_11_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1964),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_12_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1974),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_13_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1984),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_14_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1994),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_15_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n2151),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_16_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(net142),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_17_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1943),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_18_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1953),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_19_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1963),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_1_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1945),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_20_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1973),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_21_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1983),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_22_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1993),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_23_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n2150),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_24_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1932),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_25_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net125),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_26_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1952),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_27_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1962),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_28_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1972),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_29_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net101),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_2_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net137),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_30_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1992),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_31_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n2149),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_32_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1931),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[32] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_33_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1941),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[33] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_34_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1951),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[34] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_35_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1961),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[35] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_36_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1971),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[36] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_37_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1981),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[37] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_38_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net86),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[38] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_39_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2148),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[39] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_3_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net75),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_40_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1930),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[40] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_41_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1940),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[41] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_42_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1950),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[42] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_43_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1960),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[43] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_44_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1970),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[44] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_45_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1980),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[45] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_46_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(net112),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[46] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_47_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2147),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[47] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_48_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1929),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[48] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_49_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1939),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[49] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_4_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(net80),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_50_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1949),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[50] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_51_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1959),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[51] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_52_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(net77),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[52] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_53_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1979),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[53] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_54_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1989),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[54] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_55_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n2146),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[55] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_56_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1928),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[56] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_57_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1938),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[57] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_58_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1948),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[58] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_59_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(net109),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[59] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_5_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net98),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_60_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1968),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[60] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_61_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1978),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[61] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_62_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1988),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[62] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_63_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n2145),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[63] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_64_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(net139),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[64] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_65_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(net128),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[65] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_66_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(net130),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[66] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_67_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1957),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[67] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_68_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1967),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[68] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_69_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1977),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[69] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_6_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1995),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_70_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1987),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[70] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_71_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(net88),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[71] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_7_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net92),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_8_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1934),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_9_ (.CLK(clknet_leaf_8_usb_cdc_clk_48MHz),
    .D(n1944),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q[9] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_0_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2163),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[0] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_1_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2157),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_2_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2159),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_3_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2161),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q[3] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_0_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2164),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[0] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_1_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2158),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_2_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2160),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_3_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2162),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq[3] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q_reg_0_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2155),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[0] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q_reg_1_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2156),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q_reg_2_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2154),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q_reg_3_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2153),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q[3] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q_reg (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n3841),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_state_q_reg (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2166),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_state_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_valid_q_reg (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1926),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_bulk_in_valid));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1936),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1946),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_2_ (.CLK(clknet_leaf_5_HCLK),
    .D(n1956),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_3_ (.CLK(clknet_leaf_6_HCLK),
    .D(n1966),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[3] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_4_ (.CLK(clknet_leaf_6_HCLK),
    .D(n1976),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[4] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_5_ (.CLK(clknet_leaf_6_HCLK),
    .D(n1986),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[5] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_6_ (.CLK(clknet_leaf_6_HCLK),
    .D(n1996),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[6] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_7_ (.CLK(clknet_leaf_6_HCLK),
    .D(n2248),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_mask_q_reg (.CLK(clknet_leaf_5_HCLK),
    .D(n2141),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_mask_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(net330),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(net347),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_mask_q_reg (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2142),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_mask_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq_reg_0_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(net322),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq_reg_1_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(net356),
    .RESET_B(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1841),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q_reg_1_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1840),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_delay_out_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_0_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1808),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_10_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1818),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_11_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1819),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_12_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1820),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_13_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1821),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_14_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1822),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_15_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1823),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_16_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1824),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_17_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1825),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_18_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1826),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_19_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1827),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_1_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1809),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_20_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1828),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_21_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1829),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_22_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1830),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_23_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1831),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_24_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1832),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_25_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1833),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_26_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1834),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_27_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1835),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_28_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1836),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_29_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1837),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_2_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1810),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_30_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1838),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_31_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1839),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_32_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1776),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[32] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_33_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1777),
    .RESET_B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[33] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_34_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1778),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[34] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_35_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1779),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[35] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_36_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1780),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[36] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_37_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1781),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[37] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_38_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1782),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[38] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_39_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1783),
    .RESET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[39] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_3_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1811),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_40_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1784),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[40] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_41_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1785),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[41] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_42_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1786),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[42] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_43_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1787),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[43] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_44_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1788),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[44] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_45_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1789),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[45] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_46_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1790),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[46] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_47_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1791),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[47] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_48_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1792),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[48] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_49_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1793),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[49] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_4_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1812),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_50_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1794),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[50] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_51_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1795),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[51] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_52_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1796),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[52] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_53_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1797),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[53] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_54_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1798),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[54] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_55_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1799),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[55] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_56_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1800),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[56] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_57_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1801),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[57] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_58_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1802),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[58] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_59_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1803),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[59] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_5_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1813),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_60_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1804),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[60] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_61_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1805),
    .RESET_B(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[61] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_62_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1806),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[62] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_63_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1807),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[63] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_64_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1870),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[64] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_65_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1871),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[65] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_66_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1872),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[66] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_67_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1873),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[67] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_68_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1874),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[68] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_69_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1875),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[69] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_6_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1814),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_70_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1876),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[70] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_71_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1877),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[71] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_7_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1815),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_8_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1816),
    .RESET_B(net201),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_9_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1817),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q[9] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q_reg_0_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1863),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[0] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q_reg_1_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1862),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q_reg_2_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1861),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q_reg_3_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1864),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_first_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_full_q_reg (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1580),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_full_o));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1868),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q_reg_1_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1867),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q_reg_2_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1866),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q_reg_3_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1865),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_q[3] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1881),
    .RESET_B(net198),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq_reg_1_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1880),
    .RESET_B(net197),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq_reg_2_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1879),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq_reg_3_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1878),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_last_qq[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_nak_q_reg (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1869),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_bulk_out_nak));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1883),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q_reg_1_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1882),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_0_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1775),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_1_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1758),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_2_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1741),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_3_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1724),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_4_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1707),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_5_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1690),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_6_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1673),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_7_ (.CLK(clknet_leaf_1_usb_cdc_clk_48MHz),
    .D(n1656),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_out_data_o[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_mask_q_reg (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(n1860),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_mask_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(net316),
    .RESET_B(net191),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq_reg_1_ (.CLK(clknet_leaf_9_usb_cdc_clk_48MHz),
    .D(net341),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_mask_q_reg (.CLK(clknet_leaf_5_HCLK),
    .D(n1859),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_mask_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq_reg_0_ (.CLK(clknet_leaf_5_HCLK),
    .D(net332),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq_reg_1_ (.CLK(clknet_leaf_5_HCLK),
    .D(net360),
    .RESET_B(net307),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q_reg_0_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1905),
    .RESET_B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q_reg_1_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1906),
    .RESET_B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q_reg_2_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1907),
    .RESET_B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q_reg_3_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1901),
    .RESET_B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q_reg_4_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1902),
    .RESET_B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q_reg_5_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1903),
    .RESET_B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q_reg_6_ (.CLK(clknet_leaf_2_usb_cdc_clk_48MHz),
    .D(n1904),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_0_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1890),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_addr[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_1_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1889),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_addr[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_2_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1888),
    .RESET_B(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_addr[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_3_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1887),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_addr[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_4_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1886),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_addr[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_5_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1885),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_addr[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_6_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1884),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_addr[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_0_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1922),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_1_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1921),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_2_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1920),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_3_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1919),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[3] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_4_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1918),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[4] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_5_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1917),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[5] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_6_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n1923),
    .RESET_B(net195),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q_reg (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1915),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q_reg_0_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1909),
    .SET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q_reg_1_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1908),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2229),
    .RESET_B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq_reg_1_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2226),
    .RESET_B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q_reg (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1924),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_endp_q_reg (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1916),
    .RESET_B(net194),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_endp_q));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q_reg (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(inst_to_wrap_u_usb_cdc_ctrl_in_req),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_req_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1895),
    .RESET_B(net186),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_1_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1896),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_2_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1897),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_3_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n2227),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_4_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1900),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_5_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1899),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_6_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1898),
    .RESET_B(net192),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q[6] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q_reg_0_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1913),
    .RESET_B(n3860),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q_reg_1_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1914),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q_reg_0_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1911),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q_reg_1_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1910),
    .RESET_B(net200),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q_reg_2_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n1912),
    .RESET_B(net188),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q_reg_3_ (.CLK(clknet_leaf_0_usb_cdc_clk_48MHz),
    .D(n2228),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1925),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q_reg_1_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2230),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_ctrl_endp_usb_reset_q_reg (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(inst_to_wrap_u_usb_cdc_u_ctrl_endp_N109),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_ctrl_endp_usb_reset_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_0_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2174),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_1_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2175),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_2_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2176),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_3_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2177),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_4_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2178),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_5_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2179),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_6_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2180),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_addr_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2201),
    .RESET_B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_10_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2211),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_11_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2212),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[11] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_12_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2213),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_13_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2214),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_14_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2215),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_15_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2216),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_1_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2202),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_2_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2203),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_3_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2204),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_4_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2205),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_5_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2206),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_6_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2207),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_7_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2208),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_8_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2209),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_9_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2210),
    .RESET_B(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_crc16_q[9] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2185),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[0] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_10_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2195),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_11_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2196),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[3] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_12_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2197),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_13_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2198),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_14_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2199),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[6] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_15_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2200),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[7] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_1_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2186),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_2_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2187),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[2] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_3_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2188),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[3] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_4_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2189),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[4] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_5_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2190),
    .RESET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[5] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_6_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2191),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[6] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_7_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2192),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_data_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_8_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2193),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_9_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2194),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_out_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2217),
    .RESET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q_reg_1_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2218),
    .RESET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2219),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q_reg_1_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2220),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n1894),
    .RESET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_1_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1891),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_2_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1892),
    .RESET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_3_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n1893),
    .RESET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_4_ (.CLK(clknet_leaf_3_usb_cdc_clk_48MHz),
    .D(n2232),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2181),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_endp[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_1_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2182),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_endp[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_2_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2183),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_endp[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_3_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2184),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_endp[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2221),
    .RESET_B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_1_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2222),
    .RESET_B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_2_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2223),
    .RESET_B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_3_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2224),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_in_byte_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_in_data_ack_q_reg (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2165),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_in_data_ack));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_out_eop_q_reg (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2167),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_sie_out_eop_q));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_out_err_q_reg (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2231),
    .RESET_B(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_out_err));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n2225),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_1_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2168),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_2_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2169),
    .RESET_B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_3_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2233),
    .RESET_B(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_phy_state_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2170),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_1_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2171),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_2_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2172),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_3_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2173),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_pid_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n3840),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q_reg_1_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_N51),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_clk_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2269),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_10_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2261),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_11_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2262),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_12_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2263),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_13_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2264),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_14_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2265),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_15_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2266),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_16_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2267),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_17_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2268),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_1_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2252),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_2_ (.CLK(clknet_leaf_7_usb_cdc_clk_48MHz),
    .D(n2253),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_3_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2254),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_4_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2255),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[4] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_5_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2256),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_6_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2257),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_7_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2258),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_8_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2259),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q_reg_9_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2260),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1591),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_0_));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_1_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1592),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_2_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1593),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_3_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1594),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_4_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1595),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_5_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1596),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_6_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1597),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_7_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1598),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[6] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_8_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1578),
    .SET_B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_rx_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[1] ),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q_reg_1_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(net333),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q_reg_2_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(net302),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_pu_q_reg (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2250),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(net57));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[1] ),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q_reg_1_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(net334),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q_reg_2_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(net300),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1601),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q_reg_1_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1602),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q_reg_2_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1603),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q_reg_3_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1604),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_nrzi_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q_reg (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n2251),
    .RESET_B(net228),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q_reg_0_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1589),
    .RESET_B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q_reg_1_ (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1590),
    .RESET_B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q_reg_2_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1599),
    .RESET_B(n3852),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_fq_reg (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1584),
    .RESET_B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_fq));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq_reg (.CLK(clknet_leaf_5_usb_cdc_clk_48MHz),
    .D(n1588),
    .RESET_B(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q_reg_0_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1587),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q_reg_1_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1586),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q_reg_2_ (.CLK(clknet_leaf_6_usb_cdc_clk_48MHz),
    .D(n1585),
    .RESET_B(net229),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_stuffing_cnt_q[2] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2241),
    .SET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[0] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q_reg_1_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2242),
    .SET_B(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[1] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q_reg_2_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2246),
    .SET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_N30),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q_reg_1_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_N31),
    .RESET_B(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2240),
    .RESET_B(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_1_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2239),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_2_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2238),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_3_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2237),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_4_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2236),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_5_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2235),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_6_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2234),
    .RESET_B(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[6] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_7_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2243),
    .SET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q[7] ));
 sky130_fd_sc_hd__dfstp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q_reg (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n1577),
    .SET_B(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n1582),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q_reg_1_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n1581),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q_reg_2_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n1600),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q_reg_0_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2244),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q_reg_1_ (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n2245),
    .RESET_B(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q_reg (.CLK(clknet_leaf_4_usb_cdc_clk_48MHz),
    .D(n1583),
    .RESET_B(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_0_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1624),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[0] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_10_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1634),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[10] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_11_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1635),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[11] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_12_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1636),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[12] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_13_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1637),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[13] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_14_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1638),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[14] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_15_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1639),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[15] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_1_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1625),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[1] ));
 sky130_fd_sc_hd__dfrtp_2 last_HADDR_reg_2_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1626),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[2] ));
 sky130_fd_sc_hd__dfrtp_4 last_HADDR_reg_3_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1627),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[3] ));
 sky130_fd_sc_hd__dfrtp_4 last_HADDR_reg_4_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1628),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[4] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_5_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1629),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[5] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_6_ (.CLK(clknet_leaf_2_HCLK),
    .D(n1630),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[6] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_7_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1631),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[7] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_8_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1632),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[8] ));
 sky130_fd_sc_hd__dfrtp_1 last_HADDR_reg_9_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1633),
    .RESET_B(net240),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(\last_HADDR[9] ));
 sky130_fd_sc_hd__dfrtp_1 last_HSEL_reg (.CLK(clknet_leaf_1_HCLK),
    .D(n1621),
    .RESET_B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(last_HSEL));
 sky130_fd_sc_hd__dfrtp_1 last_HTRANS_reg_1_ (.CLK(clknet_leaf_1_HCLK),
    .D(n1622),
    .RESET_B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(last_HTRANS_1_));
 sky130_fd_sc_hd__dfrtp_1 last_HWRITE_reg (.CLK(clknet_leaf_1_HCLK),
    .D(n1623),
    .RESET_B(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .Q(last_HWRITE));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_84 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_88 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_89 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_112 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_115 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_140 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_143 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_151 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_166 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_167 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_168 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_169 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_170 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_171 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_172 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_173 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_174 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_175 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_176 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_177 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_178 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_179 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_180 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_181 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_182 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_183 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_184 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_185 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_186 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_187 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_188 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_189 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_190 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_191 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_192 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_193 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_194 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_195 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_196 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_197 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_198 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_199 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_200 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_201 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_202 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_203 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_204 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_205 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_206 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_207 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_208 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_209 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_210 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_211 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_212 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_213 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_214 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_215 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_216 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_217 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_218 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_219 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_220 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_221 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_222 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_223 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_224 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_225 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_226 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_227 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_228 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_229 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_230 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_231 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_232 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_233 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_234 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_235 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_236 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_237 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_238 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_239 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_240 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_241 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_242 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_243 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_244 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_245 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_246 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_247 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_248 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_249 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_250 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_251 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_252 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_253 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_254 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_255 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_256 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_257 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_258 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_259 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_260 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_261 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_262 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_263 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_264 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_265 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_266 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_267 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_268 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_269 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_270 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_271 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_272 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_273 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_274 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_275 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_276 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_277 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_278 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_279 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_280 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_281 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_282 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_283 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_284 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_285 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_286 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_287 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_288 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_289 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_290 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_291 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_292 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_293 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_294 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_295 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_296 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_297 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_298 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_299 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_300 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_301 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_302 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_303 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_304 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_305 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_306 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_307 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_308 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_309 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_310 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_311 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_312 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_313 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_314 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_315 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_316 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_317 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_318 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_319 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_320 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_321 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_322 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_323 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_324 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_325 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_326 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_327 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_328 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_329 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_330 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_331 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_332 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_333 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_334 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_335 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_336 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_337 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_338 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_339 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_340 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_341 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_342 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_343 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_344 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_345 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_346 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_347 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_348 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_349 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_350 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_351 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_352 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_353 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_354 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_355 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_356 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_357 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_358 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_359 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_360 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_361 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_362 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_363 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_364 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_365 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_366 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_367 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_368 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_369 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_370 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_371 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_372 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_373 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_374 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_375 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_376 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_377 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_378 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_379 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_380 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_381 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_382 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_383 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_384 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_385 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_386 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_387 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_388 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_389 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_390 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_391 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_392 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_393 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_394 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_395 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_396 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_397 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_398 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_399 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_400 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_401 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_402 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_403 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_404 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_405 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_406 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_407 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_408 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_409 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_410 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_411 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_412 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_413 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_414 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_415 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_416 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_417 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_418 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_419 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_420 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_421 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_422 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_423 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_424 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_425 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_426 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_427 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_428 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_429 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_430 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_431 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_432 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_433 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_434 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_435 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_436 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_437 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_438 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_439 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_440 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_441 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_442 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_443 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_444 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_445 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_446 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_447 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_448 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_449 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_450 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_451 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_452 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_453 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_454 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_455 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_456 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_457 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_458 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_459 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_460 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_461 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_462 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_463 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_464 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_465 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_466 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_467 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_468 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_469 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_470 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_471 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_472 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_473 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_474 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_475 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_476 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_477 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_478 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_479 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_480 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_481 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_482 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_483 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_484 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_485 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_486 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_487 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_488 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_489 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_490 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_491 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_492 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_493 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_494 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_495 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_496 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_497 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_498 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_499 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_500 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_501 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_502 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_503 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_504 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_505 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_506 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_507 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_508 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_509 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_510 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_511 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_512 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_513 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_514 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_515 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_516 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_517 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_518 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_519 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_520 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_521 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_522 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_523 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_524 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_525 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_526 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_527 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_528 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_529 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_530 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_531 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_532 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_533 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_534 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_535 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_536 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_537 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_538 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_539 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_540 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_541 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_542 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_543 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_544 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_545 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_546 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_547 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_548 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_549 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_550 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_551 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_552 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_553 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_554 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_555 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_556 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_557 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_558 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_559 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_560 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_561 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_562 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_563 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_564 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_565 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_566 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_567 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_568 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_569 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_570 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_571 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_572 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_573 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_574 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_575 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_576 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_577 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_578 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_579 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_580 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_581 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_582 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_583 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_584 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_585 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_586 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_587 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_588 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_589 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_590 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_591 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_592 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_593 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_594 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_595 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_596 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_597 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_598 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_599 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_600 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_601 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_602 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_603 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_604 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_605 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_606 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_607 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_608 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_609 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_610 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_611 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_612 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_613 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_614 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_615 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_616 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_617 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_618 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_619 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_620 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_621 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_622 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_623 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_624 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_625 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_626 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_627 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_628 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_629 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_630 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_631 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_632 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_633 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_634 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_635 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_636 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_637 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_638 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_639 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_640 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_641 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_642 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_643 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_644 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_645 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_646 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_647 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_648 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_649 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_650 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_651 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_652 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_653 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_654 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_655 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_656 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_657 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_658 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_659 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_660 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_661 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_662 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_663 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_664 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_665 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_666 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_667 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_668 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_669 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_670 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_671 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_672 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_673 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_674 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_675 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_676 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_677 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_678 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_679 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_680 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_681 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_682 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_683 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_684 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_685 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_686 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_687 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_688 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_689 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_690 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_691 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_692 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_693 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_694 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_695 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_696 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_697 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_698 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_699 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_700 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_701 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_702 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_703 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_704 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_705 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_706 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_707 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_708 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_709 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_710 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_711 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_712 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_713 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_714 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_715 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_716 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_717 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_718 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_719 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_720 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_721 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_722 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_723 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_724 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_725 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_726 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_727 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_728 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_729 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_730 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_731 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_732 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_733 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_734 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_735 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_736 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_737 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_738 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_739 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_740 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_741 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_742 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_743 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_744 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_745 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_746 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_747 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_748 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_749 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_750 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_751 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_752 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_753 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_754 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_755 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_756 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_757 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_758 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_759 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_760 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_761 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_762 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_763 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_764 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_765 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_766 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_767 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_768 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_769 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_770 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_771 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_772 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_773 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_774 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_775 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_776 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_777 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_778 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_779 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_780 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_781 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_782 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_783 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_784 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_785 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_786 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_787 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_788 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_789 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_790 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_791 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_792 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_793 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_794 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_795 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_796 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_797 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_798 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_799 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_800 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_801 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_802 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_803 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_804 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_805 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_806 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_807 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_808 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_809 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_810 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_811 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_812 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_813 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_814 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_815 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_816 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_817 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_818 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_819 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_820 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_821 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_822 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_823 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_824 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_825 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_826 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_827 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_828 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_829 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_830 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_831 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_832 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_833 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_834 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_835 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_836 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_837 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_838 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_839 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_840 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_841 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_842 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_843 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_844 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_845 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_846 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_847 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_848 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_849 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_850 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_851 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_852 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_853 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_854 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_855 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_856 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_857 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_858 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_859 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_860 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_861 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_862 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_863 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_864 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_865 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_866 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_867 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_868 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_869 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_870 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_871 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_872 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_873 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_874 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_875 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_876 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_877 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_878 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_879 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_880 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_881 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_882 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_883 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_884 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_885 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_886 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_887 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_888 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_889 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_890 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_891 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_892 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_893 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_894 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_895 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_896 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_897 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_898 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_899 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_900 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_901 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_902 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_903 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_904 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_905 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_906 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_907 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_908 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_909 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_910 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_911 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_912 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_913 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_914 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_915 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_916 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_917 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_918 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_919 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_920 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_921 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_922 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_923 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_924 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_925 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_926 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_927 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_928 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_929 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_930 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_931 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_932 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_933 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_934 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_935 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_936 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_937 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_938 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_939 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_940 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_941 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_942 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_943 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_944 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_945 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_946 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_947 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_948 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_949 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_950 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_951 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_952 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_953 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_954 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_955 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_956 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_957 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_958 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_959 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_960 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_961 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_962 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_963 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_964 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_965 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_966 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_967 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_968 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_969 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_970 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_971 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_972 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_973 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_974 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_975 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_976 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_977 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_978 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_979 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_980 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_981 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_982 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_983 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_984 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_985 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_986 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_987 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_988 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_989 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_990 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_991 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_992 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_993 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_994 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_995 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_996 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_997 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_998 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_999 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1000 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1001 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1002 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1003 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1004 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1005 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1006 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1007 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1008 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_1009 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1010 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1011 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1012 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1013 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1014 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1015 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1016 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1017 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1018 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1019 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1020 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1021 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_1022 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1023 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1024 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1025 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1026 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1027 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1028 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1029 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1030 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1031 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1032 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1033 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1034 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1035 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1036 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1037 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1038 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1039 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1040 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1041 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1042 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1043 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1044 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1045 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1046 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1047 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1048 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1049 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1050 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1051 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1052 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1053 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1054 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1055 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1056 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1057 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1058 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1059 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1060 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1061 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1062 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1063 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1064 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1065 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1066 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1067 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1068 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1069 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1070 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1071 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1072 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1073 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1074 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1075 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1076 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1077 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1078 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1079 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1080 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1081 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1082 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1083 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1084 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1085 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1086 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1087 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1088 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1089 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1090 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1091 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1092 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1093 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1094 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1095 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1096 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1097 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1098 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1099 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1100 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1101 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1102 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1103 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1104 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1105 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1106 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1107 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1108 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1109 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1110 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1111 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1112 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1113 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1114 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1115 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1116 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1117 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1118 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1119 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1120 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1121 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1122 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1123 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1124 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1125 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1126 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1127 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1128 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1129 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1130 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1131 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1132 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1133 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1134 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1135 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1136 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1137 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1138 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1139 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1140 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1141 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1142 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1143 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1144 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1145 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1146 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1147 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1148 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1149 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1150 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1151 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1152 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1153 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1154 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1155 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1156 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1157 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1158 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1159 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1160 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1161 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1162 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1163 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1164 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1165 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__buf_4 fanout184 (.A(n2866),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net184));
 sky130_fd_sc_hd__buf_4 fanout185 (.A(n3029),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net185));
 sky130_fd_sc_hd__clkbuf_8 fanout186 (.A(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net186));
 sky130_fd_sc_hd__buf_6 fanout187 (.A(n3862),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_8 fanout188 (.A(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net188));
 sky130_fd_sc_hd__clkbuf_8 fanout189 (.A(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net189));
 sky130_fd_sc_hd__buf_4 fanout190 (.A(n3863),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_8 fanout191 (.A(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 fanout192 (.A(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net192));
 sky130_fd_sc_hd__clkbuf_8 fanout193 (.A(n3866),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_8 fanout194 (.A(net196),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_8 fanout195 (.A(n3865),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net195));
 sky130_fd_sc_hd__buf_2 fanout196 (.A(n3865),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_8 fanout197 (.A(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_8 fanout198 (.A(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net198));
 sky130_fd_sc_hd__buf_4 fanout199 (.A(n3867),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_8 fanout200 (.A(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_4 fanout201 (.A(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net201));
 sky130_fd_sc_hd__clkbuf_8 fanout202 (.A(n3868),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_8 fanout203 (.A(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_8 fanout204 (.A(net296),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_8 fanout205 (.A(net295),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net205));
 sky130_fd_sc_hd__buf_4 fanout206 (.A(n3289),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(n2481),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net207));
 sky130_fd_sc_hd__buf_6 fanout208 (.A(net305),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net208));
 sky130_fd_sc_hd__buf_4 fanout209 (.A(n3301),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net209));
 sky130_fd_sc_hd__buf_4 fanout210 (.A(\inst_to_wrap_u_usb_cdc_out_data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_4 fanout211 (.A(\inst_to_wrap_u_usb_cdc_out_data[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_8 fanout212 (.A(\inst_to_wrap_u_usb_cdc_out_data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net212));
 sky130_fd_sc_hd__buf_2 fanout213 (.A(\inst_to_wrap_u_usb_cdc_out_data[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net213));
 sky130_fd_sc_hd__buf_4 fanout214 (.A(\inst_to_wrap_u_usb_cdc_out_data[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net214));
 sky130_fd_sc_hd__buf_4 fanout215 (.A(\inst_to_wrap_u_usb_cdc_out_data[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_8 fanout216 (.A(\inst_to_wrap_u_usb_cdc_out_data[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net216));
 sky130_fd_sc_hd__clkbuf_8 fanout217 (.A(\inst_to_wrap_u_usb_cdc_out_data[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_8 fanout218 (.A(\inst_to_wrap_u_usb_cdc_out_data[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_8 fanout219 (.A(\inst_to_wrap_u_usb_cdc_out_data[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net219));
 sky130_fd_sc_hd__buf_4 fanout220 (.A(net245),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net220));
 sky130_fd_sc_hd__clkbuf_8 fanout221 (.A(net177),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net221));
 sky130_fd_sc_hd__buf_4 fanout222 (.A(net274),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net222));
 sky130_fd_sc_hd__buf_4 fanout223 (.A(net256),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net223));
 sky130_fd_sc_hd__buf_4 fanout224 (.A(net287),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net224));
 sky130_fd_sc_hd__buf_4 fanout225 (.A(net260),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net225));
 sky130_fd_sc_hd__buf_4 fanout226 (.A(net270),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net226));
 sky130_fd_sc_hd__buf_4 fanout227 (.A(net252),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_8 fanout228 (.A(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_8 fanout229 (.A(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net229));
 sky130_fd_sc_hd__buf_4 fanout230 (.A(net306),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(n3699),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net231));
 sky130_fd_sc_hd__buf_4 fanout232 (.A(net25),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net232));
 sky130_fd_sc_hd__buf_4 fanout233 (.A(net24),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net233));
 sky130_fd_sc_hd__buf_4 fanout234 (.A(net23),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net234));
 sky130_fd_sc_hd__buf_4 fanout235 (.A(net22),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net235));
 sky130_fd_sc_hd__buf_4 fanout236 (.A(net21),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net236));
 sky130_fd_sc_hd__buf_4 fanout237 (.A(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net237));
 sky130_fd_sc_hd__buf_4 fanout238 (.A(net239),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net238));
 sky130_fd_sc_hd__buf_2 fanout239 (.A(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net239));
 sky130_fd_sc_hd__buf_4 fanout240 (.A(net241),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net240));
 sky130_fd_sc_hd__buf_2 fanout241 (.A(net154),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net241));
 sky130_fd_sc_hd__buf_4 fanout242 (.A(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net242));
 sky130_fd_sc_hd__buf_6 fanout243 (.A(net157),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_4 fanout244 (.A(net17),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net244));
 sky130_fd_sc_hd__buf_1 input1 (.A(net321),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input2 (.A(net317),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(net312),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(net311),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(net308),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(net309),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(net310),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net7));
 sky130_fd_sc_hd__buf_1 input8 (.A(net325),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(net328),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net9));
 sky130_fd_sc_hd__buf_1 input10 (.A(net327),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net10));
 sky130_fd_sc_hd__buf_1 input11 (.A(net323),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net11));
 sky130_fd_sc_hd__buf_1 input12 (.A(net319),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net12));
 sky130_fd_sc_hd__buf_1 input13 (.A(net324),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net13));
 sky130_fd_sc_hd__buf_1 input14 (.A(net320),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(net313),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(net314),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(HREADY),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input18 (.A(net315),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net18));
 sky130_fd_sc_hd__buf_1 input19 (.A(net318),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(HWDATA[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(HWDATA[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(HWDATA[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(net335),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net23));
 sky130_fd_sc_hd__buf_1 input24 (.A(HWDATA[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net24));
 sky130_fd_sc_hd__buf_1 input25 (.A(HWDATA[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net25));
 sky130_fd_sc_hd__buf_4 input26 (.A(HWDATA[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net26));
 sky130_fd_sc_hd__buf_4 input27 (.A(HWDATA[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(net326),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(net351),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(net349),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_8 output31 (.A(net31),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[0]));
 sky130_fd_sc_hd__clkbuf_8 output32 (.A(net32),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[10]));
 sky130_fd_sc_hd__clkbuf_8 output33 (.A(net33),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[11]));
 sky130_fd_sc_hd__clkbuf_8 output34 (.A(net34),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[12]));
 sky130_fd_sc_hd__clkbuf_8 output35 (.A(net35),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[13]));
 sky130_fd_sc_hd__clkbuf_8 output36 (.A(net36),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[15]));
 sky130_fd_sc_hd__clkbuf_8 output37 (.A(net37),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[16]));
 sky130_fd_sc_hd__clkbuf_8 output38 (.A(net38),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[18]));
 sky130_fd_sc_hd__clkbuf_8 output39 (.A(net39),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[19]));
 sky130_fd_sc_hd__clkbuf_8 output40 (.A(net40),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[1]));
 sky130_fd_sc_hd__clkbuf_8 output41 (.A(net41),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[21]));
 sky130_fd_sc_hd__clkbuf_8 output42 (.A(net42),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[23]));
 sky130_fd_sc_hd__clkbuf_8 output43 (.A(net43),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[25]));
 sky130_fd_sc_hd__clkbuf_8 output44 (.A(net44),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[26]));
 sky130_fd_sc_hd__clkbuf_8 output45 (.A(net45),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[27]));
 sky130_fd_sc_hd__clkbuf_8 output46 (.A(net46),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[28]));
 sky130_fd_sc_hd__clkbuf_8 output47 (.A(net47),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[2]));
 sky130_fd_sc_hd__clkbuf_8 output48 (.A(net48),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[30]));
 sky130_fd_sc_hd__clkbuf_8 output49 (.A(net49),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[31]));
 sky130_fd_sc_hd__clkbuf_8 output50 (.A(net50),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[3]));
 sky130_fd_sc_hd__clkbuf_8 output51 (.A(net51),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[4]));
 sky130_fd_sc_hd__clkbuf_8 output52 (.A(net52),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[5]));
 sky130_fd_sc_hd__clkbuf_8 output53 (.A(net53),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[6]));
 sky130_fd_sc_hd__clkbuf_8 output54 (.A(net54),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[7]));
 sky130_fd_sc_hd__clkbuf_8 output55 (.A(net55),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(HRDATA[9]));
 sky130_fd_sc_hd__clkbuf_8 output56 (.A(net56),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(dn_tx_o));
 sky130_fd_sc_hd__clkbuf_8 output57 (.A(net57),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(dp_pu_o));
 sky130_fd_sc_hd__clkbuf_8 output58 (.A(net58),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(dp_tx_o));
 sky130_fd_sc_hd__clkbuf_8 output59 (.A(net59),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(irq));
 sky130_fd_sc_hd__clkbuf_8 output60 (.A(net60),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(tx_en_o));
 sky130_fd_sc_hd__conb_1 U2292_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .LO(net61));
 sky130_fd_sc_hd__conb_1 U2293_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net62));
 sky130_fd_sc_hd__conb_1 U2294_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net63));
 sky130_fd_sc_hd__conb_1 U2295_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net64));
 sky130_fd_sc_hd__conb_1 U2296_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net65));
 sky130_fd_sc_hd__conb_1 U2297_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net66));
 sky130_fd_sc_hd__conb_1 U2298_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net67));
 sky130_fd_sc_hd__conb_1 U2299_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net68));
 sky130_fd_sc_hd__conb_1 inst_to_wrap_u_usb_cdc_rstn_sq_reg_1__69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net69));
 sky130_fd_sc_hd__conb_1 inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq_reg_1__70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(net70));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_HCLK (.A(clknet_1_1__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_HCLK (.A(clknet_1_1__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_HCLK (.A(clknet_1_1__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_HCLK (.A(clknet_1_1__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_HCLK (.A(clknet_1_1__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_HCLK (.A(clknet_1_0__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_HCLK (.A(clknet_1_0__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_HCLK (.A(clknet_1_0__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_HCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_HCLK (.A(HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_HCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_HCLK (.A(clknet_0_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_HCLK));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_HCLK (.A(clknet_0_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_HCLK));
 sky130_fd_sc_hd__clkbuf_8 clkload0 (.A(clknet_1_0__leaf_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload1 (.A(clknet_leaf_0_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload2 (.A(clknet_leaf_7_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_8 clkload3 (.A(clknet_leaf_8_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(clknet_leaf_1_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload5 (.A(clknet_leaf_2_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload6 (.A(clknet_leaf_3_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkload7 (.A(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_0_usb_cdc_clk_48MHz (.A(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_0_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_1_usb_cdc_clk_48MHz (.A(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_1_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_2_usb_cdc_clk_48MHz (.A(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_2_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_3_usb_cdc_clk_48MHz (.A(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_3_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_4_usb_cdc_clk_48MHz (.A(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_4_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_5_usb_cdc_clk_48MHz (.A(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_5_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_6_usb_cdc_clk_48MHz (.A(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_6_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_7_usb_cdc_clk_48MHz (.A(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_7_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_8_usb_cdc_clk_48MHz (.A(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_8_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_leaf_9_usb_cdc_clk_48MHz (.A(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_leaf_9_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_usb_cdc_clk_48MHz (.A(usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_0_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_usb_cdc_clk_48MHz (.A(clknet_0_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_0__leaf_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_usb_cdc_clk_48MHz (.A(clknet_0_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(clknet_1_1__leaf_usb_cdc_clk_48MHz));
 sky130_fd_sc_hd__clkbuf_4 clkload8 (.A(clknet_leaf_0_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload9 (.A(clknet_leaf_1_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkinv_16 clkload10 (.A(clknet_leaf_9_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload11 (.A(clknet_leaf_3_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload12 (.A(clknet_leaf_4_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload13 (.A(clknet_leaf_5_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__clkbuf_4 clkload14 (.A(clknet_leaf_7_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(net354),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net362),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net340),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net114),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(n1965),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net82),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(n1969),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net81),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(net83),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(n1975),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net89),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(net78),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net76),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net79),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(net118),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(n1991),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net94),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(n2247),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net93),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(net95),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(n2152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net102),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(net90),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net87),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net91),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(net104),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(n1985),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net103),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(net105),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(n1982),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(net121),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net99),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net97),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(net100),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net113),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net115),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(n1958),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net117),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net119),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(n1990),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net122),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net107),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(net74),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net108),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net123),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(net110),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net85),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net111),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(net132),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(n1942),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net131),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(net133),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(n1937),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net144),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(n1947),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net152),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net126),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(net124),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net127),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net143),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(net145),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(n1955),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net148),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(n1927),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net147),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net149),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(n1933),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(net352),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(net135),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net129),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net136),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(net151),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(net140),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net138),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net141),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net358),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net156),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(net243),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(HRESETn),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net154),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net291),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(n1723),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net281),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(n1757),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(net284),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(n1740),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net344),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(net346),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(net264),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(n1706),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net249),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(n1655),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net278),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(n1689),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(net267),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(n1774),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net181),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(n1672),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net180),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net182),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net177));
 sky130_fd_sc_hd__buf_4 hold108 (.A(net221),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(n1660),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\inst_to_wrap_out_data_o[6] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net176),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(net174),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net248),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net250),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net245));
 sky130_fd_sc_hd__buf_4 hold115 (.A(net220),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(n1643),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\inst_to_wrap_out_data_o[7] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(net183),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(net168),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(net266),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(net268),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net252));
 sky130_fd_sc_hd__buf_4 hold122 (.A(net227),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(n1768),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(net263),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(net265),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net256));
 sky130_fd_sc_hd__buf_4 hold126 (.A(net223),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(n1700),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(net283),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(net285),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net260));
 sky130_fd_sc_hd__buf_4 hold130 (.A(net225),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(n1728),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\inst_to_wrap_out_data_o[4] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(net255),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(net166),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\inst_to_wrap_out_data_o[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(net251),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(net172),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(net280),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(net282),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net270));
 sky130_fd_sc_hd__buf_4 hold140 (.A(net226),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(n1745),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(net277),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(net279),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net274));
 sky130_fd_sc_hd__buf_4 hold144 (.A(net222),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(n1681),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\inst_to_wrap_out_data_o[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(net273),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(net170),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\inst_to_wrap_out_data_o[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(net269),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(net160),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\inst_to_wrap_out_data_o[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(net259),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(net162),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(net290),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(net292),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net287));
 sky130_fd_sc_hd__buf_4 hold157 (.A(net224),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(n1716),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\inst_to_wrap_out_data_o[3] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(net286),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(net158),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_cnt_q[5] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(net304),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(n3864),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(net204),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(net348),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(net30),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(net350),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(net29),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_en_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(n1576),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(net294),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\inst_to_wrap_u_usb_cdc_rstn_sq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net306));
 sky130_fd_sc_hd__buf_4 hold176 (.A(net364),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(HADDR[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(HADDR[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(HADDR[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(HADDR[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(HADDR[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(HADDR[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(HADDR[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(HSEL),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_sq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(HADDR[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(HTRANS[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(HADDR[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(HADDR[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(HADDR[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(HADDR[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(HADDR[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(HADDR[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(HWRITE),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(HADDR[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(HADDR[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\inst_to_wrap_u_usb_cdc_rstn_sq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq[1] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dn_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_dp_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(HWDATA[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(net353),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(net355),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(net361),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(net72),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(n3838),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(net73),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(net357),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(net359),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_mask_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(net164),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(n3839),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(net165),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(dp_rx_i),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(net299),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(dn_rx_i),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(net301),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q[2] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(net363),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(net336),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(net71),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(net337),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_iready_mask_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(net342),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(net153),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(net343),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_mask_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(net338),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_mask_q),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold190_A (.DIODE(HADDR[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold186_A (.DIODE(HADDR[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold181_A (.DIODE(HADDR[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold180_A (.DIODE(HADDR[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold177_A (.DIODE(HADDR[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold178_A (.DIODE(HADDR[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold179_A (.DIODE(HADDR[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold194_A (.DIODE(HADDR[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold197_A (.DIODE(HADDR[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold196_A (.DIODE(HADDR[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold192_A (.DIODE(HADDR[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold188_A (.DIODE(HADDR[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold193_A (.DIODE(HADDR[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold189_A (.DIODE(HADDR[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold182_A (.DIODE(HADDR[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold183_A (.DIODE(HADDR[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_HCLK_A (.DIODE(HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_eco_cell_13_0_X (.DIODE(HRDATA[14]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_eco_cell_16_0_X (.DIODE(HRDATA[17]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_eco_cell_19_0_X (.DIODE(HRDATA[20]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_eco_cell_21_0_X (.DIODE(HRDATA[22]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_eco_cell_23_0_X (.DIODE(HRDATA[24]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_eco_cell_28_0_X (.DIODE(HRDATA[29]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_eco_cell_7_0_X (.DIODE(HRDATA[8]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(HREADY),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2292_Y (.DIODE(HREADYOUT),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold86_A (.DIODE(HRESETn),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold184_A (.DIODE(HSEL),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold187_A (.DIODE(HTRANS[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(HWDATA[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(HWDATA[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(HWDATA[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold204_A (.DIODE(HWDATA[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(HWDATA[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(HWDATA[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(HWDATA[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(HWDATA[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold195_A (.DIODE(HWRITE),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold219_A (.DIODE(dn_rx_i),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold217_A (.DIODE(dp_rx_i),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_usb_cdc_clk_48MHz_A (.DIODE(usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_X (.DIODE(HRDATA[0]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_X (.DIODE(HRDATA[10]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_X (.DIODE(HRDATA[11]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_X (.DIODE(HRDATA[12]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_X (.DIODE(HRDATA[13]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_X (.DIODE(HRDATA[15]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_X (.DIODE(HRDATA[16]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_X (.DIODE(HRDATA[18]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_X (.DIODE(HRDATA[19]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_X (.DIODE(HRDATA[1]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output41_X (.DIODE(HRDATA[21]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output42_X (.DIODE(HRDATA[23]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output43_X (.DIODE(HRDATA[25]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output44_X (.DIODE(HRDATA[26]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output45_X (.DIODE(HRDATA[27]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output46_X (.DIODE(HRDATA[28]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output47_X (.DIODE(HRDATA[2]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_X (.DIODE(HRDATA[30]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output49_X (.DIODE(HRDATA[31]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output50_X (.DIODE(HRDATA[3]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output51_X (.DIODE(HRDATA[4]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output52_X (.DIODE(HRDATA[5]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output53_X (.DIODE(HRDATA[6]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output54_X (.DIODE(HRDATA[7]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output55_X (.DIODE(HRDATA[9]),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output56_X (.DIODE(dn_tx_o),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output57_X (.DIODE(dp_pu_o),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output58_X (.DIODE(dp_tx_o),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output59_X (.DIODE(irq),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_X (.DIODE(tx_en_o),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q_reg_1__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_2__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_1__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_0__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q_reg_1__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_dataout_toggle_q_reg_0__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_8__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_7__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_2__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_1__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_15__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_10__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_in_dir_q_reg_RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_5__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_4__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_64__RESET_B (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2560_X (.DIODE(n3859),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2557_X (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold167_A (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_valid_q_reg_RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q_reg_2__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q_reg_1__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_stuffing_cnt_q_reg_0__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_out_eop_q_reg_RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_7__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_10__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_data_q_reg_0__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_state_q_reg_0__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_full_q_reg_RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_71__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_70__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_66__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_32__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_63__RESET_B (.DIODE(n3861),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_X (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_addr_qq_reg_6__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_2__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_5__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_0__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_in_data_ack_q_reg_RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_1__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_pid_q_reg_3__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_1__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_2__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_3__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_4__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_5__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_6__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_0__RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_nak_q_reg_RESET_B (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net187),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_X (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_3__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_3__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_0__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q_reg_0__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_1__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_11__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_12__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_15__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_3__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_4__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_3__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_3__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_14__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_4__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_1__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_2__RESET_B (.DIODE(net189),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_X (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_phy_state_q_reg_2__RESET_B (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_0__RESET_B (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_1__RESET_B (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_0__RESET_B (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_0__RESET_B (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_in_byte_q_reg_2__RESET_B (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_33__RESET_B (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout188_A (.DIODE(net190),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_X (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_1__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_2__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_3__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_req_q_reg_RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_0__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_0__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_1__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_6__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_8__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_9__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_0__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_1__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_endp_q_reg_2__RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_out_err_q_reg_RESET_B (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net193),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout199_X (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_q_reg_0__SET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q_reg_0__RESET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_datain_toggle_q_reg_1__RESET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_0__RESET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_2__RESET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_delay_cnt_q_reg_3__RESET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q_reg_1__SET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_out_fifo_q_reg_39__RESET_B (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout202_X (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_14__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_13__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_12__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_11__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_6__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_valid_q_reg_RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_9__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_6__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_5__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_4__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_crc16_q_reg_3__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_4__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_addr_q_reg_5__RESET_B (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net202),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_X (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_56__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2561_A (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_65__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_66__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_67__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_68__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_69__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_70__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_fifo_q_reg_71__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq_reg_1__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_sq_reg_0__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q_reg_0__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_last_q_reg_3__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_ovalid_mask_q_reg_RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q_reg_1__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_delay_in_cnt_q_reg_0__RESET_B (.DIODE(net203),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_X (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold165_A (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_state_q_reg_RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q_reg_0__SET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_clk_cnt_q_reg_0__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q_reg_0__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_tx_state_q_reg_1__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_qq_reg_0__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_3__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_2__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_1__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_in_first_q_reg_0__RESET_B (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(net205),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_X (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_nrzi_q_reg_SET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_bit_cnt_q_reg_2__SET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_tx_data_q_reg_7__SET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_5__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_2__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2558_A (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2560_A (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2564_A (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_byte_cnt_q_reg_4__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_class_q_reg_RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_1__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_max_length_q_reg_5__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_rec_q_reg_1__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_req_q_reg_3__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_state_q_reg_1__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_data_q_reg_13__RESET_B (.DIODE(net208),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout210_X (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3100_B1 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3106_A1 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3234_A1 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3930_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4190_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3400_A1 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3892_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3940_B1 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4000_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4118_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4128_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4138_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4148_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4159_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4170_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4180_A2 (.DIODE(net210),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_X (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3105_A1 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3235_A1 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3401_A1 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3908_B1 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3931_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4191_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3893_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3941_B1 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4001_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4119_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4129_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4139_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4149_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4160_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4171_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4181_A2 (.DIODE(net212),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_X (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3394_B1 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3927_C (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3907_A (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3890_A1 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3056_A (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3120_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3875_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4132_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4122_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4112_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3994_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4142_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4184_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4174_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4164_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4153_A2 (.DIODE(net214),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_X (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2960_A (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2962_A1 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2979_B2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3056_D (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3083_B (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3395_A1 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3229_A1 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4113_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4123_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4133_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4143_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4154_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4165_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4175_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3938_B1 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3995_A2 (.DIODE(net215),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout216_X (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2966_A (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2991_A (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3230_A1 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4186_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3396_A1 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3056_B (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3996_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4114_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4124_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4134_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4144_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4155_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4166_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4176_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3937_B1 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3891_A2 (.DIODE(net216),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout217_X (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2952_A (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2990_B (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3083_A (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4187_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3397_A1 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3231_A1 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3056_C (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3997_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4115_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4125_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4135_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4145_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4156_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4167_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4177_A2 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3936_B1 (.DIODE(net217),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_X (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2963_B2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3232_A1 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3398_A1 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2989_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2958_A (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3096_A (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3998_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4116_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4126_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4136_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4146_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4157_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4168_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4178_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4188_A2 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3124_A1 (.DIODE(net218),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_X (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_data_q_reg_8__SET_B (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_rq_reg_RESET_B (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_valid_fq_reg_RESET_B (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q_reg_1__RESET_B (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_sie_u_phy_rx_rx_state_q_reg_0__RESET_B (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq_reg_1__RESET_B (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_ctrl_endp_dev_state_qq_reg_0__RESET_B (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout228_A (.DIODE(net230),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_X (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3647_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3687_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4460_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2774_B_N (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3626_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3584_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3551_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3573_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3595_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3616_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3637_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3657_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3667_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3677_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3704_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3697_A2 (.DIODE(net232),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_X (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3648_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3688_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4461_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2773_B_N (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3627_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3585_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3552_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3574_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3596_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3617_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3638_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3658_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3668_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3678_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3705_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3698_A2 (.DIODE(net233),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout234_X (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4462_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4452_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3553_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3564_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3575_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3597_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3607_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3618_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3639_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3649_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3659_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3669_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3679_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3689_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3699_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3706_A2 (.DIODE(net234),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_X (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3630_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3588_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4464_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4454_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3555_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3577_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3599_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3620_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3641_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3651_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3661_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3671_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3681_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3691_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3701_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3708_A2 (.DIODE(net236),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_X (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4467_A0 (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4465_A2 (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4457_A1 (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U4455_A2 (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3623_A2 (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3581_A2 (.DIODE(net20),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_X (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3703_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3696_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3686_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3676_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3666_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3656_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3646_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3636_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3625_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3615_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3604_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3594_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3583_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3572_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3561_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3550_A2 (.DIODE(net26),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_X (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3695_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3685_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3675_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3665_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3655_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3645_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3635_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3624_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3614_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3603_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3593_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3582_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3571_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3560_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U3549_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_U2853_A2 (.DIODE(net27),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkload7_A (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_sq_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_level_reg_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_mask_q_reg_CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_r_ptr_reg_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_r_ptr_reg_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_r_ptr_reg_reg_3__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_iready_sq_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_2__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_in_fifo_u_ltx4_async_data_in_data_q_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_r_ptr_reg_reg_2__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_empty_reg_reg_CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_level_reg_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_u_usb_cdc_u_bulk_endp_u_out_fifo_u_ltx4_async_data_out_ovalid_mask_q_reg_CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_RXFIFOT_REG_reg_2__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_RXFIFOT_REG_reg_3__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_level_reg_reg_3__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_tx_fifo_level_reg_reg_2__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_RIS_REG_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_RXFIFOT_REG_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_RIS_REG_reg_3__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_RXFIFOT_REG_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_level_reg_reg_2__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_level_reg_reg_0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_level_reg_reg_1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_level_reg_reg_3__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_15__1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_15__3__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_13__0__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_13__4__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_13__3__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_13__5__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_13__1__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_inst_to_wrap_rx_fifo_array_reg_reg_12__2__CLK (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_HCLK_X (.DIODE(clknet_leaf_5_HCLK),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0__f_usb_cdc_clk_48MHz_X (.DIODE(clknet_1_0__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_usb_cdc_clk_48MHz_A (.DIODE(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1__f_usb_cdc_clk_48MHz_X (.DIODE(clknet_1_1__leaf_usb_cdc_clk_48MHz),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(n2440),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\inst_to_wrap_u_usb_cdc_u_bulk_endp_u_async_app_rstn_app_rstn_sq[0] ),
    .VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .X(net364));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_0_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_64 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_0_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_0_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_0_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_0_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_0_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_0_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_0_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_0_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_1_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_1_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_241 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_1_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_417 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_1_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_1_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_1_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_2_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_2_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_164 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_2_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_2_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_2_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_2_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_2_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_333 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_345 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_2_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_2_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_2_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_2_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_2_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_129 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_3_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_3_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_3_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_185 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_3_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_266 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_3_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_417 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_3_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_3_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_3_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_3_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_3_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_3_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_4_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_4_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_4_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_4_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_145 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_171 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_4_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_4_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_271 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_4_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_333 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_345 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_4_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_4_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_4_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_4_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_4_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_5_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_77 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_89 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_5_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_5_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_5_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_178 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_5_190 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_232 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_240 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_5_252 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_5_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_308 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_5_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_417 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_5_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_5_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_5_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_5_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_5_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_6_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_6_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_6_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_6_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_6_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_6_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_325 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_6_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_6_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_6_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_6_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_6_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_6_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_37 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_7_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_7_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_266 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_315 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_7_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_7_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_7_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_430 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_7_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_7_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_7_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_7_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_7_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_8_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_8_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_8_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_342 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_8_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_8_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_8_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_443 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_8_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_464 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_8_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_8_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_8_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_8_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_8_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_50 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_146 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_285 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_302 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_314 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_9_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_9_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_9_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_9_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_9_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_9_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_9_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_9_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_9_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_9_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_9_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_9_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_111 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_10_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_10_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_10_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_10_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_10_450 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_497 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_509 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_10_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_10_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_10_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_10_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_648 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_660 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_672 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_684 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_10_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_10_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_10_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_10_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_66 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_129 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_11_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_182 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_11_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_11_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_288 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_11_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_11_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_11_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_11_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_11_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_11_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_11_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_11_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_11_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_11_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_58 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_12_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_76 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_12_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_127 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_12_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_12_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_12_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_12_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_497 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_509 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_12_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_12_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_12_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_12_676 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_688 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_12_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_12_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_68 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_136 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_13_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_241 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_262 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_288 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_13_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_13_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_401 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_13_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_484 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_13_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_13_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_13_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_13_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_13_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_667 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_13_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_13_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_13_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_13_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_13_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_16 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_49 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_14_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_92 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_14_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_446 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_14_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_14_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_560 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_572 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_14_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_14_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_14_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_618 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_14_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_631 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_14_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_14_666 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_14_674 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_14_696 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_14_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_14_721 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_24 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_15_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_456 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_15_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_15_488 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_15_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_15_605 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_15_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_15_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_15_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_15_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_16_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_147 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_16_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_173 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_16_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_16_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_16_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_16_547 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_16_567 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_592 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_16_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_16_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_17_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_17_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_17_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_270 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_17_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_17_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_17_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_17_668 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_17_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_688 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_17_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_51 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_18_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_18_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_205 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_236 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_18_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_380 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_18_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_18_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_18_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_18_556 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_568 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_18_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_18_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_620 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_632 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_18_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_18_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_18_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_142 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_19_233 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_320 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_464 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_479 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_512 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_516 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_19_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_594 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_644 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_19_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_19_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_19_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_19_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_19_717 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_19_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_19_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_123 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_156 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_174 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_20_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_222 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_280 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_379 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_20_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_20_522 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_554 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_20_566 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_20_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_20_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_20_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_638 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_20_685 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_20_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_20_717 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_20_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_63 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_132 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_21_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_21_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_552 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_21_592 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_21_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_21_628 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_21_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_21_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_21_720 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_21_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_367 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_458 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_22_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_22_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_548 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_574 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_22_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_22_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_22_615 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_22_627 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_22_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_22_672 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_22_708 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_22_730 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_17 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_34 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_38 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_77 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_120 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_23_132 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_23_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_23_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_200 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_23_637 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_23_649 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_23_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_23_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_23_678 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_23_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_23_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_60 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_134 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_24_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_24_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_176 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_212 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_255 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_24_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_481 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_24_575 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_24_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_24_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_24_728 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_24_732 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_25_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_25_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_207 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_25_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_321 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_380 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_25_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_456 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_467 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_25_479 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_511 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_548 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_25_571 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_25_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_25_705 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_25_717 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_25_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_25_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_26_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_70 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_26_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_202 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_26_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_463 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_26_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_26_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_26_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_26_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_530 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_541 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_26_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_26_603 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_26_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_26_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_26_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_26_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_95 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_27_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_27_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_27_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_495 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_542 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_27_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_27_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_602 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_27_610 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_27_623 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_27_635 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_27_647 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_680 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_27_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_27_718 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_27_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_27_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_87 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_167 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_179 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_28_237 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_347 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_368 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_28_380 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_392 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_400 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_28_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_28_500 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_508 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_567 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_579 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_28_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_609 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_28_621 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_632 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_28_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_28_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_28_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_28_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_28_728 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_28_732 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_29_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_29_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_206 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_230 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_29_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_289 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_29_375 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_398 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_29_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_29_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_29_599 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_29_619 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_29_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_29_660 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_29_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_38 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_30_50 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_30_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_150 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_30_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_30_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_30_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_350 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_30_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_30_506 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_30_535 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_30_547 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_575 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_30_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_30_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_30_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_23 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_40 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_31_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_31_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_157 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_31_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_324 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_339 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_31_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_467 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_31_479 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_483 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_564 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_31_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_658 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_31_666 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_31_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_31_678 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_31_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_698 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_31_713 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_717 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_31_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_32 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_44 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_32_56 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_103 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_179 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_331 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_343 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_32_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_394 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_433 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_472 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_491 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_510 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_520 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_32_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_32_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_32_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_619 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_32_647 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_32_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_32_658 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_32_670 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_32_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_32_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_33 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_42 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_33_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_33_69 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_33_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_33_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_33_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_33_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_33_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_426 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_33_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_33_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_539 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_33_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_33_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_33_660 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_33_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_33_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_33_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_35 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_34_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_34_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_90 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_34_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_149 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_264 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_418 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_34_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_437 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_34_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_518 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_539 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_34_551 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_34_575 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_595 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_616 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_34_622 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_34_665 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_34_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_34_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_86 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_110 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_182 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_274 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_35_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_35_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_378 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_35_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_458 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_35_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_488 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_35_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_35_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_35_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_628 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_658 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_35_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_35_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_677 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_35_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_35_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_35_716 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_35_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_48 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_36_60 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_36_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_125 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_210 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_323 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_360 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_376 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_396 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_442 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_459 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_36_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_36_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_36_652 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_36_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_36_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_36_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_36_695 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_36_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_36_732 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_201 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_297 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_331 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_37_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_377 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_415 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_423 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_431 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_455 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_37_467 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_476 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_480 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_484 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_515 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_521 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_534 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_37_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_552 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_37_576 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_37_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_37_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_37_660 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_680 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_37_692 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_37_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_37_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_35 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_38_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_104 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_38_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_38_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_38_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_168 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_38_180 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_184 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_38_209 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_219 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_38_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_394 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_38_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_506 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_511 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_519 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_38_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_575 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_38_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_593 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_600 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_38_606 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_38_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_38_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_38_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_38_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_38_723 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_38_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_35 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_132 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_39_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_39_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_39_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_235 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_298 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_39_319 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_374 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_39_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_39_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_463 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_470 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_479 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_39_518 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_535 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_539 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_574 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_39_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_39_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_39_659 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_688 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_39_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_39_712 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_39_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_39_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_100 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_253 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_40_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_287 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_369 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_40_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_455 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_40_467 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_490 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_516 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_40_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_40_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_539 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_545 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_40_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_611 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_40_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_40_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_40_675 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_40_714 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_40_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_40_732 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_18 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_41_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_41_136 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_41_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_41_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_203 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_41_215 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_245 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_41_257 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_320 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_41_332 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_360 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_41_374 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_41_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_41_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_41_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_41_571 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_41_583 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_640 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_664 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_41_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_41_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_723 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_41_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_41_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_107 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_42_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_42_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_172 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_42_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_42_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_42_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_291 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_314 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_42_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_457 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_42_462 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_42_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_513 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_42_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_546 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_42_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_42_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_42_666 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_42_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_42_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_43_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_72 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_43_84 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_43_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_122 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_43_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_229 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_43_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_284 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_43_294 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_300 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_43_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_364 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_43_376 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_43_388 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_413 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_43_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_487 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_43_499 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_511 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_540 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_43_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_43_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_594 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_598 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_43_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_638 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_650 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_43_676 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_43_714 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_43_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_43_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_44_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_26 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_36 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_44_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_124 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_176 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_44_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_44_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_290 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_44_302 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_316 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_328 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_340 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_352 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_44_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_44_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_427 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_44_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_499 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_511 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_44_523 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_570 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_44_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_606 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_620 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_628 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_44_636 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_44_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_44_686 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_44_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_44_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_44_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_45_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_82 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_45_94 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_45_106 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_119 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_45_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_45_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_190 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_45_202 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_45_214 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_45_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_45_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_326 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_45_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_384 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_429 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_458 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_490 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_45_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_526 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_45_554 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_568 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_45_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_634 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_650 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_45_662 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_684 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_45_696 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_45_708 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_45_716 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_45_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_7 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_46_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_123 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_46_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_170 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_234 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_242 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_259 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_46_287 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_46_299 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_340 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_398 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_495 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_526 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_576 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_584 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_604 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_622 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_639 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_46_652 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_46_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_46_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_46_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_46_704 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_46_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_47_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_30 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_47_42 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_47_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_47_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_47_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_47_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_47_155 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_199 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_260 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_267 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_296 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_47_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_374 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_47_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_47_434 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_440 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_484 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_47_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_518 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_47_570 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_47_582 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_633 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_47_642 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_47_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_47_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_47_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_48_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_48_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_48_41 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_65 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_48_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_138 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_266 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_48_278 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_286 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_356 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_385 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_48_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_48_404 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_48_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_48_441 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_48_453 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_48_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_48_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_48_566 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_48_578 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_48_612 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_624 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_48_638 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_662 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_48_690 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_48_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_48_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_49_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_271 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_347 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_410 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_49_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_461 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_495 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_532 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_536 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_49_563 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_571 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_601 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_49_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_49_646 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_49_658 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_49_680 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_688 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_692 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_49_701 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_49_722 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_49_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_50_62 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_96 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_50_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_194 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_314 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_50_322 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_338 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_50_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_351 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_50_359 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_50_411 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_50_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_50_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_533 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_548 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_562 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_50_574 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_50_586 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_50_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_50_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_50_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_50_717 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_50_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_75 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_51_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_153 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_159 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_268 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_308 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_325 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_364 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_374 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_51_413 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_51_425 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_478 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_482 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_51_550 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_51_591 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_614 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_620 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_51_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_679 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_683 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_51_687 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_51_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_51_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_20 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_45 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_52_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_96 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_52_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_128 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_144 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_52_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_52_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_52_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_52_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_485 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_52_548 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_52_560 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_596 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_52_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_625 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_52_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_52_730 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_53_47 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_135 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_53_147 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_160 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_183 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_244 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_283 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_293 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_53_312 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_330 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_53_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_422 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_53_436 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_53_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_538 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_53_588 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_594 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_53_607 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_636 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_53_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_53_684 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_53_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_53_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_101 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_188 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_230 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_54_239 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_250 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_261 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_306 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_54_327 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_54_336 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_344 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_54_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_54_372 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_54_404 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_54_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_421 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_54_438 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_54_450 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_54_462 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_468 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_54_519 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_54_558 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_577 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_54_626 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_54_672 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_54_689 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_54_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_54_722 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_54_730 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_71 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_100 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_55_119 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_132 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_55_150 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_272 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_292 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_313 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_346 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_55_365 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_371 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_402 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_55_414 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_420 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_443 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_455 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_55_463 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_55_486 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_496 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_55_508 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_55_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_55_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_569 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_595 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_611 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_55_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_658 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_55_670 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_55_692 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_55_712 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_55_724 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_55_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_79 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_94 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_102 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_227 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_231 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_318 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_328 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_334 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_362 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_383 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_56_395 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_56_407 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_416 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_56_428 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_432 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_466 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_474 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_477 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_560 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_56_572 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_56_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_617 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_56_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_56_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_56_657 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_663 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_56_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_56_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_56_732 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_73 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_57_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_57_162 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_57_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_316 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_382 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_390 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_489 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_502 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_57_507 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_57_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_608 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_57_629 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_57_636 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_57_648 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_682 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_57_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_57_720 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_57_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_154 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_58_175 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_219 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_269 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_290 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_58_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_315 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_343 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_58_355 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_446 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_484 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_539 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_58_580 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_618 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_58_623 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_58_635 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_58_666 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_675 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_58_691 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_58_712 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_58_720 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_14 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_74 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_82 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_90 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_117 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_281 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_304 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_341 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_349 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_353 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_381 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_59_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_436 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_459 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_480 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_59_492 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_505 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_59_543 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_59_555 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_59_561 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_567 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_623 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_631 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_673 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_59_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_59_718 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_59_726 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_59_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_80 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_114 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_152 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_218 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_226 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_267 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_60_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_342 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_383 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_60_395 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_399 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_402 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_60_435 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_486 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_60_498 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_60_504 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_516 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_60_528 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_60_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_60_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_60_565 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_60_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_60_684 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_60_721 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_61_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_98 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_61_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_61_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_337 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_345 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_61_386 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_475 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_61_487 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_61_525 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_61_537 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_61_549 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_61_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_61_573 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_61_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_619 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_61_627 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_61_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_61_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_61_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_62_59 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_67 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_62_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_224 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_228 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_62_265 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_317 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_354 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_385 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_62_397 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_437 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_62_449 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_479 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_491 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_503 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_515 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_62_527 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_62_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_62_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_62_589 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_62_597 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_62_612 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_62_624 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_62_636 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_645 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_62_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_43 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_63_64 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_72 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_129 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_135 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_175 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_63_187 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_211 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_240 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_366 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_387 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_2 FILLER_63_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_63_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_63_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_63_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_63_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_63_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_63_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_63_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_63_653 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_661 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_63_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_675 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_63_681 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_63_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_63_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_63_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_59 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_71 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_64_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_64_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_126 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_64_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_166 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_64_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_186 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_255 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_64_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_64_311 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_343 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_64_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_64_393 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_64_406 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_412 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_423 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_435 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_447 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_459 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_64_471 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_64_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_64_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_64_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_64_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_64_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_64_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_64_721 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_65_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_31 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_42 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_65_49 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_65_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_83 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_65_95 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_99 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_107 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_121 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_65_181 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_65_207 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_220 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_65_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_252 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_264 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_65_276 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_283 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_65_295 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_65_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_65_405 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_409 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_432 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_65_444 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_65_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_65_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_65_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_65_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_65_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_65_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_65_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_65_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_65_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_36 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_52 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_66_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_66_141 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_178 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_66_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_255 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_267 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_279 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_291 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_66_303 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_66_309 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_333 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_345 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_66_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_66_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_66_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_66_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_66_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_67_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_11 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_67_30 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_67_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_67_70 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_80 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_67_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_67_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_177 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_192 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_67_208 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_263 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_67_275 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_417 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_67_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_67_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_67_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_67_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_67_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_68_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_45 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_68_78 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_68_92 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_120 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_68_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_131 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_68_163 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_171 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_68_204 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_269 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_68_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_333 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_345 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_68_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_68_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_68_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_68_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_68_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_44 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_69_97 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_127 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_69_158 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_69_166 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_196 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_225 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_69_243 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_69_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_417 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_69_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_69_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_69_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_69_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_69_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_70_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_73 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_70_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_70_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_70_118 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_148 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_156 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_168 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_174 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_70_191 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_213 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_70_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_333 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_345 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_70_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_70_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_70_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_70_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_70_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_34 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_71_46 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_54 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_73 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_71_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 FILLER_71_93 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_113 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_130 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_164 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_71_169 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_71_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_71_222 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_417 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_71_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_71_709 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_71_721 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_71_727 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_71_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_72_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_72_85 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_91 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_8 FILLER_72_108 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_116 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_124 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_72_136 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_148 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_160 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_172 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_184 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_72_197 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_212 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_224 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_236 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_72_248 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_333 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_345 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_72_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_72_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_72_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_72_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_72_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_27 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_39 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_4 FILLER_73_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_81 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_93 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_105 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_111 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_137 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_149 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_161 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_167 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_193 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_205 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_217 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_223 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_249 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_261 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_273 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_279 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_305 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_317 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_329 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_335 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_361 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_373 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_385 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_391 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_417 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_429 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_441 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_447 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_473 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_485 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_497 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_503 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_529 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_541 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_553 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_559 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_585 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_597 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_609 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_615 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_641 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_653 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_73_665 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_73_671 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_73_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_73_697 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_73_709 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_2 FILLER_73_731 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_74_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_53 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_65 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_77 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_83 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_109 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_121 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_133 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_139 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_165 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_177 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_189 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_195 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_221 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_233 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_245 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_251 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_277 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_289 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_301 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_307 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_333 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_345 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_357 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_363 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_389 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_401 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_413 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_419 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_445 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_457 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_469 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_475 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_501 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_513 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_525 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_531 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_557 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_569 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_581 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_587 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_613 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_625 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_637 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_643 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_669 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_681 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_6 FILLER_74_693 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_74_699 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_74_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_74_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_8 FILLER_74_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_3 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_15 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__fill_1 FILLER_75_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_29 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_41 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_53 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_57 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_69 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_81 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_85 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_97 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_109 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_113 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_125 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_137 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_141 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_153 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_165 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_169 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_181 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_193 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_197 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_209 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_221 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_225 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_237 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_249 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_253 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_265 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_277 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_281 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_293 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_305 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_309 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_321 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_333 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_337 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_349 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_361 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_365 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_377 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_389 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_393 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_405 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_417 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_421 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_433 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_445 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_449 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_461 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_473 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_477 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_489 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_501 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_505 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_517 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_529 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_533 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_545 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_557 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_561 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_573 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_585 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_589 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_601 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_613 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_617 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_629 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_641 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_645 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_657 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_669 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_673 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_685 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_697 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_ef_sc_hd__decap_12 FILLER_75_701 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_ef_sc_hd__decap_12 FILLER_75_713 (.VPWR(VPWR),
    .VGND(VGND),
    .VPB(VPWR),
    .VNB(VGND));
 sky130_fd_sc_hd__decap_3 FILLER_75_725 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_75_729 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
endmodule
