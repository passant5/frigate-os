magic
tech sky130A
magscale 1 2
timestamp 1750121950
<< viali >>
rect 1225 1989 1259 2023
rect 8217 1989 8251 2023
rect 1041 1921 1075 1955
rect 1685 1921 1719 1955
rect 1961 1921 1995 1955
rect 2329 1921 2363 1955
rect 2789 1921 2823 1955
rect 3157 1921 3191 1955
rect 3433 1921 3467 1955
rect 3709 1921 3743 1955
rect 4261 1921 4295 1955
rect 4813 1921 4847 1955
rect 5365 1921 5399 1955
rect 5733 1921 5767 1955
rect 6285 1921 6319 1955
rect 6837 1921 6871 1955
rect 7389 1921 7423 1955
rect 7941 1921 7975 1955
rect 8493 1921 8527 1955
rect 8769 1921 8803 1955
rect 9045 1921 9079 1955
rect 9321 1921 9355 1955
rect 9597 1921 9631 1955
rect 9873 1921 9907 1955
rect 10701 1921 10735 1955
rect 11529 1921 11563 1955
rect 12081 1921 12115 1955
rect 14105 1921 14139 1955
rect 15209 1921 15243 1955
rect 16681 1921 16715 1955
rect 17417 1921 17451 1955
rect 17785 1921 17819 1955
rect 18705 1921 18739 1955
rect 1409 1853 1443 1887
rect 2237 1853 2271 1887
rect 3801 1853 3835 1887
rect 5825 1853 5859 1887
rect 6377 1853 6411 1887
rect 6929 1853 6963 1887
rect 9965 1853 9999 1887
rect 10977 1853 11011 1887
rect 12633 1853 12667 1887
rect 14657 1853 14691 1887
rect 16405 1853 16439 1887
rect 18429 1853 18463 1887
rect 18981 1853 19015 1887
rect 4353 1785 4387 1819
rect 5089 1785 5123 1819
rect 7481 1785 7515 1819
rect 11253 1785 11287 1819
rect 12357 1785 12391 1819
rect 13277 1785 13311 1819
rect 13553 1785 13587 1819
rect 15853 1785 15887 1819
rect 18061 1785 18095 1819
rect 10241 1717 10275 1751
rect 11805 1717 11839 1751
rect 12909 1717 12943 1751
rect 13829 1717 13863 1751
rect 14381 1717 14415 1751
rect 14933 1717 14967 1751
rect 15485 1717 15519 1751
rect 16129 1717 16163 1751
rect 16957 1717 16991 1751
rect 17509 1717 17543 1751
rect 19257 1717 19291 1751
rect 1685 1513 1719 1547
rect 1777 1513 1811 1547
rect 2329 1513 2363 1547
rect 2881 1513 2915 1547
rect 3249 1513 3283 1547
rect 3801 1513 3835 1547
rect 4169 1513 4203 1547
rect 4353 1513 4387 1547
rect 4721 1513 4755 1547
rect 5089 1513 5123 1547
rect 5733 1513 5767 1547
rect 6285 1513 6319 1547
rect 6929 1513 6963 1547
rect 7297 1513 7331 1547
rect 7481 1513 7515 1547
rect 7849 1513 7883 1547
rect 8217 1513 8251 1547
rect 8585 1513 8619 1547
rect 9045 1513 9079 1547
rect 9505 1513 9539 1547
rect 10057 1513 10091 1547
rect 10241 1513 10275 1547
rect 10701 1513 10735 1547
rect 11529 1513 11563 1547
rect 11713 1513 11747 1547
rect 11989 1513 12023 1547
rect 12265 1513 12299 1547
rect 12633 1513 12667 1547
rect 13185 1513 13219 1547
rect 13737 1513 13771 1547
rect 14289 1513 14323 1547
rect 14841 1513 14875 1547
rect 15209 1513 15243 1547
rect 15853 1513 15887 1547
rect 16313 1513 16347 1547
rect 16865 1513 16899 1547
rect 17417 1513 17451 1547
rect 17785 1513 17819 1547
rect 18337 1513 18371 1547
rect 19165 1513 19199 1547
rect 19349 1513 19383 1547
rect 9137 1445 9171 1479
rect 10977 1445 11011 1479
rect 14013 1445 14047 1479
rect 16129 1445 16163 1479
rect 18613 1445 18647 1479
rect 2237 1377 2271 1411
rect 2789 1377 2823 1411
rect 3709 1377 3743 1411
rect 5825 1377 5859 1411
rect 6377 1377 6411 1411
rect 18981 1377 19015 1411
rect 11253 1309 11287 1343
rect 12909 1309 12943 1343
rect 14565 1309 14599 1343
rect 15485 1309 15519 1343
rect 17141 1309 17175 1343
rect 18797 1309 18831 1343
rect 6837 1241 6871 1275
rect 13461 1241 13495 1275
rect 16589 1241 16623 1275
rect 18061 1241 18095 1275
rect 9689 1173 9723 1207
rect 2513 969 2547 1003
rect 2789 969 2823 1003
rect 2973 969 3007 1003
rect 3341 969 3375 1003
rect 3525 969 3559 1003
rect 3893 969 3927 1003
rect 4261 969 4295 1003
rect 4445 969 4479 1003
rect 4629 969 4663 1003
rect 4813 969 4847 1003
rect 5273 969 5307 1003
rect 5549 969 5583 1003
rect 5917 969 5951 1003
rect 6469 969 6503 1003
rect 7021 969 7055 1003
rect 7573 969 7607 1003
rect 8217 969 8251 1003
rect 8677 969 8711 1003
rect 9413 969 9447 1003
rect 11989 969 12023 1003
rect 12541 969 12575 1003
rect 12909 969 12943 1003
rect 13829 969 13863 1003
rect 14105 969 14139 1003
rect 14749 969 14783 1003
rect 14933 969 14967 1003
rect 15577 969 15611 1003
rect 16313 969 16347 1003
rect 16681 969 16715 1003
rect 17325 969 17359 1003
rect 17693 969 17727 1003
rect 18153 969 18187 1003
rect 18613 969 18647 1003
rect 19257 969 19291 1003
rect 3985 901 4019 935
rect 6101 901 6135 935
rect 6653 901 6687 935
rect 7205 901 7239 935
rect 7757 901 7791 935
rect 8861 901 8895 935
rect 12449 901 12483 935
rect 13553 901 13587 935
rect 14565 901 14599 935
rect 15301 901 15335 935
rect 16129 901 16163 935
rect 17141 901 17175 935
rect 4997 833 5031 867
rect 9045 833 9079 867
rect 13277 833 13311 867
rect 14381 833 14415 867
rect 15393 833 15427 867
rect 16957 833 16991 867
rect 8309 765 8343 799
<< metal1 >>
rect 18046 2456 18052 2508
rect 18104 2496 18110 2508
rect 18966 2496 18972 2508
rect 18104 2468 18972 2496
rect 18104 2456 18110 2468
rect 18966 2456 18972 2468
rect 19024 2456 19030 2508
rect 1578 2320 1584 2372
rect 1636 2360 1642 2372
rect 1854 2360 1860 2372
rect 1636 2332 1860 2360
rect 1636 2320 1642 2332
rect 1854 2320 1860 2332
rect 1912 2320 1918 2372
rect 17126 2320 17132 2372
rect 17184 2360 17190 2372
rect 18322 2360 18328 2372
rect 17184 2332 18328 2360
rect 17184 2320 17190 2332
rect 18322 2320 18328 2332
rect 18380 2320 18386 2372
rect 276 2202 19780 2224
rect 276 2150 1122 2202
rect 1174 2150 1186 2202
rect 1238 2150 1250 2202
rect 1302 2150 1314 2202
rect 1366 2150 1378 2202
rect 1430 2150 9122 2202
rect 9174 2150 9186 2202
rect 9238 2150 9250 2202
rect 9302 2150 9314 2202
rect 9366 2150 9378 2202
rect 9430 2150 17122 2202
rect 17174 2150 17186 2202
rect 17238 2150 17250 2202
rect 17302 2150 17314 2202
rect 17366 2150 17378 2202
rect 17430 2150 19780 2202
rect 276 2128 19780 2150
rect 13446 2048 13452 2100
rect 13504 2088 13510 2100
rect 14274 2088 14280 2100
rect 13504 2060 14280 2088
rect 13504 2048 13510 2060
rect 14274 2048 14280 2060
rect 14332 2048 14338 2100
rect 14550 2048 14556 2100
rect 14608 2088 14614 2100
rect 15194 2088 15200 2100
rect 14608 2060 15200 2088
rect 14608 2048 14614 2060
rect 15194 2048 15200 2060
rect 15252 2048 15258 2100
rect 16942 2048 16948 2100
rect 17000 2088 17006 2100
rect 17000 2060 17816 2088
rect 17000 2048 17006 2060
rect 1213 2023 1271 2029
rect 1213 1989 1225 2023
rect 1259 2020 1271 2023
rect 8205 2023 8263 2029
rect 1259 1992 1992 2020
rect 1259 1989 1271 1992
rect 1213 1983 1271 1989
rect 1029 1955 1087 1961
rect 1029 1921 1041 1955
rect 1075 1952 1087 1955
rect 1578 1952 1584 1964
rect 1075 1924 1584 1952
rect 1075 1921 1087 1924
rect 1029 1915 1087 1921
rect 1578 1912 1584 1924
rect 1636 1952 1642 1964
rect 1964 1961 1992 1992
rect 8205 1989 8217 2023
rect 8251 2020 8263 2023
rect 8251 1992 8800 2020
rect 8251 1989 8263 1992
rect 8205 1983 8263 1989
rect 1673 1955 1731 1961
rect 1673 1952 1685 1955
rect 1636 1924 1685 1952
rect 1636 1912 1642 1924
rect 1673 1921 1685 1924
rect 1719 1921 1731 1955
rect 1673 1915 1731 1921
rect 1949 1955 2007 1961
rect 1949 1921 1961 1955
rect 1995 1952 2007 1955
rect 2130 1952 2136 1964
rect 1995 1924 2136 1952
rect 1995 1921 2007 1924
rect 1949 1915 2007 1921
rect 2130 1912 2136 1924
rect 2188 1912 2194 1964
rect 2317 1955 2375 1961
rect 2317 1921 2329 1955
rect 2363 1952 2375 1955
rect 2590 1952 2596 1964
rect 2363 1924 2596 1952
rect 2363 1921 2375 1924
rect 2317 1915 2375 1921
rect 2590 1912 2596 1924
rect 2648 1912 2654 1964
rect 2777 1955 2835 1961
rect 2777 1921 2789 1955
rect 2823 1952 2835 1955
rect 2958 1952 2964 1964
rect 2823 1924 2964 1952
rect 2823 1921 2835 1924
rect 2777 1915 2835 1921
rect 2958 1912 2964 1924
rect 3016 1912 3022 1964
rect 3145 1955 3203 1961
rect 3145 1921 3157 1955
rect 3191 1952 3203 1955
rect 3326 1952 3332 1964
rect 3191 1924 3332 1952
rect 3191 1921 3203 1924
rect 3145 1915 3203 1921
rect 3326 1912 3332 1924
rect 3384 1912 3390 1964
rect 3421 1955 3479 1961
rect 3421 1921 3433 1955
rect 3467 1952 3479 1955
rect 3510 1952 3516 1964
rect 3467 1924 3516 1952
rect 3467 1921 3479 1924
rect 3421 1915 3479 1921
rect 3510 1912 3516 1924
rect 3568 1912 3574 1964
rect 3697 1955 3755 1961
rect 3697 1921 3709 1955
rect 3743 1952 3755 1955
rect 3878 1952 3884 1964
rect 3743 1924 3884 1952
rect 3743 1921 3755 1924
rect 3697 1915 3755 1921
rect 3878 1912 3884 1924
rect 3936 1912 3942 1964
rect 4249 1955 4307 1961
rect 4249 1921 4261 1955
rect 4295 1952 4307 1955
rect 4430 1952 4436 1964
rect 4295 1924 4436 1952
rect 4295 1921 4307 1924
rect 4249 1915 4307 1921
rect 4430 1912 4436 1924
rect 4488 1912 4494 1964
rect 4801 1955 4859 1961
rect 4801 1921 4813 1955
rect 4847 1952 4859 1955
rect 5166 1952 5172 1964
rect 4847 1924 5172 1952
rect 4847 1921 4859 1924
rect 4801 1915 4859 1921
rect 5166 1912 5172 1924
rect 5224 1912 5230 1964
rect 5353 1955 5411 1961
rect 5353 1921 5365 1955
rect 5399 1952 5411 1955
rect 5534 1952 5540 1964
rect 5399 1924 5540 1952
rect 5399 1921 5411 1924
rect 5353 1915 5411 1921
rect 5534 1912 5540 1924
rect 5592 1912 5598 1964
rect 5721 1955 5779 1961
rect 5721 1921 5733 1955
rect 5767 1952 5779 1955
rect 5902 1952 5908 1964
rect 5767 1924 5908 1952
rect 5767 1921 5779 1924
rect 5721 1915 5779 1921
rect 5902 1912 5908 1924
rect 5960 1912 5966 1964
rect 6273 1955 6331 1961
rect 6273 1921 6285 1955
rect 6319 1952 6331 1955
rect 6454 1952 6460 1964
rect 6319 1924 6460 1952
rect 6319 1921 6331 1924
rect 6273 1915 6331 1921
rect 6454 1912 6460 1924
rect 6512 1912 6518 1964
rect 6825 1955 6883 1961
rect 6825 1921 6837 1955
rect 6871 1952 6883 1955
rect 7006 1952 7012 1964
rect 6871 1924 7012 1952
rect 6871 1921 6883 1924
rect 6825 1915 6883 1921
rect 7006 1912 7012 1924
rect 7064 1912 7070 1964
rect 7377 1955 7435 1961
rect 7377 1921 7389 1955
rect 7423 1952 7435 1955
rect 7558 1952 7564 1964
rect 7423 1924 7564 1952
rect 7423 1921 7435 1924
rect 7377 1915 7435 1921
rect 7558 1912 7564 1924
rect 7616 1912 7622 1964
rect 7929 1955 7987 1961
rect 7929 1921 7941 1955
rect 7975 1952 7987 1955
rect 8294 1952 8300 1964
rect 7975 1924 8300 1952
rect 7975 1921 7987 1924
rect 7929 1915 7987 1921
rect 8294 1912 8300 1924
rect 8352 1912 8358 1964
rect 8481 1955 8539 1961
rect 8481 1921 8493 1955
rect 8527 1952 8539 1955
rect 8662 1952 8668 1964
rect 8527 1924 8668 1952
rect 8527 1921 8539 1924
rect 8481 1915 8539 1921
rect 8662 1912 8668 1924
rect 8720 1912 8726 1964
rect 8772 1961 8800 1992
rect 11238 1980 11244 2032
rect 11296 2020 11302 2032
rect 11296 1992 12112 2020
rect 11296 1980 11302 1992
rect 12084 1964 12112 1992
rect 12710 1980 12716 2032
rect 12768 2020 12774 2032
rect 13538 2020 13544 2032
rect 12768 1992 13544 2020
rect 12768 1980 12774 1992
rect 13538 1980 13544 1992
rect 13596 1980 13602 2032
rect 16390 1980 16396 2032
rect 16448 2020 16454 2032
rect 17788 2020 17816 2060
rect 18782 2020 18788 2032
rect 16448 1992 17448 2020
rect 16448 1980 16454 1992
rect 8757 1955 8815 1961
rect 8757 1921 8769 1955
rect 8803 1952 8815 1955
rect 8846 1952 8852 1964
rect 8803 1924 8852 1952
rect 8803 1921 8815 1924
rect 8757 1915 8815 1921
rect 8846 1912 8852 1924
rect 8904 1912 8910 1964
rect 9030 1912 9036 1964
rect 9088 1912 9094 1964
rect 9309 1955 9367 1961
rect 9309 1921 9321 1955
rect 9355 1952 9367 1955
rect 9490 1952 9496 1964
rect 9355 1924 9496 1952
rect 9355 1921 9367 1924
rect 9309 1915 9367 1921
rect 9490 1912 9496 1924
rect 9548 1912 9554 1964
rect 9582 1912 9588 1964
rect 9640 1912 9646 1964
rect 9861 1955 9919 1961
rect 9861 1921 9873 1955
rect 9907 1952 9919 1955
rect 10134 1952 10140 1964
rect 9907 1924 10140 1952
rect 9907 1921 9919 1924
rect 9861 1915 9919 1921
rect 10134 1912 10140 1924
rect 10192 1912 10198 1964
rect 10410 1912 10416 1964
rect 10468 1952 10474 1964
rect 10689 1955 10747 1961
rect 10689 1952 10701 1955
rect 10468 1924 10701 1952
rect 10468 1912 10474 1924
rect 10689 1921 10701 1924
rect 10735 1921 10747 1955
rect 10689 1915 10747 1921
rect 10870 1912 10876 1964
rect 10928 1952 10934 1964
rect 11517 1955 11575 1961
rect 11517 1952 11529 1955
rect 10928 1924 11529 1952
rect 10928 1912 10934 1924
rect 11517 1921 11529 1924
rect 11563 1952 11575 1955
rect 11974 1952 11980 1964
rect 11563 1924 11980 1952
rect 11563 1921 11575 1924
rect 11517 1915 11575 1921
rect 11974 1912 11980 1924
rect 12032 1912 12038 1964
rect 12066 1912 12072 1964
rect 12124 1912 12130 1964
rect 13262 1912 13268 1964
rect 13320 1952 13326 1964
rect 14093 1955 14151 1961
rect 14093 1952 14105 1955
rect 13320 1924 14105 1952
rect 13320 1912 13326 1924
rect 14093 1921 14105 1924
rect 14139 1952 14151 1955
rect 14366 1952 14372 1964
rect 14139 1924 14372 1952
rect 14139 1921 14151 1924
rect 14093 1915 14151 1921
rect 14366 1912 14372 1924
rect 14424 1912 14430 1964
rect 14458 1912 14464 1964
rect 14516 1952 14522 1964
rect 15197 1955 15255 1961
rect 15197 1952 15209 1955
rect 14516 1924 15209 1952
rect 14516 1912 14522 1924
rect 15197 1921 15209 1924
rect 15243 1952 15255 1955
rect 15746 1952 15752 1964
rect 15243 1924 15752 1952
rect 15243 1921 15255 1924
rect 15197 1915 15255 1921
rect 15746 1912 15752 1924
rect 15804 1912 15810 1964
rect 15838 1912 15844 1964
rect 15896 1952 15902 1964
rect 16669 1955 16727 1961
rect 16669 1952 16681 1955
rect 15896 1924 16681 1952
rect 15896 1912 15902 1924
rect 16669 1921 16681 1924
rect 16715 1952 16727 1955
rect 16942 1952 16948 1964
rect 16715 1924 16948 1952
rect 16715 1921 16727 1924
rect 16669 1915 16727 1921
rect 16942 1912 16948 1924
rect 17000 1912 17006 1964
rect 17420 1961 17448 1992
rect 17788 1992 18788 2020
rect 17788 1961 17816 1992
rect 18782 1980 18788 1992
rect 18840 1980 18846 2032
rect 17405 1955 17463 1961
rect 17405 1921 17417 1955
rect 17451 1921 17463 1955
rect 17405 1915 17463 1921
rect 17773 1955 17831 1961
rect 17773 1921 17785 1955
rect 17819 1921 17831 1955
rect 17773 1915 17831 1921
rect 1397 1887 1455 1893
rect 1397 1853 1409 1887
rect 1443 1884 1455 1887
rect 2225 1887 2283 1893
rect 2225 1884 2237 1887
rect 1443 1856 2237 1884
rect 1443 1853 1455 1856
rect 1397 1847 1455 1853
rect 2225 1853 2237 1856
rect 2271 1884 2283 1887
rect 2406 1884 2412 1896
rect 2271 1856 2412 1884
rect 2271 1853 2283 1856
rect 2225 1847 2283 1853
rect 2406 1844 2412 1856
rect 2464 1844 2470 1896
rect 3789 1887 3847 1893
rect 3789 1853 3801 1887
rect 3835 1884 3847 1887
rect 4062 1884 4068 1896
rect 3835 1856 4068 1884
rect 3835 1853 3847 1856
rect 3789 1847 3847 1853
rect 4062 1844 4068 1856
rect 4120 1844 4126 1896
rect 5813 1887 5871 1893
rect 5813 1853 5825 1887
rect 5859 1884 5871 1887
rect 6086 1884 6092 1896
rect 5859 1856 6092 1884
rect 5859 1853 5871 1856
rect 5813 1847 5871 1853
rect 6086 1844 6092 1856
rect 6144 1844 6150 1896
rect 6365 1887 6423 1893
rect 6365 1853 6377 1887
rect 6411 1884 6423 1887
rect 6638 1884 6644 1896
rect 6411 1856 6644 1884
rect 6411 1853 6423 1856
rect 6365 1847 6423 1853
rect 6638 1844 6644 1856
rect 6696 1844 6702 1896
rect 6917 1887 6975 1893
rect 6917 1853 6929 1887
rect 6963 1884 6975 1887
rect 7190 1884 7196 1896
rect 6963 1856 7196 1884
rect 6963 1853 6975 1856
rect 6917 1847 6975 1853
rect 7190 1844 7196 1856
rect 7248 1844 7254 1896
rect 9953 1887 10011 1893
rect 9953 1853 9965 1887
rect 9999 1884 10011 1887
rect 10226 1884 10232 1896
rect 9999 1856 10232 1884
rect 9999 1853 10011 1856
rect 9953 1847 10011 1853
rect 10226 1844 10232 1856
rect 10284 1844 10290 1896
rect 10502 1844 10508 1896
rect 10560 1884 10566 1896
rect 10962 1884 10968 1896
rect 10560 1856 10968 1884
rect 10560 1844 10566 1856
rect 10962 1844 10968 1856
rect 11020 1844 11026 1896
rect 11790 1844 11796 1896
rect 11848 1884 11854 1896
rect 12621 1887 12679 1893
rect 12621 1884 12633 1887
rect 11848 1856 12633 1884
rect 11848 1844 11854 1856
rect 12621 1853 12633 1856
rect 12667 1884 12679 1887
rect 12894 1884 12900 1896
rect 12667 1856 12900 1884
rect 12667 1853 12679 1856
rect 12621 1847 12679 1853
rect 12894 1844 12900 1856
rect 12952 1844 12958 1896
rect 12986 1844 12992 1896
rect 13044 1884 13050 1896
rect 13044 1856 13676 1884
rect 13044 1844 13050 1856
rect 4154 1776 4160 1828
rect 4212 1816 4218 1828
rect 4341 1819 4399 1825
rect 4341 1816 4353 1819
rect 4212 1788 4353 1816
rect 4212 1776 4218 1788
rect 4341 1785 4353 1788
rect 4387 1816 4399 1819
rect 4798 1816 4804 1828
rect 4387 1788 4804 1816
rect 4387 1785 4399 1788
rect 4341 1779 4399 1785
rect 4798 1776 4804 1788
rect 4856 1776 4862 1828
rect 5077 1819 5135 1825
rect 5077 1785 5089 1819
rect 5123 1816 5135 1819
rect 5350 1816 5356 1828
rect 5123 1788 5356 1816
rect 5123 1785 5135 1788
rect 5077 1779 5135 1785
rect 5350 1776 5356 1788
rect 5408 1776 5414 1828
rect 7282 1776 7288 1828
rect 7340 1816 7346 1828
rect 7469 1819 7527 1825
rect 7469 1816 7481 1819
rect 7340 1788 7481 1816
rect 7340 1776 7346 1788
rect 7469 1785 7481 1788
rect 7515 1816 7527 1819
rect 7926 1816 7932 1828
rect 7515 1788 7932 1816
rect 7515 1785 7527 1788
rect 7469 1779 7527 1785
rect 7926 1776 7932 1788
rect 7984 1776 7990 1828
rect 10686 1776 10692 1828
rect 10744 1816 10750 1828
rect 11238 1816 11244 1828
rect 10744 1788 11244 1816
rect 10744 1776 10750 1788
rect 11238 1776 11244 1788
rect 11296 1776 11302 1828
rect 11422 1776 11428 1828
rect 11480 1816 11486 1828
rect 12250 1816 12256 1828
rect 11480 1788 12256 1816
rect 11480 1776 11486 1788
rect 12250 1776 12256 1788
rect 12308 1816 12314 1828
rect 12345 1819 12403 1825
rect 12345 1816 12357 1819
rect 12308 1788 12357 1816
rect 12308 1776 12314 1788
rect 12345 1785 12357 1788
rect 12391 1785 12403 1819
rect 12345 1779 12403 1785
rect 12434 1776 12440 1828
rect 12492 1816 12498 1828
rect 13265 1819 13323 1825
rect 13265 1816 13277 1819
rect 12492 1788 13277 1816
rect 12492 1776 12498 1788
rect 13265 1785 13277 1788
rect 13311 1816 13323 1819
rect 13446 1816 13452 1828
rect 13311 1788 13452 1816
rect 13311 1785 13323 1788
rect 13265 1779 13323 1785
rect 13446 1776 13452 1788
rect 13504 1776 13510 1828
rect 13538 1776 13544 1828
rect 13596 1776 13602 1828
rect 10229 1751 10287 1757
rect 10229 1717 10241 1751
rect 10275 1748 10287 1751
rect 10318 1748 10324 1760
rect 10275 1720 10324 1748
rect 10275 1717 10287 1720
rect 10229 1711 10287 1717
rect 10318 1708 10324 1720
rect 10376 1708 10382 1760
rect 11054 1708 11060 1760
rect 11112 1748 11118 1760
rect 11790 1748 11796 1760
rect 11112 1720 11796 1748
rect 11112 1708 11118 1720
rect 11790 1708 11796 1720
rect 11848 1708 11854 1760
rect 11882 1708 11888 1760
rect 11940 1748 11946 1760
rect 12897 1751 12955 1757
rect 12897 1748 12909 1751
rect 11940 1720 12909 1748
rect 11940 1708 11946 1720
rect 12897 1717 12909 1720
rect 12943 1748 12955 1751
rect 13354 1748 13360 1760
rect 12943 1720 13360 1748
rect 12943 1717 12955 1720
rect 12897 1711 12955 1717
rect 13354 1708 13360 1720
rect 13412 1708 13418 1760
rect 13648 1748 13676 1856
rect 13814 1844 13820 1896
rect 13872 1884 13878 1896
rect 14645 1887 14703 1893
rect 14645 1884 14657 1887
rect 13872 1856 14657 1884
rect 13872 1844 13878 1856
rect 14645 1853 14657 1856
rect 14691 1884 14703 1887
rect 14918 1884 14924 1896
rect 14691 1856 14924 1884
rect 14691 1853 14703 1856
rect 14645 1847 14703 1853
rect 14918 1844 14924 1856
rect 14976 1844 14982 1896
rect 15470 1844 15476 1896
rect 15528 1884 15534 1896
rect 16390 1884 16396 1896
rect 15528 1856 16396 1884
rect 15528 1844 15534 1856
rect 16390 1844 16396 1856
rect 16448 1844 16454 1896
rect 13998 1776 14004 1828
rect 14056 1816 14062 1828
rect 14826 1816 14832 1828
rect 14056 1788 14832 1816
rect 14056 1776 14062 1788
rect 14826 1776 14832 1788
rect 14884 1816 14890 1828
rect 14884 1788 14964 1816
rect 14884 1776 14890 1788
rect 13817 1751 13875 1757
rect 13817 1748 13829 1751
rect 13648 1720 13829 1748
rect 13817 1717 13829 1720
rect 13863 1748 13875 1751
rect 14090 1748 14096 1760
rect 13863 1720 14096 1748
rect 13863 1717 13875 1720
rect 13817 1711 13875 1717
rect 14090 1708 14096 1720
rect 14148 1708 14154 1760
rect 14274 1708 14280 1760
rect 14332 1748 14338 1760
rect 14936 1757 14964 1788
rect 15010 1776 15016 1828
rect 15068 1816 15074 1828
rect 15838 1816 15844 1828
rect 15068 1788 15844 1816
rect 15068 1776 15074 1788
rect 15838 1776 15844 1788
rect 15896 1776 15902 1828
rect 16022 1776 16028 1828
rect 16080 1816 16086 1828
rect 16080 1788 16528 1816
rect 16080 1776 16086 1788
rect 14369 1751 14427 1757
rect 14369 1748 14381 1751
rect 14332 1720 14381 1748
rect 14332 1708 14338 1720
rect 14369 1717 14381 1720
rect 14415 1717 14427 1751
rect 14369 1711 14427 1717
rect 14921 1751 14979 1757
rect 14921 1717 14933 1751
rect 14967 1717 14979 1751
rect 14921 1711 14979 1717
rect 15194 1708 15200 1760
rect 15252 1748 15258 1760
rect 15473 1751 15531 1757
rect 15473 1748 15485 1751
rect 15252 1720 15485 1748
rect 15252 1708 15258 1720
rect 15473 1717 15485 1720
rect 15519 1717 15531 1751
rect 15473 1711 15531 1717
rect 15562 1708 15568 1760
rect 15620 1748 15626 1760
rect 16114 1748 16120 1760
rect 15620 1720 16120 1748
rect 15620 1708 15626 1720
rect 16114 1708 16120 1720
rect 16172 1708 16178 1760
rect 16500 1748 16528 1788
rect 16574 1776 16580 1828
rect 16632 1816 16638 1828
rect 17420 1816 17448 1915
rect 18138 1912 18144 1964
rect 18196 1952 18202 1964
rect 18693 1955 18751 1961
rect 18693 1952 18705 1955
rect 18196 1924 18705 1952
rect 18196 1912 18202 1924
rect 18693 1921 18705 1924
rect 18739 1952 18751 1955
rect 19334 1952 19340 1964
rect 18739 1924 19340 1952
rect 18739 1921 18751 1924
rect 18693 1915 18751 1921
rect 19334 1912 19340 1924
rect 19392 1912 19398 1964
rect 17586 1844 17592 1896
rect 17644 1884 17650 1896
rect 18414 1884 18420 1896
rect 17644 1856 18420 1884
rect 17644 1844 17650 1856
rect 18414 1844 18420 1856
rect 18472 1844 18478 1896
rect 18966 1844 18972 1896
rect 19024 1844 19030 1896
rect 18049 1819 18107 1825
rect 16632 1788 17356 1816
rect 17420 1788 17724 1816
rect 16632 1776 16638 1788
rect 16850 1748 16856 1760
rect 16500 1720 16856 1748
rect 16850 1708 16856 1720
rect 16908 1748 16914 1760
rect 16945 1751 17003 1757
rect 16945 1748 16957 1751
rect 16908 1720 16957 1748
rect 16908 1708 16914 1720
rect 16945 1717 16957 1720
rect 16991 1717 17003 1751
rect 17328 1748 17356 1788
rect 17497 1751 17555 1757
rect 17497 1748 17509 1751
rect 17328 1720 17509 1748
rect 16945 1711 17003 1717
rect 17497 1717 17509 1720
rect 17543 1717 17555 1751
rect 17696 1748 17724 1788
rect 18049 1785 18061 1819
rect 18095 1816 18107 1819
rect 18322 1816 18328 1828
rect 18095 1788 18328 1816
rect 18095 1785 18107 1788
rect 18049 1779 18107 1785
rect 18322 1776 18328 1788
rect 18380 1776 18386 1828
rect 19245 1751 19303 1757
rect 19245 1748 19257 1751
rect 17696 1720 19257 1748
rect 17497 1711 17555 1717
rect 19245 1717 19257 1720
rect 19291 1717 19303 1751
rect 19245 1711 19303 1717
rect 276 1658 19780 1680
rect 276 1606 1762 1658
rect 1814 1606 1826 1658
rect 1878 1606 1890 1658
rect 1942 1606 1954 1658
rect 2006 1606 2018 1658
rect 2070 1606 9762 1658
rect 9814 1606 9826 1658
rect 9878 1606 9890 1658
rect 9942 1606 9954 1658
rect 10006 1606 10018 1658
rect 10070 1606 17762 1658
rect 17814 1606 17826 1658
rect 17878 1606 17890 1658
rect 17942 1606 17954 1658
rect 18006 1606 18018 1658
rect 18070 1606 19780 1658
rect 276 1584 19780 1606
rect 1670 1504 1676 1556
rect 1728 1544 1734 1556
rect 1765 1547 1823 1553
rect 1765 1544 1777 1547
rect 1728 1516 1777 1544
rect 1728 1504 1734 1516
rect 1765 1513 1777 1516
rect 1811 1513 1823 1547
rect 1765 1507 1823 1513
rect 2222 1504 2228 1556
rect 2280 1544 2286 1556
rect 2317 1547 2375 1553
rect 2317 1544 2329 1547
rect 2280 1516 2329 1544
rect 2280 1504 2286 1516
rect 2317 1513 2329 1516
rect 2363 1513 2375 1547
rect 2317 1507 2375 1513
rect 2774 1504 2780 1556
rect 2832 1544 2838 1556
rect 2869 1547 2927 1553
rect 2869 1544 2881 1547
rect 2832 1516 2881 1544
rect 2832 1504 2838 1516
rect 2869 1513 2881 1516
rect 2915 1513 2927 1547
rect 2869 1507 2927 1513
rect 3142 1504 3148 1556
rect 3200 1544 3206 1556
rect 3237 1547 3295 1553
rect 3237 1544 3249 1547
rect 3200 1516 3249 1544
rect 3200 1504 3206 1516
rect 3237 1513 3249 1516
rect 3283 1513 3295 1547
rect 3237 1507 3295 1513
rect 3694 1504 3700 1556
rect 3752 1544 3758 1556
rect 3789 1547 3847 1553
rect 3789 1544 3801 1547
rect 3752 1516 3801 1544
rect 3752 1504 3758 1516
rect 3789 1513 3801 1516
rect 3835 1513 3847 1547
rect 3789 1507 3847 1513
rect 4154 1504 4160 1556
rect 4212 1504 4218 1556
rect 4246 1504 4252 1556
rect 4304 1544 4310 1556
rect 4341 1547 4399 1553
rect 4341 1544 4353 1547
rect 4304 1516 4353 1544
rect 4304 1504 4310 1516
rect 4341 1513 4353 1516
rect 4387 1513 4399 1547
rect 4341 1507 4399 1513
rect 4614 1504 4620 1556
rect 4672 1544 4678 1556
rect 4709 1547 4767 1553
rect 4709 1544 4721 1547
rect 4672 1516 4721 1544
rect 4672 1504 4678 1516
rect 4709 1513 4721 1516
rect 4755 1513 4767 1547
rect 4709 1507 4767 1513
rect 4982 1504 4988 1556
rect 5040 1544 5046 1556
rect 5077 1547 5135 1553
rect 5077 1544 5089 1547
rect 5040 1516 5089 1544
rect 5040 1504 5046 1516
rect 5077 1513 5089 1516
rect 5123 1513 5135 1547
rect 5077 1507 5135 1513
rect 5721 1547 5779 1553
rect 5721 1513 5733 1547
rect 5767 1544 5779 1547
rect 6086 1544 6092 1556
rect 5767 1516 6092 1544
rect 5767 1513 5779 1516
rect 5721 1507 5779 1513
rect 6086 1504 6092 1516
rect 6144 1504 6150 1556
rect 6273 1547 6331 1553
rect 6273 1513 6285 1547
rect 6319 1544 6331 1547
rect 6638 1544 6644 1556
rect 6319 1516 6644 1544
rect 6319 1513 6331 1516
rect 6273 1507 6331 1513
rect 6638 1504 6644 1516
rect 6696 1504 6702 1556
rect 6822 1504 6828 1556
rect 6880 1544 6886 1556
rect 6917 1547 6975 1553
rect 6917 1544 6929 1547
rect 6880 1516 6929 1544
rect 6880 1504 6886 1516
rect 6917 1513 6929 1516
rect 6963 1513 6975 1547
rect 6917 1507 6975 1513
rect 7282 1504 7288 1556
rect 7340 1504 7346 1556
rect 7374 1504 7380 1556
rect 7432 1544 7438 1556
rect 7469 1547 7527 1553
rect 7469 1544 7481 1547
rect 7432 1516 7481 1544
rect 7432 1504 7438 1516
rect 7469 1513 7481 1516
rect 7515 1513 7527 1547
rect 7469 1507 7527 1513
rect 7742 1504 7748 1556
rect 7800 1544 7806 1556
rect 7837 1547 7895 1553
rect 7837 1544 7849 1547
rect 7800 1516 7849 1544
rect 7800 1504 7806 1516
rect 7837 1513 7849 1516
rect 7883 1513 7895 1547
rect 7837 1507 7895 1513
rect 8110 1504 8116 1556
rect 8168 1544 8174 1556
rect 8205 1547 8263 1553
rect 8205 1544 8217 1547
rect 8168 1516 8217 1544
rect 8168 1504 8174 1516
rect 8205 1513 8217 1516
rect 8251 1513 8263 1547
rect 8205 1507 8263 1513
rect 8478 1504 8484 1556
rect 8536 1544 8542 1556
rect 8573 1547 8631 1553
rect 8573 1544 8585 1547
rect 8536 1516 8585 1544
rect 8536 1504 8542 1516
rect 8573 1513 8585 1516
rect 8619 1513 8631 1547
rect 8573 1507 8631 1513
rect 9030 1504 9036 1556
rect 9088 1504 9094 1556
rect 9490 1504 9496 1556
rect 9548 1504 9554 1556
rect 10045 1547 10103 1553
rect 10045 1513 10057 1547
rect 10091 1544 10103 1547
rect 10134 1544 10140 1556
rect 10091 1516 10140 1544
rect 10091 1513 10103 1516
rect 10045 1507 10103 1513
rect 10134 1504 10140 1516
rect 10192 1504 10198 1556
rect 10226 1504 10232 1556
rect 10284 1504 10290 1556
rect 10318 1504 10324 1556
rect 10376 1544 10382 1556
rect 10689 1547 10747 1553
rect 10689 1544 10701 1547
rect 10376 1516 10701 1544
rect 10376 1504 10382 1516
rect 10689 1513 10701 1516
rect 10735 1513 10747 1547
rect 10689 1507 10747 1513
rect 11238 1504 11244 1556
rect 11296 1544 11302 1556
rect 11517 1547 11575 1553
rect 11517 1544 11529 1547
rect 11296 1516 11529 1544
rect 11296 1504 11302 1516
rect 11517 1513 11529 1516
rect 11563 1513 11575 1547
rect 11517 1507 11575 1513
rect 11606 1504 11612 1556
rect 11664 1544 11670 1556
rect 11701 1547 11759 1553
rect 11701 1544 11713 1547
rect 11664 1516 11713 1544
rect 11664 1504 11670 1516
rect 11701 1513 11713 1516
rect 11747 1513 11759 1547
rect 11701 1507 11759 1513
rect 11974 1504 11980 1556
rect 12032 1504 12038 1556
rect 12158 1504 12164 1556
rect 12216 1544 12222 1556
rect 12253 1547 12311 1553
rect 12253 1544 12265 1547
rect 12216 1516 12265 1544
rect 12216 1504 12222 1516
rect 12253 1513 12265 1516
rect 12299 1513 12311 1547
rect 12253 1507 12311 1513
rect 12526 1504 12532 1556
rect 12584 1544 12590 1556
rect 12621 1547 12679 1553
rect 12621 1544 12633 1547
rect 12584 1516 12633 1544
rect 12584 1504 12590 1516
rect 12621 1513 12633 1516
rect 12667 1513 12679 1547
rect 12621 1507 12679 1513
rect 13078 1504 13084 1556
rect 13136 1544 13142 1556
rect 13173 1547 13231 1553
rect 13173 1544 13185 1547
rect 13136 1516 13185 1544
rect 13136 1504 13142 1516
rect 13173 1513 13185 1516
rect 13219 1513 13231 1547
rect 13173 1507 13231 1513
rect 13630 1504 13636 1556
rect 13688 1544 13694 1556
rect 13725 1547 13783 1553
rect 13725 1544 13737 1547
rect 13688 1516 13737 1544
rect 13688 1504 13694 1516
rect 13725 1513 13737 1516
rect 13771 1513 13783 1547
rect 13725 1507 13783 1513
rect 14182 1504 14188 1556
rect 14240 1544 14246 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 14240 1516 14289 1544
rect 14240 1504 14246 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 14734 1504 14740 1556
rect 14792 1544 14798 1556
rect 14829 1547 14887 1553
rect 14829 1544 14841 1547
rect 14792 1516 14841 1544
rect 14792 1504 14798 1516
rect 14829 1513 14841 1516
rect 14875 1513 14887 1547
rect 14829 1507 14887 1513
rect 15102 1504 15108 1556
rect 15160 1544 15166 1556
rect 15197 1547 15255 1553
rect 15197 1544 15209 1547
rect 15160 1516 15209 1544
rect 15160 1504 15166 1516
rect 15197 1513 15209 1516
rect 15243 1513 15255 1547
rect 15197 1507 15255 1513
rect 15654 1504 15660 1556
rect 15712 1544 15718 1556
rect 15841 1547 15899 1553
rect 15841 1544 15853 1547
rect 15712 1516 15853 1544
rect 15712 1504 15718 1516
rect 15841 1513 15853 1516
rect 15887 1513 15899 1547
rect 15841 1507 15899 1513
rect 16206 1504 16212 1556
rect 16264 1544 16270 1556
rect 16301 1547 16359 1553
rect 16301 1544 16313 1547
rect 16264 1516 16313 1544
rect 16264 1504 16270 1516
rect 16301 1513 16313 1516
rect 16347 1513 16359 1547
rect 16301 1507 16359 1513
rect 16758 1504 16764 1556
rect 16816 1544 16822 1556
rect 16853 1547 16911 1553
rect 16853 1544 16865 1547
rect 16816 1516 16865 1544
rect 16816 1504 16822 1516
rect 16853 1513 16865 1516
rect 16899 1513 16911 1547
rect 16853 1507 16911 1513
rect 17405 1547 17463 1553
rect 17405 1513 17417 1547
rect 17451 1544 17463 1547
rect 17494 1544 17500 1556
rect 17451 1516 17500 1544
rect 17451 1513 17463 1516
rect 17405 1507 17463 1513
rect 17494 1504 17500 1516
rect 17552 1504 17558 1556
rect 17586 1504 17592 1556
rect 17644 1544 17650 1556
rect 17773 1547 17831 1553
rect 17773 1544 17785 1547
rect 17644 1516 17785 1544
rect 17644 1504 17650 1516
rect 17773 1513 17785 1516
rect 17819 1544 17831 1547
rect 18138 1544 18144 1556
rect 17819 1516 18144 1544
rect 17819 1513 17831 1516
rect 17773 1507 17831 1513
rect 18138 1504 18144 1516
rect 18196 1504 18202 1556
rect 18230 1504 18236 1556
rect 18288 1544 18294 1556
rect 18325 1547 18383 1553
rect 18325 1544 18337 1547
rect 18288 1516 18337 1544
rect 18288 1504 18294 1516
rect 18325 1513 18337 1516
rect 18371 1513 18383 1547
rect 18325 1507 18383 1513
rect 18414 1504 18420 1556
rect 18472 1544 18478 1556
rect 19153 1547 19211 1553
rect 19153 1544 19165 1547
rect 18472 1516 19165 1544
rect 18472 1504 18478 1516
rect 19153 1513 19165 1516
rect 19199 1513 19211 1547
rect 19153 1507 19211 1513
rect 19334 1504 19340 1556
rect 19392 1504 19398 1556
rect 2225 1411 2283 1417
rect 2225 1377 2237 1411
rect 2271 1408 2283 1411
rect 2590 1408 2596 1420
rect 2271 1380 2596 1408
rect 2271 1377 2283 1380
rect 2225 1371 2283 1377
rect 2590 1368 2596 1380
rect 2648 1368 2654 1420
rect 2777 1411 2835 1417
rect 2777 1377 2789 1411
rect 2823 1408 2835 1411
rect 3160 1408 3188 1504
rect 8938 1436 8944 1488
rect 8996 1476 9002 1488
rect 9125 1479 9183 1485
rect 9125 1476 9137 1479
rect 8996 1448 9137 1476
rect 8996 1436 9002 1448
rect 9125 1445 9137 1448
rect 9171 1445 9183 1479
rect 9125 1439 9183 1445
rect 10410 1436 10416 1488
rect 10468 1476 10474 1488
rect 10965 1479 11023 1485
rect 10965 1476 10977 1479
rect 10468 1448 10977 1476
rect 10468 1436 10474 1448
rect 10965 1445 10977 1448
rect 11011 1445 11023 1479
rect 10965 1439 11023 1445
rect 13354 1436 13360 1488
rect 13412 1476 13418 1488
rect 14001 1479 14059 1485
rect 14001 1476 14013 1479
rect 13412 1448 14013 1476
rect 13412 1436 13418 1448
rect 14001 1445 14013 1448
rect 14047 1445 14059 1479
rect 14001 1439 14059 1445
rect 15746 1436 15752 1488
rect 15804 1476 15810 1488
rect 16117 1479 16175 1485
rect 16117 1476 16129 1479
rect 15804 1448 16129 1476
rect 15804 1436 15810 1448
rect 16117 1445 16129 1448
rect 16163 1445 16175 1479
rect 16117 1439 16175 1445
rect 16574 1436 16580 1488
rect 16632 1476 16638 1488
rect 18601 1479 18659 1485
rect 18601 1476 18613 1479
rect 16632 1448 18613 1476
rect 16632 1436 16638 1448
rect 18601 1445 18613 1448
rect 18647 1445 18659 1479
rect 18601 1439 18659 1445
rect 2823 1380 3188 1408
rect 3697 1411 3755 1417
rect 2823 1377 2835 1380
rect 2777 1371 2835 1377
rect 3697 1377 3709 1411
rect 3743 1408 3755 1411
rect 4062 1408 4068 1420
rect 3743 1380 4068 1408
rect 3743 1377 3755 1380
rect 3697 1371 3755 1377
rect 4062 1368 4068 1380
rect 4120 1368 4126 1420
rect 5718 1368 5724 1420
rect 5776 1408 5782 1420
rect 5813 1411 5871 1417
rect 5813 1408 5825 1411
rect 5776 1380 5825 1408
rect 5776 1368 5782 1380
rect 5813 1377 5825 1380
rect 5859 1377 5871 1411
rect 5813 1371 5871 1377
rect 6270 1368 6276 1420
rect 6328 1408 6334 1420
rect 6365 1411 6423 1417
rect 6365 1408 6377 1411
rect 6328 1380 6377 1408
rect 6328 1368 6334 1380
rect 6365 1377 6377 1380
rect 6411 1377 6423 1411
rect 6365 1371 6423 1377
rect 14274 1368 14280 1420
rect 14332 1408 14338 1420
rect 14332 1380 15516 1408
rect 14332 1368 14338 1380
rect 10962 1300 10968 1352
rect 11020 1340 11026 1352
rect 11241 1343 11299 1349
rect 11241 1340 11253 1343
rect 11020 1312 11253 1340
rect 11020 1300 11026 1312
rect 11241 1309 11253 1312
rect 11287 1309 11299 1343
rect 11241 1303 11299 1309
rect 11790 1300 11796 1352
rect 11848 1340 11854 1352
rect 12897 1343 12955 1349
rect 12897 1340 12909 1343
rect 11848 1312 12909 1340
rect 11848 1300 11854 1312
rect 12897 1309 12909 1312
rect 12943 1309 12955 1343
rect 12897 1303 12955 1309
rect 13538 1300 13544 1352
rect 13596 1340 13602 1352
rect 15488 1349 15516 1380
rect 18322 1368 18328 1420
rect 18380 1408 18386 1420
rect 18969 1411 19027 1417
rect 18969 1408 18981 1411
rect 18380 1380 18981 1408
rect 18380 1368 18386 1380
rect 18969 1377 18981 1380
rect 19015 1377 19027 1411
rect 18969 1371 19027 1377
rect 14553 1343 14611 1349
rect 14553 1340 14565 1343
rect 13596 1312 14565 1340
rect 13596 1300 13602 1312
rect 14553 1309 14565 1312
rect 14599 1309 14611 1343
rect 14553 1303 14611 1309
rect 15473 1343 15531 1349
rect 15473 1309 15485 1343
rect 15519 1309 15531 1343
rect 15473 1303 15531 1309
rect 16114 1300 16120 1352
rect 16172 1340 16178 1352
rect 17129 1343 17187 1349
rect 17129 1340 17141 1343
rect 16172 1312 17141 1340
rect 16172 1300 16178 1312
rect 17129 1309 17141 1312
rect 17175 1309 17187 1343
rect 17129 1303 17187 1309
rect 18782 1300 18788 1352
rect 18840 1300 18846 1352
rect 6825 1275 6883 1281
rect 6825 1241 6837 1275
rect 6871 1272 6883 1275
rect 7190 1272 7196 1284
rect 6871 1244 7196 1272
rect 6871 1241 6883 1244
rect 6825 1235 6883 1241
rect 7190 1232 7196 1244
rect 7248 1232 7254 1284
rect 12250 1232 12256 1284
rect 12308 1272 12314 1284
rect 13449 1275 13507 1281
rect 13449 1272 13461 1275
rect 12308 1244 13461 1272
rect 12308 1232 12314 1244
rect 13449 1241 13461 1244
rect 13495 1241 13507 1275
rect 13449 1235 13507 1241
rect 15286 1232 15292 1284
rect 15344 1272 15350 1284
rect 16577 1275 16635 1281
rect 16577 1272 16589 1275
rect 15344 1244 16589 1272
rect 15344 1232 15350 1244
rect 16577 1241 16589 1244
rect 16623 1241 16635 1275
rect 16577 1235 16635 1241
rect 16850 1232 16856 1284
rect 16908 1272 16914 1284
rect 18049 1275 18107 1281
rect 18049 1272 18061 1275
rect 16908 1244 18061 1272
rect 16908 1232 16914 1244
rect 18049 1241 18061 1244
rect 18095 1241 18107 1275
rect 18049 1235 18107 1241
rect 9582 1204 9588 1216
rect 9541 1176 9588 1204
rect 9582 1164 9588 1176
rect 9640 1204 9646 1216
rect 9677 1207 9735 1213
rect 9677 1204 9689 1207
rect 9640 1176 9689 1204
rect 9640 1164 9646 1176
rect 9677 1173 9689 1176
rect 9723 1173 9735 1207
rect 9677 1167 9735 1173
rect 276 1114 19780 1136
rect 276 1062 1122 1114
rect 1174 1062 1186 1114
rect 1238 1062 1250 1114
rect 1302 1062 1314 1114
rect 1366 1062 1378 1114
rect 1430 1062 9122 1114
rect 9174 1062 9186 1114
rect 9238 1062 9250 1114
rect 9302 1062 9314 1114
rect 9366 1062 9378 1114
rect 9430 1062 17122 1114
rect 17174 1062 17186 1114
rect 17238 1062 17250 1114
rect 17302 1062 17314 1114
rect 17366 1062 17378 1114
rect 17430 1062 19780 1114
rect 276 1040 19780 1062
rect 2222 960 2228 1012
rect 2280 1000 2286 1012
rect 2501 1003 2559 1009
rect 2501 1000 2513 1003
rect 2280 972 2513 1000
rect 2280 960 2286 972
rect 2501 969 2513 972
rect 2547 969 2559 1003
rect 2501 963 2559 969
rect 2774 960 2780 1012
rect 2832 960 2838 1012
rect 2958 960 2964 1012
rect 3016 960 3022 1012
rect 3326 960 3332 1012
rect 3384 960 3390 1012
rect 3510 960 3516 1012
rect 3568 960 3574 1012
rect 3878 960 3884 1012
rect 3936 960 3942 1012
rect 4246 960 4252 1012
rect 4304 960 4310 1012
rect 4430 960 4436 1012
rect 4488 960 4494 1012
rect 4614 960 4620 1012
rect 4672 960 4678 1012
rect 4801 1003 4859 1009
rect 4801 969 4813 1003
rect 4847 1000 4859 1003
rect 4982 1000 4988 1012
rect 4847 972 4988 1000
rect 4847 969 4859 972
rect 4801 963 4859 969
rect 4982 960 4988 972
rect 5040 960 5046 1012
rect 5261 1003 5319 1009
rect 5261 969 5273 1003
rect 5307 1000 5319 1003
rect 5350 1000 5356 1012
rect 5307 972 5356 1000
rect 5307 969 5319 972
rect 5261 963 5319 969
rect 5350 960 5356 972
rect 5408 960 5414 1012
rect 5534 960 5540 1012
rect 5592 960 5598 1012
rect 5902 960 5908 1012
rect 5960 960 5966 1012
rect 6454 960 6460 1012
rect 6512 960 6518 1012
rect 7006 960 7012 1012
rect 7064 960 7070 1012
rect 7558 960 7564 1012
rect 7616 960 7622 1012
rect 8202 960 8208 1012
rect 8260 960 8266 1012
rect 8662 960 8668 1012
rect 8720 960 8726 1012
rect 8938 960 8944 1012
rect 8996 1000 9002 1012
rect 9401 1003 9459 1009
rect 9401 1000 9413 1003
rect 8996 972 9413 1000
rect 8996 960 9002 972
rect 9401 969 9413 972
rect 9447 969 9459 1003
rect 9401 963 9459 969
rect 11606 960 11612 1012
rect 11664 1000 11670 1012
rect 11977 1003 12035 1009
rect 11977 1000 11989 1003
rect 11664 972 11989 1000
rect 11664 960 11670 972
rect 11977 969 11989 972
rect 12023 969 12035 1003
rect 11977 963 12035 969
rect 12158 960 12164 1012
rect 12216 1000 12222 1012
rect 12529 1003 12587 1009
rect 12529 1000 12541 1003
rect 12216 972 12541 1000
rect 12216 960 12222 972
rect 12529 969 12541 972
rect 12575 969 12587 1003
rect 12529 963 12587 969
rect 12894 960 12900 1012
rect 12952 960 12958 1012
rect 13078 960 13084 1012
rect 13136 1000 13142 1012
rect 13817 1003 13875 1009
rect 13817 1000 13829 1003
rect 13136 972 13829 1000
rect 13136 960 13142 972
rect 13817 969 13829 972
rect 13863 969 13875 1003
rect 13817 963 13875 969
rect 14090 960 14096 1012
rect 14148 960 14154 1012
rect 14182 960 14188 1012
rect 14240 1000 14246 1012
rect 14737 1003 14795 1009
rect 14737 1000 14749 1003
rect 14240 972 14749 1000
rect 14240 960 14246 972
rect 14737 969 14749 972
rect 14783 969 14795 1003
rect 14737 963 14795 969
rect 14918 960 14924 1012
rect 14976 960 14982 1012
rect 15194 960 15200 1012
rect 15252 1000 15258 1012
rect 15565 1003 15623 1009
rect 15565 1000 15577 1003
rect 15252 972 15577 1000
rect 15252 960 15258 972
rect 15565 969 15577 972
rect 15611 969 15623 1003
rect 15565 963 15623 969
rect 15654 960 15660 1012
rect 15712 1000 15718 1012
rect 16301 1003 16359 1009
rect 16301 1000 16313 1003
rect 15712 972 16313 1000
rect 15712 960 15718 972
rect 16301 969 16313 972
rect 16347 969 16359 1003
rect 16301 963 16359 969
rect 16390 960 16396 1012
rect 16448 1000 16454 1012
rect 16669 1003 16727 1009
rect 16669 1000 16681 1003
rect 16448 972 16681 1000
rect 16448 960 16454 972
rect 16669 969 16681 972
rect 16715 969 16727 1003
rect 16669 963 16727 969
rect 16758 960 16764 1012
rect 16816 1000 16822 1012
rect 17313 1003 17371 1009
rect 17313 1000 17325 1003
rect 16816 972 17325 1000
rect 16816 960 16822 972
rect 17313 969 17325 972
rect 17359 969 17371 1003
rect 17313 963 17371 969
rect 17494 960 17500 1012
rect 17552 1000 17558 1012
rect 17681 1003 17739 1009
rect 17681 1000 17693 1003
rect 17552 972 17693 1000
rect 17552 960 17558 972
rect 17681 969 17693 972
rect 17727 969 17739 1003
rect 17681 963 17739 969
rect 18138 960 18144 1012
rect 18196 960 18202 1012
rect 18230 960 18236 1012
rect 18288 1000 18294 1012
rect 18601 1003 18659 1009
rect 18601 1000 18613 1003
rect 18288 972 18613 1000
rect 18288 960 18294 972
rect 18601 969 18613 972
rect 18647 969 18659 1003
rect 18601 963 18659 969
rect 18966 960 18972 1012
rect 19024 1000 19030 1012
rect 19245 1003 19303 1009
rect 19245 1000 19257 1003
rect 19024 972 19257 1000
rect 19024 960 19030 972
rect 19245 969 19257 972
rect 19291 969 19303 1003
rect 19245 963 19303 969
rect 3694 892 3700 944
rect 3752 932 3758 944
rect 3973 935 4031 941
rect 3973 932 3985 935
rect 3752 904 3985 932
rect 3752 892 3758 904
rect 3973 901 3985 904
rect 4019 901 4031 935
rect 3973 895 4031 901
rect 5718 892 5724 944
rect 5776 932 5782 944
rect 6089 935 6147 941
rect 6089 932 6101 935
rect 5776 904 6101 932
rect 5776 892 5782 904
rect 6089 901 6101 904
rect 6135 901 6147 935
rect 6089 895 6147 901
rect 6270 892 6276 944
rect 6328 932 6334 944
rect 6641 935 6699 941
rect 6641 932 6653 935
rect 6328 904 6653 932
rect 6328 892 6334 904
rect 6641 901 6653 904
rect 6687 901 6699 935
rect 6641 895 6699 901
rect 6914 892 6920 944
rect 6972 932 6978 944
rect 7193 935 7251 941
rect 7193 932 7205 935
rect 6972 904 7205 932
rect 6972 892 6978 904
rect 7193 901 7205 904
rect 7239 901 7251 935
rect 7193 895 7251 901
rect 7374 892 7380 944
rect 7432 932 7438 944
rect 7745 935 7803 941
rect 7745 932 7757 935
rect 7432 904 7757 932
rect 7432 892 7438 904
rect 7745 901 7757 904
rect 7791 901 7803 935
rect 7745 895 7803 901
rect 8478 892 8484 944
rect 8536 932 8542 944
rect 8849 935 8907 941
rect 8849 932 8861 935
rect 8536 904 8861 932
rect 8536 892 8542 904
rect 8849 901 8861 904
rect 8895 901 8907 935
rect 8849 895 8907 901
rect 12066 892 12072 944
rect 12124 932 12130 944
rect 12437 935 12495 941
rect 12437 932 12449 935
rect 12124 904 12449 932
rect 12124 892 12130 904
rect 12437 901 12449 904
rect 12483 901 12495 935
rect 12437 895 12495 901
rect 13446 892 13452 944
rect 13504 932 13510 944
rect 13541 935 13599 941
rect 13541 932 13553 935
rect 13504 904 13553 932
rect 13504 892 13510 904
rect 13541 901 13553 904
rect 13587 901 13599 935
rect 13541 895 13599 901
rect 13630 892 13636 944
rect 13688 932 13694 944
rect 14553 935 14611 941
rect 14553 932 14565 935
rect 13688 904 14565 932
rect 13688 892 13694 904
rect 14553 901 14565 904
rect 14599 901 14611 935
rect 14553 895 14611 901
rect 14826 892 14832 944
rect 14884 932 14890 944
rect 15289 935 15347 941
rect 15289 932 15301 935
rect 14884 904 15301 932
rect 14884 892 14890 904
rect 15289 901 15301 904
rect 15335 901 15347 935
rect 15289 895 15347 901
rect 15838 892 15844 944
rect 15896 932 15902 944
rect 16117 935 16175 941
rect 16117 932 16129 935
rect 15896 904 16129 932
rect 15896 892 15902 904
rect 16117 901 16129 904
rect 16163 901 16175 935
rect 16117 895 16175 901
rect 16206 892 16212 944
rect 16264 932 16270 944
rect 17129 935 17187 941
rect 17129 932 17141 935
rect 16264 904 17141 932
rect 16264 892 16270 904
rect 17129 901 17141 904
rect 17175 901 17187 935
rect 17129 895 17187 901
rect 4985 867 5043 873
rect 4985 833 4997 867
rect 5031 864 5043 867
rect 5166 864 5172 876
rect 5031 836 5172 864
rect 5031 833 5043 836
rect 4985 827 5043 833
rect 5166 824 5172 836
rect 5224 824 5230 876
rect 8110 824 8116 876
rect 8168 864 8174 876
rect 9033 867 9091 873
rect 9033 864 9045 867
rect 8168 836 9045 864
rect 8168 824 8174 836
rect 9033 833 9045 836
rect 9079 833 9091 867
rect 9033 827 9091 833
rect 12526 824 12532 876
rect 12584 864 12590 876
rect 13265 867 13323 873
rect 13265 864 13277 867
rect 12584 836 13277 864
rect 12584 824 12590 836
rect 13265 833 13277 836
rect 13311 833 13323 867
rect 13265 827 13323 833
rect 14366 824 14372 876
rect 14424 824 14430 876
rect 14734 824 14740 876
rect 14792 864 14798 876
rect 15381 867 15439 873
rect 15381 864 15393 867
rect 14792 836 15393 864
rect 14792 824 14798 836
rect 15381 833 15393 836
rect 15427 833 15439 867
rect 15381 827 15439 833
rect 16942 824 16948 876
rect 17000 824 17006 876
rect 7742 756 7748 808
rect 7800 796 7806 808
rect 8297 799 8355 805
rect 8297 796 8309 799
rect 7800 768 8309 796
rect 7800 756 7806 768
rect 8297 765 8309 768
rect 8343 765 8355 799
rect 8297 759 8355 765
rect 276 570 19780 592
rect 276 518 1762 570
rect 1814 518 1826 570
rect 1878 518 1890 570
rect 1942 518 1954 570
rect 2006 518 2018 570
rect 2070 518 9762 570
rect 9814 518 9826 570
rect 9878 518 9890 570
rect 9942 518 9954 570
rect 10006 518 10018 570
rect 10070 518 17762 570
rect 17814 518 17826 570
rect 17878 518 17890 570
rect 17942 518 17954 570
rect 18006 518 18018 570
rect 18070 518 19780 570
rect 276 496 19780 518
<< via1 >>
rect 18052 2456 18104 2508
rect 18972 2456 19024 2508
rect 1584 2320 1636 2372
rect 1860 2320 1912 2372
rect 17132 2320 17184 2372
rect 18328 2320 18380 2372
rect 1122 2150 1174 2202
rect 1186 2150 1238 2202
rect 1250 2150 1302 2202
rect 1314 2150 1366 2202
rect 1378 2150 1430 2202
rect 9122 2150 9174 2202
rect 9186 2150 9238 2202
rect 9250 2150 9302 2202
rect 9314 2150 9366 2202
rect 9378 2150 9430 2202
rect 17122 2150 17174 2202
rect 17186 2150 17238 2202
rect 17250 2150 17302 2202
rect 17314 2150 17366 2202
rect 17378 2150 17430 2202
rect 13452 2048 13504 2100
rect 14280 2048 14332 2100
rect 14556 2048 14608 2100
rect 15200 2048 15252 2100
rect 16948 2048 17000 2100
rect 1584 1912 1636 1964
rect 2136 1912 2188 1964
rect 2596 1912 2648 1964
rect 2964 1912 3016 1964
rect 3332 1912 3384 1964
rect 3516 1912 3568 1964
rect 3884 1912 3936 1964
rect 4436 1912 4488 1964
rect 5172 1912 5224 1964
rect 5540 1912 5592 1964
rect 5908 1912 5960 1964
rect 6460 1912 6512 1964
rect 7012 1912 7064 1964
rect 7564 1912 7616 1964
rect 8300 1912 8352 1964
rect 8668 1912 8720 1964
rect 11244 1980 11296 2032
rect 12716 1980 12768 2032
rect 13544 1980 13596 2032
rect 16396 1980 16448 2032
rect 8852 1912 8904 1964
rect 9036 1955 9088 1964
rect 9036 1921 9045 1955
rect 9045 1921 9079 1955
rect 9079 1921 9088 1955
rect 9036 1912 9088 1921
rect 9496 1912 9548 1964
rect 9588 1955 9640 1964
rect 9588 1921 9597 1955
rect 9597 1921 9631 1955
rect 9631 1921 9640 1955
rect 9588 1912 9640 1921
rect 10140 1912 10192 1964
rect 10416 1912 10468 1964
rect 10876 1912 10928 1964
rect 11980 1912 12032 1964
rect 12072 1955 12124 1964
rect 12072 1921 12081 1955
rect 12081 1921 12115 1955
rect 12115 1921 12124 1955
rect 12072 1912 12124 1921
rect 13268 1912 13320 1964
rect 14372 1912 14424 1964
rect 14464 1912 14516 1964
rect 15752 1912 15804 1964
rect 15844 1912 15896 1964
rect 16948 1912 17000 1964
rect 18788 1980 18840 2032
rect 2412 1844 2464 1896
rect 4068 1844 4120 1896
rect 6092 1844 6144 1896
rect 6644 1844 6696 1896
rect 7196 1844 7248 1896
rect 10232 1844 10284 1896
rect 10508 1844 10560 1896
rect 10968 1887 11020 1896
rect 10968 1853 10977 1887
rect 10977 1853 11011 1887
rect 11011 1853 11020 1887
rect 10968 1844 11020 1853
rect 11796 1844 11848 1896
rect 12900 1844 12952 1896
rect 12992 1844 13044 1896
rect 4160 1776 4212 1828
rect 4804 1776 4856 1828
rect 5356 1776 5408 1828
rect 7288 1776 7340 1828
rect 7932 1776 7984 1828
rect 10692 1776 10744 1828
rect 11244 1819 11296 1828
rect 11244 1785 11253 1819
rect 11253 1785 11287 1819
rect 11287 1785 11296 1819
rect 11244 1776 11296 1785
rect 11428 1776 11480 1828
rect 12256 1776 12308 1828
rect 12440 1776 12492 1828
rect 13452 1776 13504 1828
rect 13544 1819 13596 1828
rect 13544 1785 13553 1819
rect 13553 1785 13587 1819
rect 13587 1785 13596 1819
rect 13544 1776 13596 1785
rect 10324 1708 10376 1760
rect 11060 1708 11112 1760
rect 11796 1751 11848 1760
rect 11796 1717 11805 1751
rect 11805 1717 11839 1751
rect 11839 1717 11848 1751
rect 11796 1708 11848 1717
rect 11888 1708 11940 1760
rect 13360 1708 13412 1760
rect 13820 1844 13872 1896
rect 14924 1844 14976 1896
rect 15476 1844 15528 1896
rect 16396 1887 16448 1896
rect 16396 1853 16405 1887
rect 16405 1853 16439 1887
rect 16439 1853 16448 1887
rect 16396 1844 16448 1853
rect 14004 1776 14056 1828
rect 14832 1776 14884 1828
rect 14096 1708 14148 1760
rect 14280 1708 14332 1760
rect 15016 1776 15068 1828
rect 15844 1819 15896 1828
rect 15844 1785 15853 1819
rect 15853 1785 15887 1819
rect 15887 1785 15896 1819
rect 15844 1776 15896 1785
rect 16028 1776 16080 1828
rect 15200 1708 15252 1760
rect 15568 1708 15620 1760
rect 16120 1751 16172 1760
rect 16120 1717 16129 1751
rect 16129 1717 16163 1751
rect 16163 1717 16172 1751
rect 16120 1708 16172 1717
rect 16580 1776 16632 1828
rect 18144 1912 18196 1964
rect 19340 1912 19392 1964
rect 17592 1844 17644 1896
rect 18420 1887 18472 1896
rect 18420 1853 18429 1887
rect 18429 1853 18463 1887
rect 18463 1853 18472 1887
rect 18420 1844 18472 1853
rect 18972 1887 19024 1896
rect 18972 1853 18981 1887
rect 18981 1853 19015 1887
rect 19015 1853 19024 1887
rect 18972 1844 19024 1853
rect 16856 1708 16908 1760
rect 18328 1776 18380 1828
rect 1762 1606 1814 1658
rect 1826 1606 1878 1658
rect 1890 1606 1942 1658
rect 1954 1606 2006 1658
rect 2018 1606 2070 1658
rect 9762 1606 9814 1658
rect 9826 1606 9878 1658
rect 9890 1606 9942 1658
rect 9954 1606 10006 1658
rect 10018 1606 10070 1658
rect 17762 1606 17814 1658
rect 17826 1606 17878 1658
rect 17890 1606 17942 1658
rect 17954 1606 18006 1658
rect 18018 1606 18070 1658
rect 1676 1547 1728 1556
rect 1676 1513 1685 1547
rect 1685 1513 1719 1547
rect 1719 1513 1728 1547
rect 1676 1504 1728 1513
rect 2228 1504 2280 1556
rect 2780 1504 2832 1556
rect 3148 1504 3200 1556
rect 3700 1504 3752 1556
rect 4160 1547 4212 1556
rect 4160 1513 4169 1547
rect 4169 1513 4203 1547
rect 4203 1513 4212 1547
rect 4160 1504 4212 1513
rect 4252 1504 4304 1556
rect 4620 1504 4672 1556
rect 4988 1504 5040 1556
rect 6092 1504 6144 1556
rect 6644 1504 6696 1556
rect 6828 1504 6880 1556
rect 7288 1547 7340 1556
rect 7288 1513 7297 1547
rect 7297 1513 7331 1547
rect 7331 1513 7340 1547
rect 7288 1504 7340 1513
rect 7380 1504 7432 1556
rect 7748 1504 7800 1556
rect 8116 1504 8168 1556
rect 8484 1504 8536 1556
rect 9036 1547 9088 1556
rect 9036 1513 9045 1547
rect 9045 1513 9079 1547
rect 9079 1513 9088 1547
rect 9036 1504 9088 1513
rect 9496 1547 9548 1556
rect 9496 1513 9505 1547
rect 9505 1513 9539 1547
rect 9539 1513 9548 1547
rect 9496 1504 9548 1513
rect 10140 1504 10192 1556
rect 10232 1547 10284 1556
rect 10232 1513 10241 1547
rect 10241 1513 10275 1547
rect 10275 1513 10284 1547
rect 10232 1504 10284 1513
rect 10324 1504 10376 1556
rect 11244 1504 11296 1556
rect 11612 1504 11664 1556
rect 11980 1547 12032 1556
rect 11980 1513 11989 1547
rect 11989 1513 12023 1547
rect 12023 1513 12032 1547
rect 11980 1504 12032 1513
rect 12164 1504 12216 1556
rect 12532 1504 12584 1556
rect 13084 1504 13136 1556
rect 13636 1504 13688 1556
rect 14188 1504 14240 1556
rect 14740 1504 14792 1556
rect 15108 1504 15160 1556
rect 15660 1504 15712 1556
rect 16212 1504 16264 1556
rect 16764 1504 16816 1556
rect 17500 1504 17552 1556
rect 17592 1504 17644 1556
rect 18144 1504 18196 1556
rect 18236 1504 18288 1556
rect 18420 1504 18472 1556
rect 19340 1547 19392 1556
rect 19340 1513 19349 1547
rect 19349 1513 19383 1547
rect 19383 1513 19392 1547
rect 19340 1504 19392 1513
rect 2596 1368 2648 1420
rect 8944 1436 8996 1488
rect 10416 1436 10468 1488
rect 13360 1436 13412 1488
rect 15752 1436 15804 1488
rect 16580 1436 16632 1488
rect 4068 1368 4120 1420
rect 5724 1368 5776 1420
rect 6276 1368 6328 1420
rect 14280 1368 14332 1420
rect 10968 1300 11020 1352
rect 11796 1300 11848 1352
rect 13544 1300 13596 1352
rect 18328 1368 18380 1420
rect 16120 1300 16172 1352
rect 18788 1343 18840 1352
rect 18788 1309 18797 1343
rect 18797 1309 18831 1343
rect 18831 1309 18840 1343
rect 18788 1300 18840 1309
rect 7196 1232 7248 1284
rect 12256 1232 12308 1284
rect 15292 1232 15344 1284
rect 16856 1232 16908 1284
rect 9588 1164 9640 1216
rect 1122 1062 1174 1114
rect 1186 1062 1238 1114
rect 1250 1062 1302 1114
rect 1314 1062 1366 1114
rect 1378 1062 1430 1114
rect 9122 1062 9174 1114
rect 9186 1062 9238 1114
rect 9250 1062 9302 1114
rect 9314 1062 9366 1114
rect 9378 1062 9430 1114
rect 17122 1062 17174 1114
rect 17186 1062 17238 1114
rect 17250 1062 17302 1114
rect 17314 1062 17366 1114
rect 17378 1062 17430 1114
rect 2228 960 2280 1012
rect 2780 1003 2832 1012
rect 2780 969 2789 1003
rect 2789 969 2823 1003
rect 2823 969 2832 1003
rect 2780 960 2832 969
rect 2964 1003 3016 1012
rect 2964 969 2973 1003
rect 2973 969 3007 1003
rect 3007 969 3016 1003
rect 2964 960 3016 969
rect 3332 1003 3384 1012
rect 3332 969 3341 1003
rect 3341 969 3375 1003
rect 3375 969 3384 1003
rect 3332 960 3384 969
rect 3516 1003 3568 1012
rect 3516 969 3525 1003
rect 3525 969 3559 1003
rect 3559 969 3568 1003
rect 3516 960 3568 969
rect 3884 1003 3936 1012
rect 3884 969 3893 1003
rect 3893 969 3927 1003
rect 3927 969 3936 1003
rect 3884 960 3936 969
rect 4252 1003 4304 1012
rect 4252 969 4261 1003
rect 4261 969 4295 1003
rect 4295 969 4304 1003
rect 4252 960 4304 969
rect 4436 1003 4488 1012
rect 4436 969 4445 1003
rect 4445 969 4479 1003
rect 4479 969 4488 1003
rect 4436 960 4488 969
rect 4620 1003 4672 1012
rect 4620 969 4629 1003
rect 4629 969 4663 1003
rect 4663 969 4672 1003
rect 4620 960 4672 969
rect 4988 960 5040 1012
rect 5356 960 5408 1012
rect 5540 1003 5592 1012
rect 5540 969 5549 1003
rect 5549 969 5583 1003
rect 5583 969 5592 1003
rect 5540 960 5592 969
rect 5908 1003 5960 1012
rect 5908 969 5917 1003
rect 5917 969 5951 1003
rect 5951 969 5960 1003
rect 5908 960 5960 969
rect 6460 1003 6512 1012
rect 6460 969 6469 1003
rect 6469 969 6503 1003
rect 6503 969 6512 1003
rect 6460 960 6512 969
rect 7012 1003 7064 1012
rect 7012 969 7021 1003
rect 7021 969 7055 1003
rect 7055 969 7064 1003
rect 7012 960 7064 969
rect 7564 1003 7616 1012
rect 7564 969 7573 1003
rect 7573 969 7607 1003
rect 7607 969 7616 1003
rect 7564 960 7616 969
rect 8208 1003 8260 1012
rect 8208 969 8217 1003
rect 8217 969 8251 1003
rect 8251 969 8260 1003
rect 8208 960 8260 969
rect 8668 1003 8720 1012
rect 8668 969 8677 1003
rect 8677 969 8711 1003
rect 8711 969 8720 1003
rect 8668 960 8720 969
rect 8944 960 8996 1012
rect 11612 960 11664 1012
rect 12164 960 12216 1012
rect 12900 1003 12952 1012
rect 12900 969 12909 1003
rect 12909 969 12943 1003
rect 12943 969 12952 1003
rect 12900 960 12952 969
rect 13084 960 13136 1012
rect 14096 1003 14148 1012
rect 14096 969 14105 1003
rect 14105 969 14139 1003
rect 14139 969 14148 1003
rect 14096 960 14148 969
rect 14188 960 14240 1012
rect 14924 1003 14976 1012
rect 14924 969 14933 1003
rect 14933 969 14967 1003
rect 14967 969 14976 1003
rect 14924 960 14976 969
rect 15200 960 15252 1012
rect 15660 960 15712 1012
rect 16396 960 16448 1012
rect 16764 960 16816 1012
rect 17500 960 17552 1012
rect 18144 1003 18196 1012
rect 18144 969 18153 1003
rect 18153 969 18187 1003
rect 18187 969 18196 1003
rect 18144 960 18196 969
rect 18236 960 18288 1012
rect 18972 960 19024 1012
rect 3700 892 3752 944
rect 5724 892 5776 944
rect 6276 892 6328 944
rect 6920 892 6972 944
rect 7380 892 7432 944
rect 8484 892 8536 944
rect 12072 892 12124 944
rect 13452 892 13504 944
rect 13636 892 13688 944
rect 14832 892 14884 944
rect 15844 892 15896 944
rect 16212 892 16264 944
rect 5172 824 5224 876
rect 8116 824 8168 876
rect 12532 824 12584 876
rect 14372 867 14424 876
rect 14372 833 14381 867
rect 14381 833 14415 867
rect 14415 833 14424 867
rect 14372 824 14424 833
rect 14740 824 14792 876
rect 16948 867 17000 876
rect 16948 833 16957 867
rect 16957 833 16991 867
rect 16991 833 17000 867
rect 16948 824 17000 833
rect 7748 756 7800 808
rect 1762 518 1814 570
rect 1826 518 1878 570
rect 1890 518 1942 570
rect 1954 518 2006 570
rect 2018 518 2070 570
rect 9762 518 9814 570
rect 9826 518 9878 570
rect 9890 518 9942 570
rect 9954 518 10006 570
rect 10018 518 10070 570
rect 17762 518 17814 570
rect 17826 518 17878 570
rect 17890 518 17942 570
rect 17954 518 18006 570
rect 18018 518 18070 570
<< metal2 >>
rect 1674 3000 1730 3400
rect 1858 3000 1914 3400
rect 2042 3000 2098 3400
rect 2226 3000 2282 3400
rect 2410 3000 2466 3400
rect 2594 3000 2650 3400
rect 2778 3000 2834 3400
rect 2962 3000 3018 3400
rect 3146 3000 3202 3400
rect 3330 3000 3386 3400
rect 3514 3000 3570 3400
rect 3698 3000 3754 3400
rect 3882 3000 3938 3400
rect 4066 3000 4122 3400
rect 4250 3000 4306 3400
rect 4434 3000 4490 3400
rect 4618 3000 4674 3400
rect 4802 3000 4858 3400
rect 4986 3000 5042 3400
rect 5170 3000 5226 3400
rect 5354 3000 5410 3400
rect 5538 3000 5594 3400
rect 5722 3000 5778 3400
rect 5906 3000 5962 3400
rect 6090 3000 6146 3400
rect 6274 3000 6330 3400
rect 6458 3000 6514 3400
rect 6642 3000 6698 3400
rect 6826 3000 6882 3400
rect 7010 3000 7066 3400
rect 7194 3000 7250 3400
rect 7378 3000 7434 3400
rect 7562 3000 7618 3400
rect 7746 3000 7802 3400
rect 7930 3000 7986 3400
rect 8114 3000 8170 3400
rect 8298 3000 8354 3400
rect 8482 3000 8538 3400
rect 8666 3000 8722 3400
rect 8850 3000 8906 3400
rect 9034 3000 9090 3400
rect 9218 3000 9274 3400
rect 9402 3000 9458 3400
rect 9586 3000 9642 3400
rect 9770 3000 9826 3400
rect 9954 3000 10010 3400
rect 10138 3000 10194 3400
rect 10322 3000 10378 3400
rect 10506 3000 10562 3400
rect 10690 3000 10746 3400
rect 10874 3000 10930 3400
rect 11058 3000 11114 3400
rect 11242 3000 11298 3400
rect 11426 3000 11482 3400
rect 11610 3000 11666 3400
rect 11794 3000 11850 3400
rect 11978 3000 12034 3400
rect 12162 3000 12218 3400
rect 12346 3000 12402 3400
rect 12530 3000 12586 3400
rect 12714 3000 12770 3400
rect 12898 3000 12954 3400
rect 13082 3000 13138 3400
rect 13266 3000 13322 3400
rect 13450 3000 13506 3400
rect 13634 3000 13690 3400
rect 13818 3000 13874 3400
rect 14002 3000 14058 3400
rect 14186 3000 14242 3400
rect 14370 3000 14426 3400
rect 14554 3000 14610 3400
rect 14738 3000 14794 3400
rect 14922 3000 14978 3400
rect 15106 3000 15162 3400
rect 15290 3000 15346 3400
rect 15474 3000 15530 3400
rect 15658 3000 15714 3400
rect 15842 3000 15898 3400
rect 16026 3000 16082 3400
rect 16210 3000 16266 3400
rect 16394 3000 16450 3400
rect 16578 3000 16634 3400
rect 16762 3000 16818 3400
rect 16946 3000 17002 3400
rect 17130 3000 17186 3400
rect 17314 3000 17370 3400
rect 17498 3000 17554 3400
rect 17682 3000 17738 3400
rect 17866 3000 17922 3400
rect 18050 3000 18106 3400
rect 18234 3000 18290 3400
rect 1584 2372 1636 2378
rect 1584 2314 1636 2320
rect 1116 2202 1436 2224
rect 1116 2150 1122 2202
rect 1174 2150 1186 2202
rect 1238 2150 1250 2202
rect 1302 2150 1314 2202
rect 1366 2150 1378 2202
rect 1430 2150 1436 2202
rect 1116 1188 1436 2150
rect 1596 1970 1624 2314
rect 1584 1964 1636 1970
rect 1584 1906 1636 1912
rect 1688 1562 1716 3000
rect 1872 2378 1900 3000
rect 2056 2394 2084 3000
rect 1860 2372 1912 2378
rect 2056 2366 2176 2394
rect 1860 2314 1912 2320
rect 1756 1828 2076 2224
rect 2148 1970 2176 2366
rect 2136 1964 2188 1970
rect 2136 1906 2188 1912
rect 1756 1772 1768 1828
rect 1824 1772 1848 1828
rect 1904 1772 1928 1828
rect 1984 1772 2008 1828
rect 2064 1772 2076 1828
rect 1756 1748 2076 1772
rect 1756 1692 1768 1748
rect 1824 1692 1848 1748
rect 1904 1692 1928 1748
rect 1984 1692 2008 1748
rect 2064 1692 2076 1748
rect 1756 1668 2076 1692
rect 1756 1658 1768 1668
rect 1824 1658 1848 1668
rect 1904 1658 1928 1668
rect 1984 1658 2008 1668
rect 2064 1658 2076 1668
rect 1756 1606 1762 1658
rect 1824 1612 1826 1658
rect 2006 1612 2008 1658
rect 1814 1606 1826 1612
rect 1878 1606 1890 1612
rect 1942 1606 1954 1612
rect 2006 1606 2018 1612
rect 2070 1606 2076 1658
rect 1756 1588 2076 1606
rect 1676 1556 1728 1562
rect 1676 1498 1728 1504
rect 1756 1532 1768 1588
rect 1824 1532 1848 1588
rect 1904 1532 1928 1588
rect 1984 1532 2008 1588
rect 2064 1532 2076 1588
rect 2240 1562 2268 3000
rect 2424 1902 2452 3000
rect 2608 1970 2636 3000
rect 2596 1964 2648 1970
rect 2596 1906 2648 1912
rect 2412 1896 2464 1902
rect 2412 1838 2464 1844
rect 1116 1132 1128 1188
rect 1184 1132 1208 1188
rect 1264 1132 1288 1188
rect 1344 1132 1368 1188
rect 1424 1132 1436 1188
rect 1116 1114 1436 1132
rect 1116 1062 1122 1114
rect 1174 1108 1186 1114
rect 1238 1108 1250 1114
rect 1302 1108 1314 1114
rect 1366 1108 1378 1114
rect 1184 1062 1186 1108
rect 1366 1062 1368 1108
rect 1430 1062 1436 1114
rect 1116 1052 1128 1062
rect 1184 1052 1208 1062
rect 1264 1052 1288 1062
rect 1344 1052 1368 1062
rect 1424 1052 1436 1062
rect 1116 1028 1436 1052
rect 1116 972 1128 1028
rect 1184 972 1208 1028
rect 1264 972 1288 1028
rect 1344 972 1368 1028
rect 1424 972 1436 1028
rect 1116 948 1436 972
rect 1116 892 1128 948
rect 1184 892 1208 948
rect 1264 892 1288 948
rect 1344 892 1368 948
rect 1424 892 1436 948
rect 1116 496 1436 892
rect 1756 570 2076 1532
rect 2228 1556 2280 1562
rect 2228 1498 2280 1504
rect 2240 1018 2268 1498
rect 2608 1426 2636 1906
rect 2792 1562 2820 3000
rect 2976 1970 3004 3000
rect 2964 1964 3016 1970
rect 2964 1906 3016 1912
rect 2780 1556 2832 1562
rect 2780 1498 2832 1504
rect 2596 1420 2648 1426
rect 2596 1362 2648 1368
rect 2792 1018 2820 1498
rect 2976 1018 3004 1906
rect 3160 1562 3188 3000
rect 3344 1970 3372 3000
rect 3528 1970 3556 3000
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3516 1964 3568 1970
rect 3516 1906 3568 1912
rect 3148 1556 3200 1562
rect 3148 1498 3200 1504
rect 3344 1018 3372 1906
rect 3528 1018 3556 1906
rect 3712 1562 3740 3000
rect 3896 1970 3924 3000
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 3700 1556 3752 1562
rect 3700 1498 3752 1504
rect 2228 1012 2280 1018
rect 2228 954 2280 960
rect 2780 1012 2832 1018
rect 2780 954 2832 960
rect 2964 1012 3016 1018
rect 2964 954 3016 960
rect 3332 1012 3384 1018
rect 3332 954 3384 960
rect 3516 1012 3568 1018
rect 3516 954 3568 960
rect 3712 950 3740 1498
rect 3896 1018 3924 1906
rect 4080 1902 4108 3000
rect 4068 1896 4120 1902
rect 4068 1838 4120 1844
rect 4080 1426 4108 1838
rect 4160 1828 4212 1834
rect 4160 1770 4212 1776
rect 4172 1562 4200 1770
rect 4264 1562 4292 3000
rect 4448 1970 4476 3000
rect 4436 1964 4488 1970
rect 4436 1906 4488 1912
rect 4160 1556 4212 1562
rect 4160 1498 4212 1504
rect 4252 1556 4304 1562
rect 4252 1498 4304 1504
rect 4068 1420 4120 1426
rect 4068 1362 4120 1368
rect 4264 1018 4292 1498
rect 4448 1018 4476 1906
rect 4632 1562 4660 3000
rect 4816 1834 4844 3000
rect 4804 1828 4856 1834
rect 4804 1770 4856 1776
rect 5000 1562 5028 3000
rect 5184 1970 5212 3000
rect 5172 1964 5224 1970
rect 5172 1906 5224 1912
rect 4620 1556 4672 1562
rect 4620 1498 4672 1504
rect 4988 1556 5040 1562
rect 4988 1498 5040 1504
rect 4632 1018 4660 1498
rect 5000 1018 5028 1498
rect 3884 1012 3936 1018
rect 3884 954 3936 960
rect 4252 1012 4304 1018
rect 4252 954 4304 960
rect 4436 1012 4488 1018
rect 4436 954 4488 960
rect 4620 1012 4672 1018
rect 4620 954 4672 960
rect 4988 1012 5040 1018
rect 4988 954 5040 960
rect 3700 944 3752 950
rect 3700 886 3752 892
rect 5184 882 5212 1906
rect 5368 1834 5396 3000
rect 5552 1970 5580 3000
rect 5540 1964 5592 1970
rect 5540 1906 5592 1912
rect 5356 1828 5408 1834
rect 5356 1770 5408 1776
rect 5368 1018 5396 1770
rect 5552 1018 5580 1906
rect 5736 1426 5764 3000
rect 5920 1970 5948 3000
rect 5908 1964 5960 1970
rect 5908 1906 5960 1912
rect 5724 1420 5776 1426
rect 5724 1362 5776 1368
rect 5356 1012 5408 1018
rect 5356 954 5408 960
rect 5540 1012 5592 1018
rect 5540 954 5592 960
rect 5736 950 5764 1362
rect 5920 1018 5948 1906
rect 6104 1902 6132 3000
rect 6092 1896 6144 1902
rect 6092 1838 6144 1844
rect 6104 1562 6132 1838
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 6288 1426 6316 3000
rect 6472 1970 6500 3000
rect 6460 1964 6512 1970
rect 6460 1906 6512 1912
rect 6276 1420 6328 1426
rect 6276 1362 6328 1368
rect 5908 1012 5960 1018
rect 5908 954 5960 960
rect 6288 950 6316 1362
rect 6472 1018 6500 1906
rect 6656 1902 6684 3000
rect 6644 1896 6696 1902
rect 6644 1838 6696 1844
rect 6656 1562 6684 1838
rect 6840 1562 6868 3000
rect 7024 1970 7052 3000
rect 7012 1964 7064 1970
rect 7012 1906 7064 1912
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 6828 1556 6880 1562
rect 6828 1498 6880 1504
rect 6840 1442 6868 1498
rect 6840 1414 6960 1442
rect 6460 1012 6512 1018
rect 6460 954 6512 960
rect 6932 950 6960 1414
rect 7024 1018 7052 1906
rect 7208 1902 7236 3000
rect 7196 1896 7248 1902
rect 7196 1838 7248 1844
rect 7208 1290 7236 1838
rect 7288 1828 7340 1834
rect 7288 1770 7340 1776
rect 7300 1562 7328 1770
rect 7392 1562 7420 3000
rect 7576 1970 7604 3000
rect 7564 1964 7616 1970
rect 7564 1906 7616 1912
rect 7288 1556 7340 1562
rect 7288 1498 7340 1504
rect 7380 1556 7432 1562
rect 7380 1498 7432 1504
rect 7196 1284 7248 1290
rect 7196 1226 7248 1232
rect 7012 1012 7064 1018
rect 7012 954 7064 960
rect 7392 950 7420 1498
rect 7576 1018 7604 1906
rect 7760 1562 7788 3000
rect 7944 1834 7972 3000
rect 7932 1828 7984 1834
rect 7932 1770 7984 1776
rect 8128 1562 8156 3000
rect 8312 1970 8340 3000
rect 8300 1964 8352 1970
rect 8300 1906 8352 1912
rect 8312 1850 8340 1906
rect 8220 1822 8340 1850
rect 7748 1556 7800 1562
rect 7748 1498 7800 1504
rect 8116 1556 8168 1562
rect 8116 1498 8168 1504
rect 7564 1012 7616 1018
rect 7564 954 7616 960
rect 5724 944 5776 950
rect 5724 886 5776 892
rect 6276 944 6328 950
rect 6276 886 6328 892
rect 6920 944 6972 950
rect 6920 886 6972 892
rect 7380 944 7432 950
rect 7380 886 7432 892
rect 5172 876 5224 882
rect 5172 818 5224 824
rect 7760 814 7788 1498
rect 8128 882 8156 1498
rect 8220 1018 8248 1822
rect 8496 1562 8524 3000
rect 8680 1970 8708 3000
rect 8864 1970 8892 3000
rect 9048 2530 9076 3000
rect 8956 2502 9076 2530
rect 8668 1964 8720 1970
rect 8668 1906 8720 1912
rect 8852 1964 8904 1970
rect 8852 1906 8904 1912
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8208 1012 8260 1018
rect 8208 954 8260 960
rect 8496 950 8524 1498
rect 8680 1018 8708 1906
rect 8956 1494 8984 2502
rect 9232 2394 9260 3000
rect 9048 2366 9260 2394
rect 9416 2394 9444 3000
rect 9416 2366 9536 2394
rect 9048 1970 9076 2366
rect 9116 2202 9436 2224
rect 9116 2150 9122 2202
rect 9174 2150 9186 2202
rect 9238 2150 9250 2202
rect 9302 2150 9314 2202
rect 9366 2150 9378 2202
rect 9430 2150 9436 2202
rect 9036 1964 9088 1970
rect 9036 1906 9088 1912
rect 9048 1562 9076 1906
rect 9036 1556 9088 1562
rect 9036 1498 9088 1504
rect 8944 1488 8996 1494
rect 8944 1430 8996 1436
rect 8956 1018 8984 1430
rect 9116 1188 9436 2150
rect 9508 1970 9536 2366
rect 9600 1970 9628 3000
rect 9784 2394 9812 3000
rect 9968 2530 9996 3000
rect 10152 2666 10180 3000
rect 10336 2802 10364 3000
rect 10336 2774 10456 2802
rect 10152 2638 10364 2666
rect 9968 2502 10272 2530
rect 9784 2366 10180 2394
rect 9496 1964 9548 1970
rect 9496 1906 9548 1912
rect 9588 1964 9640 1970
rect 9588 1906 9640 1912
rect 9508 1562 9536 1906
rect 9496 1556 9548 1562
rect 9496 1498 9548 1504
rect 9600 1222 9628 1906
rect 9756 1828 10076 2224
rect 10152 1970 10180 2366
rect 10140 1964 10192 1970
rect 10140 1906 10192 1912
rect 9756 1772 9768 1828
rect 9824 1772 9848 1828
rect 9904 1772 9928 1828
rect 9984 1772 10008 1828
rect 10064 1772 10076 1828
rect 9756 1748 10076 1772
rect 9756 1692 9768 1748
rect 9824 1692 9848 1748
rect 9904 1692 9928 1748
rect 9984 1692 10008 1748
rect 10064 1692 10076 1748
rect 9756 1668 10076 1692
rect 9756 1658 9768 1668
rect 9824 1658 9848 1668
rect 9904 1658 9928 1668
rect 9984 1658 10008 1668
rect 10064 1658 10076 1668
rect 9756 1606 9762 1658
rect 9824 1612 9826 1658
rect 10006 1612 10008 1658
rect 9814 1606 9826 1612
rect 9878 1606 9890 1612
rect 9942 1606 9954 1612
rect 10006 1606 10018 1612
rect 10070 1606 10076 1658
rect 9756 1588 10076 1606
rect 9756 1532 9768 1588
rect 9824 1532 9848 1588
rect 9904 1532 9928 1588
rect 9984 1532 10008 1588
rect 10064 1532 10076 1588
rect 10152 1562 10180 1906
rect 10244 1902 10272 2502
rect 10232 1896 10284 1902
rect 10232 1838 10284 1844
rect 10244 1562 10272 1838
rect 10336 1766 10364 2638
rect 10428 1970 10456 2774
rect 10416 1964 10468 1970
rect 10416 1906 10468 1912
rect 10324 1760 10376 1766
rect 10324 1702 10376 1708
rect 10336 1562 10364 1702
rect 9116 1132 9128 1188
rect 9184 1132 9208 1188
rect 9264 1132 9288 1188
rect 9344 1132 9368 1188
rect 9424 1132 9436 1188
rect 9588 1216 9640 1222
rect 9588 1158 9640 1164
rect 9116 1114 9436 1132
rect 9116 1062 9122 1114
rect 9174 1108 9186 1114
rect 9238 1108 9250 1114
rect 9302 1108 9314 1114
rect 9366 1108 9378 1114
rect 9184 1062 9186 1108
rect 9366 1062 9368 1108
rect 9430 1062 9436 1114
rect 9116 1052 9128 1062
rect 9184 1052 9208 1062
rect 9264 1052 9288 1062
rect 9344 1052 9368 1062
rect 9424 1052 9436 1062
rect 9116 1028 9436 1052
rect 8668 1012 8720 1018
rect 8668 954 8720 960
rect 8944 1012 8996 1018
rect 8944 954 8996 960
rect 9116 972 9128 1028
rect 9184 972 9208 1028
rect 9264 972 9288 1028
rect 9344 972 9368 1028
rect 9424 972 9436 1028
rect 8484 944 8536 950
rect 8484 886 8536 892
rect 9116 948 9436 972
rect 9116 892 9128 948
rect 9184 892 9208 948
rect 9264 892 9288 948
rect 9344 892 9368 948
rect 9424 892 9436 948
rect 8116 876 8168 882
rect 8116 818 8168 824
rect 7748 808 7800 814
rect 7748 750 7800 756
rect 1756 518 1762 570
rect 1814 518 1826 570
rect 1878 518 1890 570
rect 1942 518 1954 570
rect 2006 518 2018 570
rect 2070 518 2076 570
rect 1756 496 2076 518
rect 9116 496 9436 892
rect 9756 570 10076 1532
rect 10140 1556 10192 1562
rect 10140 1498 10192 1504
rect 10232 1556 10284 1562
rect 10232 1498 10284 1504
rect 10324 1556 10376 1562
rect 10324 1498 10376 1504
rect 10428 1494 10456 1906
rect 10520 1902 10548 3000
rect 10508 1896 10560 1902
rect 10508 1838 10560 1844
rect 10704 1834 10732 3000
rect 10888 1970 10916 3000
rect 10876 1964 10928 1970
rect 10876 1906 10928 1912
rect 10968 1896 11020 1902
rect 10968 1838 11020 1844
rect 10692 1828 10744 1834
rect 10692 1770 10744 1776
rect 10416 1488 10468 1494
rect 10416 1430 10468 1436
rect 10980 1358 11008 1838
rect 11072 1766 11100 3000
rect 11256 2038 11284 3000
rect 11244 2032 11296 2038
rect 11244 1974 11296 1980
rect 11440 1834 11468 3000
rect 11244 1828 11296 1834
rect 11244 1770 11296 1776
rect 11428 1828 11480 1834
rect 11428 1770 11480 1776
rect 11060 1760 11112 1766
rect 11060 1702 11112 1708
rect 11256 1562 11284 1770
rect 11624 1562 11652 3000
rect 11808 1902 11836 3000
rect 11992 2122 12020 3000
rect 11900 2094 12020 2122
rect 11796 1896 11848 1902
rect 11796 1838 11848 1844
rect 11900 1766 11928 2094
rect 11980 1964 12032 1970
rect 11980 1906 12032 1912
rect 12072 1964 12124 1970
rect 12072 1906 12124 1912
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11888 1760 11940 1766
rect 11888 1702 11940 1708
rect 11244 1556 11296 1562
rect 11244 1498 11296 1504
rect 11612 1556 11664 1562
rect 11612 1498 11664 1504
rect 10968 1352 11020 1358
rect 10968 1294 11020 1300
rect 11624 1018 11652 1498
rect 11808 1358 11836 1702
rect 11992 1562 12020 1906
rect 11980 1556 12032 1562
rect 11980 1498 12032 1504
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 11612 1012 11664 1018
rect 11612 954 11664 960
rect 12084 950 12112 1906
rect 12176 1562 12204 3000
rect 12360 1850 12388 3000
rect 12360 1834 12480 1850
rect 12256 1828 12308 1834
rect 12360 1828 12492 1834
rect 12360 1822 12440 1828
rect 12256 1770 12308 1776
rect 12440 1770 12492 1776
rect 12164 1556 12216 1562
rect 12164 1498 12216 1504
rect 12176 1018 12204 1498
rect 12268 1290 12296 1770
rect 12544 1562 12572 3000
rect 12728 2038 12756 3000
rect 12716 2032 12768 2038
rect 12716 1974 12768 1980
rect 12912 1986 12940 3000
rect 12912 1958 13032 1986
rect 13004 1902 13032 1958
rect 12900 1896 12952 1902
rect 12900 1838 12952 1844
rect 12992 1896 13044 1902
rect 12992 1838 13044 1844
rect 12532 1556 12584 1562
rect 12532 1498 12584 1504
rect 12256 1284 12308 1290
rect 12256 1226 12308 1232
rect 12164 1012 12216 1018
rect 12164 954 12216 960
rect 12072 944 12124 950
rect 12072 886 12124 892
rect 12544 882 12572 1498
rect 12912 1018 12940 1838
rect 13096 1562 13124 3000
rect 13280 1970 13308 3000
rect 13464 2106 13492 3000
rect 13452 2100 13504 2106
rect 13452 2042 13504 2048
rect 13544 2032 13596 2038
rect 13544 1974 13596 1980
rect 13268 1964 13320 1970
rect 13268 1906 13320 1912
rect 13556 1834 13584 1974
rect 13452 1828 13504 1834
rect 13452 1770 13504 1776
rect 13544 1828 13596 1834
rect 13544 1770 13596 1776
rect 13360 1760 13412 1766
rect 13360 1702 13412 1708
rect 13084 1556 13136 1562
rect 13084 1498 13136 1504
rect 13096 1018 13124 1498
rect 13372 1494 13400 1702
rect 13360 1488 13412 1494
rect 13360 1430 13412 1436
rect 12900 1012 12952 1018
rect 12900 954 12952 960
rect 13084 1012 13136 1018
rect 13084 954 13136 960
rect 13464 950 13492 1770
rect 13556 1358 13584 1770
rect 13648 1562 13676 3000
rect 13832 1902 13860 3000
rect 13820 1896 13872 1902
rect 13820 1838 13872 1844
rect 14016 1834 14044 3000
rect 14004 1828 14056 1834
rect 14004 1770 14056 1776
rect 14096 1760 14148 1766
rect 14096 1702 14148 1708
rect 13636 1556 13688 1562
rect 13636 1498 13688 1504
rect 13544 1352 13596 1358
rect 13544 1294 13596 1300
rect 13648 950 13676 1498
rect 14108 1018 14136 1702
rect 14200 1562 14228 3000
rect 14384 2122 14412 3000
rect 14280 2100 14332 2106
rect 14384 2094 14504 2122
rect 14568 2106 14596 3000
rect 14280 2042 14332 2048
rect 14292 1766 14320 2042
rect 14476 1970 14504 2094
rect 14556 2100 14608 2106
rect 14556 2042 14608 2048
rect 14372 1964 14424 1970
rect 14372 1906 14424 1912
rect 14464 1964 14516 1970
rect 14464 1906 14516 1912
rect 14280 1760 14332 1766
rect 14280 1702 14332 1708
rect 14188 1556 14240 1562
rect 14188 1498 14240 1504
rect 14200 1018 14228 1498
rect 14292 1426 14320 1702
rect 14280 1420 14332 1426
rect 14280 1362 14332 1368
rect 14096 1012 14148 1018
rect 14096 954 14148 960
rect 14188 1012 14240 1018
rect 14188 954 14240 960
rect 13452 944 13504 950
rect 13452 886 13504 892
rect 13636 944 13688 950
rect 13636 886 13688 892
rect 14384 882 14412 1906
rect 14752 1562 14780 3000
rect 14936 1986 14964 3000
rect 14936 1958 15056 1986
rect 14924 1896 14976 1902
rect 14924 1838 14976 1844
rect 14832 1828 14884 1834
rect 14832 1770 14884 1776
rect 14740 1556 14792 1562
rect 14740 1498 14792 1504
rect 14752 882 14780 1498
rect 14844 950 14872 1770
rect 14936 1018 14964 1838
rect 15028 1834 15056 1958
rect 15016 1828 15068 1834
rect 15016 1770 15068 1776
rect 15120 1562 15148 3000
rect 15200 2100 15252 2106
rect 15200 2042 15252 2048
rect 15212 1766 15240 2042
rect 15304 1850 15332 3000
rect 15488 1902 15516 3000
rect 15476 1896 15528 1902
rect 15304 1822 15424 1850
rect 15476 1838 15528 1844
rect 15200 1760 15252 1766
rect 15396 1714 15424 1822
rect 15568 1760 15620 1766
rect 15252 1708 15332 1714
rect 15200 1702 15332 1708
rect 15212 1686 15332 1702
rect 15396 1708 15568 1714
rect 15396 1702 15620 1708
rect 15396 1686 15608 1702
rect 15108 1556 15160 1562
rect 15160 1516 15240 1544
rect 15108 1498 15160 1504
rect 15212 1018 15240 1516
rect 15304 1290 15332 1686
rect 15672 1562 15700 3000
rect 15856 1970 15884 3000
rect 15752 1964 15804 1970
rect 15752 1906 15804 1912
rect 15844 1964 15896 1970
rect 15844 1906 15896 1912
rect 15660 1556 15712 1562
rect 15660 1498 15712 1504
rect 15292 1284 15344 1290
rect 15292 1226 15344 1232
rect 15672 1018 15700 1498
rect 15764 1494 15792 1906
rect 16040 1834 16068 3000
rect 15844 1828 15896 1834
rect 15844 1770 15896 1776
rect 16028 1828 16080 1834
rect 16028 1770 16080 1776
rect 15752 1488 15804 1494
rect 15752 1430 15804 1436
rect 14924 1012 14976 1018
rect 14924 954 14976 960
rect 15200 1012 15252 1018
rect 15200 954 15252 960
rect 15660 1012 15712 1018
rect 15660 954 15712 960
rect 15856 950 15884 1770
rect 16120 1760 16172 1766
rect 16120 1702 16172 1708
rect 16132 1358 16160 1702
rect 16224 1562 16252 3000
rect 16408 2038 16436 3000
rect 16396 2032 16448 2038
rect 16396 1974 16448 1980
rect 16396 1896 16448 1902
rect 16396 1838 16448 1844
rect 16212 1556 16264 1562
rect 16212 1498 16264 1504
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 16224 950 16252 1498
rect 16408 1018 16436 1838
rect 16592 1834 16620 3000
rect 16580 1828 16632 1834
rect 16580 1770 16632 1776
rect 16592 1494 16620 1770
rect 16776 1562 16804 3000
rect 16960 2106 16988 3000
rect 17144 2378 17172 3000
rect 17328 2394 17356 3000
rect 17512 2530 17540 3000
rect 17512 2502 17632 2530
rect 17132 2372 17184 2378
rect 17328 2366 17540 2394
rect 17132 2314 17184 2320
rect 17116 2202 17436 2224
rect 17116 2150 17122 2202
rect 17174 2150 17186 2202
rect 17238 2150 17250 2202
rect 17302 2150 17314 2202
rect 17366 2150 17378 2202
rect 17430 2150 17436 2202
rect 16948 2100 17000 2106
rect 16948 2042 17000 2048
rect 16948 1964 17000 1970
rect 16948 1906 17000 1912
rect 16856 1760 16908 1766
rect 16856 1702 16908 1708
rect 16764 1556 16816 1562
rect 16764 1498 16816 1504
rect 16580 1488 16632 1494
rect 16580 1430 16632 1436
rect 16776 1018 16804 1498
rect 16868 1290 16896 1702
rect 16856 1284 16908 1290
rect 16856 1226 16908 1232
rect 16396 1012 16448 1018
rect 16396 954 16448 960
rect 16764 1012 16816 1018
rect 16764 954 16816 960
rect 14832 944 14884 950
rect 14832 886 14884 892
rect 15844 944 15896 950
rect 15844 886 15896 892
rect 16212 944 16264 950
rect 16212 886 16264 892
rect 16960 882 16988 1906
rect 17116 1188 17436 2150
rect 17512 1562 17540 2366
rect 17604 1902 17632 2502
rect 17592 1896 17644 1902
rect 17592 1838 17644 1844
rect 17500 1556 17552 1562
rect 17500 1498 17552 1504
rect 17592 1556 17644 1562
rect 17696 1544 17724 3000
rect 17880 2394 17908 3000
rect 18064 2514 18092 3000
rect 18052 2508 18104 2514
rect 18052 2450 18104 2456
rect 17880 2366 18184 2394
rect 17644 1516 17724 1544
rect 17756 1828 18076 2224
rect 18156 1970 18184 2366
rect 18144 1964 18196 1970
rect 18144 1906 18196 1912
rect 17756 1772 17768 1828
rect 17824 1772 17848 1828
rect 17904 1772 17928 1828
rect 17984 1772 18008 1828
rect 18064 1772 18076 1828
rect 17756 1748 18076 1772
rect 17756 1692 17768 1748
rect 17824 1692 17848 1748
rect 17904 1692 17928 1748
rect 17984 1692 18008 1748
rect 18064 1692 18076 1748
rect 17756 1668 18076 1692
rect 17756 1658 17768 1668
rect 17824 1658 17848 1668
rect 17904 1658 17928 1668
rect 17984 1658 18008 1668
rect 18064 1658 18076 1668
rect 17756 1606 17762 1658
rect 17824 1612 17826 1658
rect 18006 1612 18008 1658
rect 17814 1606 17826 1612
rect 17878 1606 17890 1612
rect 17942 1606 17954 1612
rect 18006 1606 18018 1612
rect 18070 1606 18076 1658
rect 17756 1588 18076 1606
rect 17756 1532 17768 1588
rect 17824 1532 17848 1588
rect 17904 1532 17928 1588
rect 17984 1532 18008 1588
rect 18064 1532 18076 1588
rect 18248 1562 18276 3000
rect 18972 2508 19024 2514
rect 18972 2450 19024 2456
rect 18328 2372 18380 2378
rect 18328 2314 18380 2320
rect 18340 1834 18368 2314
rect 18788 2032 18840 2038
rect 18788 1974 18840 1980
rect 18420 1896 18472 1902
rect 18420 1838 18472 1844
rect 18328 1828 18380 1834
rect 18328 1770 18380 1776
rect 17592 1498 17644 1504
rect 17116 1132 17128 1188
rect 17184 1132 17208 1188
rect 17264 1132 17288 1188
rect 17344 1132 17368 1188
rect 17424 1132 17436 1188
rect 17116 1114 17436 1132
rect 17116 1062 17122 1114
rect 17174 1108 17186 1114
rect 17238 1108 17250 1114
rect 17302 1108 17314 1114
rect 17366 1108 17378 1114
rect 17184 1062 17186 1108
rect 17366 1062 17368 1108
rect 17430 1062 17436 1114
rect 17116 1052 17128 1062
rect 17184 1052 17208 1062
rect 17264 1052 17288 1062
rect 17344 1052 17368 1062
rect 17424 1052 17436 1062
rect 17116 1028 17436 1052
rect 17116 972 17128 1028
rect 17184 972 17208 1028
rect 17264 972 17288 1028
rect 17344 972 17368 1028
rect 17424 972 17436 1028
rect 17512 1018 17540 1498
rect 17116 948 17436 972
rect 17500 1012 17552 1018
rect 17500 954 17552 960
rect 17116 892 17128 948
rect 17184 892 17208 948
rect 17264 892 17288 948
rect 17344 892 17368 948
rect 17424 892 17436 948
rect 12532 876 12584 882
rect 12532 818 12584 824
rect 14372 876 14424 882
rect 14372 818 14424 824
rect 14740 876 14792 882
rect 14740 818 14792 824
rect 16948 876 17000 882
rect 16948 818 17000 824
rect 9756 518 9762 570
rect 9814 518 9826 570
rect 9878 518 9890 570
rect 9942 518 9954 570
rect 10006 518 10018 570
rect 10070 518 10076 570
rect 9756 496 10076 518
rect 17116 496 17436 892
rect 17756 570 18076 1532
rect 18144 1556 18196 1562
rect 18144 1498 18196 1504
rect 18236 1556 18288 1562
rect 18236 1498 18288 1504
rect 18156 1018 18184 1498
rect 18248 1018 18276 1498
rect 18340 1426 18368 1770
rect 18432 1562 18460 1838
rect 18420 1556 18472 1562
rect 18420 1498 18472 1504
rect 18328 1420 18380 1426
rect 18328 1362 18380 1368
rect 18800 1358 18828 1974
rect 18984 1902 19012 2450
rect 19340 1964 19392 1970
rect 19340 1906 19392 1912
rect 18972 1896 19024 1902
rect 18972 1838 19024 1844
rect 18788 1352 18840 1358
rect 18788 1294 18840 1300
rect 18984 1018 19012 1838
rect 19352 1562 19380 1906
rect 19340 1556 19392 1562
rect 19340 1498 19392 1504
rect 18144 1012 18196 1018
rect 18144 954 18196 960
rect 18236 1012 18288 1018
rect 18236 954 18288 960
rect 18972 1012 19024 1018
rect 18972 954 19024 960
rect 17756 518 17762 570
rect 17814 518 17826 570
rect 17878 518 17890 570
rect 17942 518 17954 570
rect 18006 518 18018 570
rect 18070 518 18076 570
rect 17756 496 18076 518
<< via2 >>
rect 1768 1772 1824 1828
rect 1848 1772 1904 1828
rect 1928 1772 1984 1828
rect 2008 1772 2064 1828
rect 1768 1692 1824 1748
rect 1848 1692 1904 1748
rect 1928 1692 1984 1748
rect 2008 1692 2064 1748
rect 1768 1658 1824 1668
rect 1848 1658 1904 1668
rect 1928 1658 1984 1668
rect 2008 1658 2064 1668
rect 1768 1612 1814 1658
rect 1814 1612 1824 1658
rect 1848 1612 1878 1658
rect 1878 1612 1890 1658
rect 1890 1612 1904 1658
rect 1928 1612 1942 1658
rect 1942 1612 1954 1658
rect 1954 1612 1984 1658
rect 2008 1612 2018 1658
rect 2018 1612 2064 1658
rect 1768 1532 1824 1588
rect 1848 1532 1904 1588
rect 1928 1532 1984 1588
rect 2008 1532 2064 1588
rect 1128 1132 1184 1188
rect 1208 1132 1264 1188
rect 1288 1132 1344 1188
rect 1368 1132 1424 1188
rect 1128 1062 1174 1108
rect 1174 1062 1184 1108
rect 1208 1062 1238 1108
rect 1238 1062 1250 1108
rect 1250 1062 1264 1108
rect 1288 1062 1302 1108
rect 1302 1062 1314 1108
rect 1314 1062 1344 1108
rect 1368 1062 1378 1108
rect 1378 1062 1424 1108
rect 1128 1052 1184 1062
rect 1208 1052 1264 1062
rect 1288 1052 1344 1062
rect 1368 1052 1424 1062
rect 1128 972 1184 1028
rect 1208 972 1264 1028
rect 1288 972 1344 1028
rect 1368 972 1424 1028
rect 1128 892 1184 948
rect 1208 892 1264 948
rect 1288 892 1344 948
rect 1368 892 1424 948
rect 9768 1772 9824 1828
rect 9848 1772 9904 1828
rect 9928 1772 9984 1828
rect 10008 1772 10064 1828
rect 9768 1692 9824 1748
rect 9848 1692 9904 1748
rect 9928 1692 9984 1748
rect 10008 1692 10064 1748
rect 9768 1658 9824 1668
rect 9848 1658 9904 1668
rect 9928 1658 9984 1668
rect 10008 1658 10064 1668
rect 9768 1612 9814 1658
rect 9814 1612 9824 1658
rect 9848 1612 9878 1658
rect 9878 1612 9890 1658
rect 9890 1612 9904 1658
rect 9928 1612 9942 1658
rect 9942 1612 9954 1658
rect 9954 1612 9984 1658
rect 10008 1612 10018 1658
rect 10018 1612 10064 1658
rect 9768 1532 9824 1588
rect 9848 1532 9904 1588
rect 9928 1532 9984 1588
rect 10008 1532 10064 1588
rect 9128 1132 9184 1188
rect 9208 1132 9264 1188
rect 9288 1132 9344 1188
rect 9368 1132 9424 1188
rect 9128 1062 9174 1108
rect 9174 1062 9184 1108
rect 9208 1062 9238 1108
rect 9238 1062 9250 1108
rect 9250 1062 9264 1108
rect 9288 1062 9302 1108
rect 9302 1062 9314 1108
rect 9314 1062 9344 1108
rect 9368 1062 9378 1108
rect 9378 1062 9424 1108
rect 9128 1052 9184 1062
rect 9208 1052 9264 1062
rect 9288 1052 9344 1062
rect 9368 1052 9424 1062
rect 9128 972 9184 1028
rect 9208 972 9264 1028
rect 9288 972 9344 1028
rect 9368 972 9424 1028
rect 9128 892 9184 948
rect 9208 892 9264 948
rect 9288 892 9344 948
rect 9368 892 9424 948
rect 17768 1772 17824 1828
rect 17848 1772 17904 1828
rect 17928 1772 17984 1828
rect 18008 1772 18064 1828
rect 17768 1692 17824 1748
rect 17848 1692 17904 1748
rect 17928 1692 17984 1748
rect 18008 1692 18064 1748
rect 17768 1658 17824 1668
rect 17848 1658 17904 1668
rect 17928 1658 17984 1668
rect 18008 1658 18064 1668
rect 17768 1612 17814 1658
rect 17814 1612 17824 1658
rect 17848 1612 17878 1658
rect 17878 1612 17890 1658
rect 17890 1612 17904 1658
rect 17928 1612 17942 1658
rect 17942 1612 17954 1658
rect 17954 1612 17984 1658
rect 18008 1612 18018 1658
rect 18018 1612 18064 1658
rect 17768 1532 17824 1588
rect 17848 1532 17904 1588
rect 17928 1532 17984 1588
rect 18008 1532 18064 1588
rect 17128 1132 17184 1188
rect 17208 1132 17264 1188
rect 17288 1132 17344 1188
rect 17368 1132 17424 1188
rect 17128 1062 17174 1108
rect 17174 1062 17184 1108
rect 17208 1062 17238 1108
rect 17238 1062 17250 1108
rect 17250 1062 17264 1108
rect 17288 1062 17302 1108
rect 17302 1062 17314 1108
rect 17314 1062 17344 1108
rect 17368 1062 17378 1108
rect 17378 1062 17424 1108
rect 17128 1052 17184 1062
rect 17208 1052 17264 1062
rect 17288 1052 17344 1062
rect 17368 1052 17424 1062
rect 17128 972 17184 1028
rect 17208 972 17264 1028
rect 17288 972 17344 1028
rect 17368 972 17424 1028
rect 17128 892 17184 948
rect 17208 892 17264 948
rect 17288 892 17344 948
rect 17368 892 17424 948
<< metal3 >>
rect 228 1828 19828 1840
rect 228 1772 1768 1828
rect 1824 1772 1848 1828
rect 1904 1772 1928 1828
rect 1984 1772 2008 1828
rect 2064 1772 9768 1828
rect 9824 1772 9848 1828
rect 9904 1772 9928 1828
rect 9984 1772 10008 1828
rect 10064 1772 17768 1828
rect 17824 1772 17848 1828
rect 17904 1772 17928 1828
rect 17984 1772 18008 1828
rect 18064 1772 19828 1828
rect 228 1748 19828 1772
rect 228 1692 1768 1748
rect 1824 1692 1848 1748
rect 1904 1692 1928 1748
rect 1984 1692 2008 1748
rect 2064 1692 9768 1748
rect 9824 1692 9848 1748
rect 9904 1692 9928 1748
rect 9984 1692 10008 1748
rect 10064 1692 17768 1748
rect 17824 1692 17848 1748
rect 17904 1692 17928 1748
rect 17984 1692 18008 1748
rect 18064 1692 19828 1748
rect 228 1668 19828 1692
rect 228 1612 1768 1668
rect 1824 1612 1848 1668
rect 1904 1612 1928 1668
rect 1984 1612 2008 1668
rect 2064 1612 9768 1668
rect 9824 1612 9848 1668
rect 9904 1612 9928 1668
rect 9984 1612 10008 1668
rect 10064 1612 17768 1668
rect 17824 1612 17848 1668
rect 17904 1612 17928 1668
rect 17984 1612 18008 1668
rect 18064 1612 19828 1668
rect 228 1588 19828 1612
rect 228 1532 1768 1588
rect 1824 1532 1848 1588
rect 1904 1532 1928 1588
rect 1984 1532 2008 1588
rect 2064 1532 9768 1588
rect 9824 1532 9848 1588
rect 9904 1532 9928 1588
rect 9984 1532 10008 1588
rect 10064 1532 17768 1588
rect 17824 1532 17848 1588
rect 17904 1532 17928 1588
rect 17984 1532 18008 1588
rect 18064 1532 19828 1588
rect 228 1520 19828 1532
rect 228 1188 19828 1200
rect 228 1132 1128 1188
rect 1184 1132 1208 1188
rect 1264 1132 1288 1188
rect 1344 1132 1368 1188
rect 1424 1132 9128 1188
rect 9184 1132 9208 1188
rect 9264 1132 9288 1188
rect 9344 1132 9368 1188
rect 9424 1132 17128 1188
rect 17184 1132 17208 1188
rect 17264 1132 17288 1188
rect 17344 1132 17368 1188
rect 17424 1132 19828 1188
rect 228 1108 19828 1132
rect 228 1052 1128 1108
rect 1184 1052 1208 1108
rect 1264 1052 1288 1108
rect 1344 1052 1368 1108
rect 1424 1052 9128 1108
rect 9184 1052 9208 1108
rect 9264 1052 9288 1108
rect 9344 1052 9368 1108
rect 9424 1052 17128 1108
rect 17184 1052 17208 1108
rect 17264 1052 17288 1108
rect 17344 1052 17368 1108
rect 17424 1052 19828 1108
rect 228 1028 19828 1052
rect 228 972 1128 1028
rect 1184 972 1208 1028
rect 1264 972 1288 1028
rect 1344 972 1368 1028
rect 1424 972 9128 1028
rect 9184 972 9208 1028
rect 9264 972 9288 1028
rect 9344 972 9368 1028
rect 9424 972 17128 1028
rect 17184 972 17208 1028
rect 17264 972 17288 1028
rect 17344 972 17368 1028
rect 17424 972 19828 1028
rect 228 948 19828 972
rect 228 892 1128 948
rect 1184 892 1208 948
rect 1264 892 1288 948
rect 1344 892 1368 948
rect 1424 892 9128 948
rect 9184 892 9208 948
rect 9264 892 9288 948
rect 9344 892 9368 948
rect 9424 892 17128 948
rect 17184 892 17208 948
rect 17264 892 17288 948
rect 17344 892 17368 948
rect 17424 892 19828 948
rect 228 880 19828 892
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_1_HI
timestamp 21601
transform -1 0 1748 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_2_HI
timestamp 21601
transform -1 0 3680 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_3_HI
timestamp 21601
transform -1 0 4140 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_4_HI
timestamp 21601
transform -1 0 3956 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_5_HI
timestamp 21601
transform -1 0 3772 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_6_HI
timestamp 21601
transform -1 0 4324 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_7_HI
timestamp 21601
transform -1 0 4508 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_8_HI
timestamp 21601
transform -1 0 4692 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_9_HI
timestamp 21601
transform -1 0 4324 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_10_HI
timestamp 21601
transform -1 0 4876 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_11_HI
timestamp 21601
transform -1 0 5060 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_12_HI
timestamp 21601
transform -1 0 1104 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_13_HI
timestamp 21601
transform -1 0 5336 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_14_HI
timestamp 21601
transform -1 0 5704 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_15_HI
timestamp 21601
transform -1 0 6256 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_16_HI
timestamp 21601
transform -1 0 5980 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_17_HI
timestamp 21601
transform -1 0 5796 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_18_HI
timestamp 21601
transform -1 0 6808 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_19_HI
timestamp 21601
transform -1 0 6532 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_20_HI
timestamp 21601
transform -1 0 6348 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_21_HI
timestamp 21601
transform -1 0 7360 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_22_HI
timestamp 21601
transform -1 0 7084 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_23_HI
timestamp 21601
transform -1 0 1288 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_24_HI
timestamp 21601
transform -1 0 6900 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_25_HI
timestamp 21601
transform -1 0 7912 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_26_HI
timestamp 21601
transform -1 0 7636 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_27_HI
timestamp 21601
transform -1 0 8464 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_28_HI
timestamp 21601
transform -1 0 7452 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_29_HI
timestamp 21601
transform -1 0 9200 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_30_HI
timestamp 21601
transform -1 0 8280 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_31_HI
timestamp 21601
transform -1 0 9016 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_32_HI
timestamp 21601
transform -1 0 8740 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_33_HI
timestamp 21601
transform -1 0 8280 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_34_HI
timestamp 21601
transform -1 0 2668 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_35_HI
timestamp 21601
transform -1 0 9568 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_36_HI
timestamp 21601
transform -1 0 9108 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_37_HI
timestamp 21601
transform -1 0 9568 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_38_HI
timestamp 21601
transform -1 0 9844 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_39_HI
timestamp 21601
transform -1 0 10120 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_40_HI
timestamp 21601
transform -1 0 10396 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_41_HI
timestamp 21601
transform -1 0 10856 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_42_HI
timestamp 21601
transform -1 0 11132 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_43_HI
timestamp 21601
transform -1 0 11408 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_44_HI
timestamp 21601
transform -1 0 11684 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_45_HI
timestamp 21601
transform -1 0 1472 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_46_HI
timestamp 21601
transform -1 0 12144 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_47_HI
timestamp 21601
transform -1 0 13064 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_48_HI
timestamp 21601
transform -1 0 12512 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_49_HI
timestamp 21601
transform -1 0 13616 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_50_HI
timestamp 21601
transform -1 0 12144 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_51_HI
timestamp 21601
transform -1 0 13064 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_52_HI
timestamp 21601
transform -1 0 14168 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_53_HI
timestamp 21601
transform -1 0 12696 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_54_HI
timestamp 21601
transform -1 0 13708 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_55_HI
timestamp 21601
transform -1 0 13432 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_56_HI
timestamp 21601
transform -1 0 2300 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_57_HI
timestamp 21601
transform -1 0 14720 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_58_HI
timestamp 21601
transform -1 0 14260 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_59_HI
timestamp 21601
transform -1 0 13892 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_60_HI
timestamp 21601
transform -1 0 14536 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_61_HI
timestamp 21601
transform -1 0 15640 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_62_HI
timestamp 21601
transform -1 0 14720 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_63_HI
timestamp 21601
transform -1 0 15088 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_64_HI
timestamp 21601
transform -1 0 15364 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_65_HI
timestamp 21601
transform -1 0 14904 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_66_HI
timestamp 21601
transform -1 0 16284 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_67_HI
timestamp 21601
transform -1 0 2852 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_68_HI
timestamp 21601
transform -1 0 16744 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_69_HI
timestamp 21601
transform -1 0 15548 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_70_HI
timestamp 21601
transform -1 0 16284 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_71_HI
timestamp 21601
transform -1 0 15732 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_72_HI
timestamp 21601
transform -1 0 17296 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_73_HI
timestamp 21601
transform -1 0 16836 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_74_HI
timestamp 21601
transform -1 0 16468 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_75_HI
timestamp 21601
transform -1 0 17112 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_76_HI
timestamp 21601
transform -1 0 18216 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_77_HI
timestamp 21601
transform -1 0 17296 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_78_HI
timestamp 21601
transform -1 0 3128 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_79_HI
timestamp 21601
transform -1 0 19412 0 1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_80_HI
timestamp 21601
transform -1 0 18768 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_81_HI
timestamp 21601
transform -1 0 17480 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_82_HI
timestamp 21601
transform -1 0 18952 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_83_HI
timestamp 21601
transform -1 0 19136 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_84_HI
timestamp 21601
transform -1 0 17848 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_85_HI
timestamp 21601
transform -1 0 19320 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_86_HI
timestamp 21601
transform -1 0 18216 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_87_HI
timestamp 21601
transform -1 0 19504 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_88_HI
timestamp 21601
transform -1 0 19412 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_89_HI
timestamp 21601
transform -1 0 2852 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_90_HI
timestamp 21601
transform -1 0 18768 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_vccd1_tie_high_91_HI
timestamp 21601
transform -1 0 3404 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3
timestamp 21601
transform 1 0 552 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6
timestamp 21601
transform 1 0 828 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9
timestamp 21601
transform 1 0 1104 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12
timestamp 21601
transform 1 0 1380 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15
timestamp 21601
transform 1 0 1656 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18
timestamp 21601
transform 1 0 1932 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21
timestamp 21601
transform 1 0 2208 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31
timestamp 21601
transform 1 0 3128 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34
timestamp 21601
transform 1 0 3404 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37
timestamp 21601
transform 1 0 3680 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52
timestamp 21601
transform 1 0 5060 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55
timestamp 21601
transform 1 0 5336 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59
timestamp 21601
transform 1 0 5704 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62
timestamp 21601
transform 1 0 5980 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65
timestamp 21601
transform 1 0 6256 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68
timestamp 21601
transform 1 0 6532 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71
timestamp 21601
transform 1 0 6808 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74
timestamp 21601
transform 1 0 7084 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77
timestamp 21601
transform 1 0 7360 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_80
timestamp 21601
transform 1 0 7636 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 21601
transform 1 0 7912 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_89
timestamp 21601
transform 1 0 8464 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 21601
transform 1 0 8740 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_97
timestamp 21601
transform 1 0 9200 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_101
timestamp 21601
transform 1 0 9568 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_104
timestamp 21601
transform 1 0 9844 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_107
timestamp 21601
transform 1 0 10120 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_110
timestamp 21601
transform 1 0 10396 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_113
timestamp 21601
transform 1 0 10672 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_116
timestamp 21601
transform 1 0 10948 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_119
timestamp 21601
transform 1 0 11224 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_122
timestamp 21601
transform 1 0 11500 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_125
timestamp 21601
transform 1 0 11776 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_129
timestamp 21601
transform 1 0 12144 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_135
timestamp 21601
transform 1 0 12696 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 21601
transform 1 0 13064 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_143
timestamp 21601
transform 1 0 13432 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_148
timestamp 21601
transform 1 0 13892 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_152
timestamp 21601
transform 1 0 14260 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_161
timestamp 21601
transform 1 0 15088 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_169
timestamp 21601
transform 1 0 15824 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_176
timestamp 21601
transform 1 0 16468 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_180
timestamp 21601
transform 1 0 16836 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_187
timestamp 21601
transform 1 0 17480 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_191
timestamp 21601
transform 1 0 17848 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 21601
transform 1 0 18216 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 21601
transform 1 0 18400 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_201
timestamp 21601
transform 1 0 18768 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_204
timestamp 21601
transform 1 0 19044 0 1 544
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_208
timestamp 21601
transform 1 0 19412 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_3
timestamp 21601
transform 1 0 552 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_6
timestamp 21601
transform 1 0 828 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_9
timestamp 21601
transform 1 0 1104 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_12
timestamp 21601
transform 1 0 1380 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_19
timestamp 21601
transform 1 0 2024 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 21601
transform 1 0 2576 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_31
timestamp 21601
transform 1 0 3128 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp 21601
transform 1 0 3496 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_41
timestamp 21601
transform 1 0 4048 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_47
timestamp 21601
transform 1 0 4600 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_51
timestamp 21601
transform 1 0 4968 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 21601
transform 1 0 5336 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_57
timestamp 21601
transform 1 0 5520 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_63
timestamp 21601
transform 1 0 6072 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_69
timestamp 21601
transform 1 0 6624 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 21601
transform 1 0 7176 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_81
timestamp 21601
transform 1 0 7728 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_85
timestamp 21601
transform 1 0 8096 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_89
timestamp 21601
transform 1 0 8464 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 21601
transform 1 0 8832 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_101
timestamp 21601
transform 1 0 9568 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_104
timestamp 21601
transform 1 0 9844 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_107
timestamp 21601
transform 1 0 10120 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_110
timestamp 21601
transform 1 0 10396 0 -1 1632
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_1_115
timestamp 21601
transform 1 0 10856 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_118
timestamp 21601
transform 1 0 11132 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_121
timestamp 21601
transform 1 0 11408 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_129
timestamp 21601
transform 1 0 12144 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_133
timestamp 21601
transform 1 0 12512 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_139
timestamp 21601
transform 1 0 13064 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_145
timestamp 21601
transform 1 0 13616 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_151
timestamp 21601
transform 1 0 14168 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_157
timestamp 21601
transform 1 0 14720 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_161
timestamp 21601
transform 1 0 15088 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 21601
transform 1 0 15640 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_179
timestamp 21601
transform 1 0 16744 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_185
timestamp 21601
transform 1 0 17296 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_189
timestamp 21601
transform 1 0 17664 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_195
timestamp 21601
transform 1 0 18216 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_3
timestamp 21601
transform 1 0 552 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_2_6
timestamp 21601
transform 1 0 828 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_111
timestamp 21601
transform 1 0 10488 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_208
timestamp 21601
transform 1 0 19412 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_3
timestamp 21601
transform 1 0 276 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 21601
transform -1 0 19780 0 1 544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_4
timestamp 21601
transform 1 0 276 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 21601
transform -1 0 19780 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_5
timestamp 21601
transform 1 0 276 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 21601
transform -1 0 19780 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_6
timestamp 21601
transform 1 0 2852 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_7
timestamp 21601
transform 1 0 5428 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_8
timestamp 21601
transform 1 0 8004 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_9
timestamp 21601
transform 1 0 10580 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_10
timestamp 21601
transform 1 0 13156 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_11
timestamp 21601
transform 1 0 15732 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_12
timestamp 21601
transform 1 0 18308 0 1 544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_13
timestamp 21601
transform 1 0 5428 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_14
timestamp 21601
transform 1 0 10580 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_15
timestamp 21601
transform 1 0 15732 0 -1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_16
timestamp 21601
transform 1 0 2852 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_17
timestamp 21601
transform 1 0 5428 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_18
timestamp 21601
transform 1 0 8004 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_19
timestamp 21601
transform 1 0 10580 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_20
timestamp 21601
transform 1 0 13156 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_21
timestamp 21601
transform 1 0 15732 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_22
timestamp 21601
transform 1 0 18308 0 1 1632
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_1
timestamp 1562557784
transform 1 0 1748 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_2
timestamp 1562557784
transform -1 0 3496 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_3
timestamp 1562557784
transform 1 0 3772 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_4
timestamp 1562557784
transform -1 0 3772 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_5
timestamp 1562557784
transform 1 0 3772 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_6
timestamp 1562557784
transform 1 0 4324 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_7
timestamp 1562557784
transform -1 0 4324 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_8
timestamp 1562557784
transform 1 0 4692 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_9
timestamp 1562557784
transform 1 0 4324 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_10
timestamp 1562557784
transform 1 0 5060 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_11
timestamp 1562557784
transform -1 0 4876 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_12
timestamp 1562557784
transform -1 0 1748 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_13
timestamp 1562557784
transform -1 0 5152 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_14
timestamp 1562557784
transform -1 0 5428 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_15
timestamp 1562557784
transform 1 0 5796 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_16
timestamp 1562557784
transform -1 0 5796 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_17
timestamp 1562557784
transform 1 0 5796 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_18
timestamp 1562557784
transform 1 0 6348 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_19
timestamp 1562557784
transform -1 0 6348 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_20
timestamp 1562557784
transform 1 0 6348 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_21
timestamp 1562557784
transform 1 0 6900 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_22
timestamp 1562557784
transform -1 0 6900 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_23
timestamp 1562557784
transform -1 0 2024 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_24
timestamp 1562557784
transform 1 0 6900 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_25
timestamp 1562557784
transform 1 0 7452 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_26
timestamp 1562557784
transform -1 0 7452 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_27
timestamp 1562557784
transform 1 0 7820 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_28
timestamp 1562557784
transform 1 0 7452 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_29
timestamp 1562557784
transform 1 0 8188 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_30
timestamp 1562557784
transform -1 0 8004 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_31
timestamp 1562557784
transform 1 0 8556 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_32
timestamp 1562557784
transform -1 0 8556 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_33
timestamp 1562557784
transform -1 0 8832 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_34
timestamp 1562557784
transform 1 0 2300 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_35
timestamp 1562557784
transform 1 0 9108 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_36
timestamp 1562557784
transform -1 0 9108 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_37
timestamp 1562557784
transform -1 0 9384 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_38
timestamp 1562557784
transform -1 0 9660 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_39
timestamp 1562557784
transform -1 0 9936 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_40
timestamp 1562557784
transform 1 0 9936 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_41
timestamp 1562557784
transform 1 0 10212 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_42
timestamp 1562557784
transform 1 0 10672 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_43
timestamp 1562557784
transform 1 0 10948 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_44
timestamp 1562557784
transform 1 0 11224 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_45
timestamp 1562557784
transform -1 0 2300 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_46
timestamp 1562557784
transform 1 0 11500 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_47
timestamp 1562557784
transform 1 0 11776 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_48
timestamp 1562557784
transform 1 0 12052 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_49
timestamp 1562557784
transform 1 0 12328 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_50
timestamp 1562557784
transform 1 0 11684 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_51
timestamp 1562557784
transform 1 0 12604 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_52
timestamp 1562557784
transform 1 0 12880 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_53
timestamp 1562557784
transform 1 0 12236 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_54
timestamp 1562557784
transform 1 0 13248 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_55
timestamp 1562557784
transform 1 0 12604 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_56
timestamp 1562557784
transform 1 0 2300 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_57
timestamp 1562557784
transform 1 0 13524 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_58
timestamp 1562557784
transform 1 0 13800 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_59
timestamp 1562557784
transform 1 0 13156 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_60
timestamp 1562557784
transform 1 0 14076 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_61
timestamp 1562557784
transform 1 0 14352 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_62
timestamp 1562557784
transform 1 0 13708 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_63
timestamp 1562557784
transform 1 0 14628 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_64
timestamp 1562557784
transform 1 0 14904 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_65
timestamp 1562557784
transform 1 0 14260 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_66
timestamp 1562557784
transform 1 0 15180 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_67
timestamp 1562557784
transform 1 0 2852 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_68
timestamp 1562557784
transform 1 0 15456 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_69
timestamp 1562557784
transform 1 0 14812 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_70
timestamp 1562557784
transform 1 0 15824 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_71
timestamp 1562557784
transform 1 0 15180 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_72
timestamp 1562557784
transform 1 0 16100 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_73
timestamp 1562557784
transform 1 0 16376 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_74
timestamp 1562557784
transform 1 0 15824 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_75
timestamp 1562557784
transform 1 0 16652 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_76
timestamp 1562557784
transform 1 0 16928 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_77
timestamp 1562557784
transform 1 0 16284 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_78
timestamp 1562557784
transform -1 0 2852 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_79
timestamp 1562557784
transform -1 0 17480 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_80
timestamp 1562557784
transform 1 0 17480 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_81
timestamp 1562557784
transform 1 0 16836 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_82
timestamp 1562557784
transform 1 0 17756 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_83
timestamp 1562557784
transform 1 0 18032 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_84
timestamp 1562557784
transform 1 0 17388 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_85
timestamp 1562557784
transform 1 0 18400 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_86
timestamp 1562557784
transform 1 0 17756 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_87
timestamp 1562557784
transform 1 0 18676 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_88
timestamp 1562557784
transform 1 0 18952 0 1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_89
timestamp 1562557784
transform 1 0 3220 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_90
timestamp 1562557784
transform 1 0 18308 0 -1 1632
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  vccd1_tie_high_91
timestamp 1562557784
transform -1 0 3220 0 1 1632
box -38 -48 314 592
<< labels >>
flabel metal2 s 1674 3000 1730 3400 0 FreeSans 224 90 0 0 HI[0]
port 0 nsew signal output
flabel metal2 s 3514 3000 3570 3400 0 FreeSans 224 90 0 0 HI[10]
port 1 nsew signal output
flabel metal2 s 3698 3000 3754 3400 0 FreeSans 224 90 0 0 HI[11]
port 2 nsew signal output
flabel metal2 s 3882 3000 3938 3400 0 FreeSans 224 90 0 0 HI[12]
port 3 nsew signal output
flabel metal2 s 4066 3000 4122 3400 0 FreeSans 224 90 0 0 HI[13]
port 4 nsew signal output
flabel metal2 s 4250 3000 4306 3400 0 FreeSans 224 90 0 0 HI[14]
port 5 nsew signal output
flabel metal2 s 4434 3000 4490 3400 0 FreeSans 224 90 0 0 HI[15]
port 6 nsew signal output
flabel metal2 s 4618 3000 4674 3400 0 FreeSans 224 90 0 0 HI[16]
port 7 nsew signal output
flabel metal2 s 4802 3000 4858 3400 0 FreeSans 224 90 0 0 HI[17]
port 8 nsew signal output
flabel metal2 s 4986 3000 5042 3400 0 FreeSans 224 90 0 0 HI[18]
port 9 nsew signal output
flabel metal2 s 5170 3000 5226 3400 0 FreeSans 224 90 0 0 HI[19]
port 10 nsew signal output
flabel metal2 s 1858 3000 1914 3400 0 FreeSans 224 90 0 0 HI[1]
port 11 nsew signal output
flabel metal2 s 5354 3000 5410 3400 0 FreeSans 224 90 0 0 HI[20]
port 12 nsew signal output
flabel metal2 s 5538 3000 5594 3400 0 FreeSans 224 90 0 0 HI[21]
port 13 nsew signal output
flabel metal2 s 5722 3000 5778 3400 0 FreeSans 224 90 0 0 HI[22]
port 14 nsew signal output
flabel metal2 s 5906 3000 5962 3400 0 FreeSans 224 90 0 0 HI[23]
port 15 nsew signal output
flabel metal2 s 6090 3000 6146 3400 0 FreeSans 224 90 0 0 HI[24]
port 16 nsew signal output
flabel metal2 s 6274 3000 6330 3400 0 FreeSans 224 90 0 0 HI[25]
port 17 nsew signal output
flabel metal2 s 6458 3000 6514 3400 0 FreeSans 224 90 0 0 HI[26]
port 18 nsew signal output
flabel metal2 s 6642 3000 6698 3400 0 FreeSans 224 90 0 0 HI[27]
port 19 nsew signal output
flabel metal2 s 6826 3000 6882 3400 0 FreeSans 224 90 0 0 HI[28]
port 20 nsew signal output
flabel metal2 s 7010 3000 7066 3400 0 FreeSans 224 90 0 0 HI[29]
port 21 nsew signal output
flabel metal2 s 2042 3000 2098 3400 0 FreeSans 224 90 0 0 HI[2]
port 22 nsew signal output
flabel metal2 s 7194 3000 7250 3400 0 FreeSans 224 90 0 0 HI[30]
port 23 nsew signal output
flabel metal2 s 7378 3000 7434 3400 0 FreeSans 224 90 0 0 HI[31]
port 24 nsew signal output
flabel metal2 s 7562 3000 7618 3400 0 FreeSans 224 90 0 0 HI[32]
port 25 nsew signal output
flabel metal2 s 7746 3000 7802 3400 0 FreeSans 224 90 0 0 HI[33]
port 26 nsew signal output
flabel metal2 s 7930 3000 7986 3400 0 FreeSans 224 90 0 0 HI[34]
port 27 nsew signal output
flabel metal2 s 8114 3000 8170 3400 0 FreeSans 224 90 0 0 HI[35]
port 28 nsew signal output
flabel metal2 s 8298 3000 8354 3400 0 FreeSans 224 90 0 0 HI[36]
port 29 nsew signal output
flabel metal2 s 8482 3000 8538 3400 0 FreeSans 224 90 0 0 HI[37]
port 30 nsew signal output
flabel metal2 s 8666 3000 8722 3400 0 FreeSans 224 90 0 0 HI[38]
port 31 nsew signal output
flabel metal2 s 8850 3000 8906 3400 0 FreeSans 224 90 0 0 HI[39]
port 32 nsew signal output
flabel metal2 s 2226 3000 2282 3400 0 FreeSans 224 90 0 0 HI[3]
port 33 nsew signal output
flabel metal2 s 9034 3000 9090 3400 0 FreeSans 224 90 0 0 HI[40]
port 34 nsew signal output
flabel metal2 s 9218 3000 9274 3400 0 FreeSans 224 90 0 0 HI[41]
port 35 nsew signal output
flabel metal2 s 9402 3000 9458 3400 0 FreeSans 224 90 0 0 HI[42]
port 36 nsew signal output
flabel metal2 s 9586 3000 9642 3400 0 FreeSans 224 90 0 0 HI[43]
port 37 nsew signal output
flabel metal2 s 9770 3000 9826 3400 0 FreeSans 224 90 0 0 HI[44]
port 38 nsew signal output
flabel metal2 s 9954 3000 10010 3400 0 FreeSans 224 90 0 0 HI[45]
port 39 nsew signal output
flabel metal2 s 10138 3000 10194 3400 0 FreeSans 224 90 0 0 HI[46]
port 40 nsew signal output
flabel metal2 s 10322 3000 10378 3400 0 FreeSans 224 90 0 0 HI[47]
port 41 nsew signal output
flabel metal2 s 10506 3000 10562 3400 0 FreeSans 224 90 0 0 HI[48]
port 42 nsew signal output
flabel metal2 s 10690 3000 10746 3400 0 FreeSans 224 90 0 0 HI[49]
port 43 nsew signal output
flabel metal2 s 2410 3000 2466 3400 0 FreeSans 224 90 0 0 HI[4]
port 44 nsew signal output
flabel metal2 s 10874 3000 10930 3400 0 FreeSans 224 90 0 0 HI[50]
port 45 nsew signal output
flabel metal2 s 11058 3000 11114 3400 0 FreeSans 224 90 0 0 HI[51]
port 46 nsew signal output
flabel metal2 s 11242 3000 11298 3400 0 FreeSans 224 90 0 0 HI[52]
port 47 nsew signal output
flabel metal2 s 11426 3000 11482 3400 0 FreeSans 224 90 0 0 HI[53]
port 48 nsew signal output
flabel metal2 s 11610 3000 11666 3400 0 FreeSans 224 90 0 0 HI[54]
port 49 nsew signal output
flabel metal2 s 11794 3000 11850 3400 0 FreeSans 224 90 0 0 HI[55]
port 50 nsew signal output
flabel metal2 s 11978 3000 12034 3400 0 FreeSans 224 90 0 0 HI[56]
port 51 nsew signal output
flabel metal2 s 12162 3000 12218 3400 0 FreeSans 224 90 0 0 HI[57]
port 52 nsew signal output
flabel metal2 s 12346 3000 12402 3400 0 FreeSans 224 90 0 0 HI[58]
port 53 nsew signal output
flabel metal2 s 12530 3000 12586 3400 0 FreeSans 224 90 0 0 HI[59]
port 54 nsew signal output
flabel metal2 s 2594 3000 2650 3400 0 FreeSans 224 90 0 0 HI[5]
port 55 nsew signal output
flabel metal2 s 12714 3000 12770 3400 0 FreeSans 224 90 0 0 HI[60]
port 56 nsew signal output
flabel metal2 s 12898 3000 12954 3400 0 FreeSans 224 90 0 0 HI[61]
port 57 nsew signal output
flabel metal2 s 13082 3000 13138 3400 0 FreeSans 224 90 0 0 HI[62]
port 58 nsew signal output
flabel metal2 s 13266 3000 13322 3400 0 FreeSans 224 90 0 0 HI[63]
port 59 nsew signal output
flabel metal2 s 13450 3000 13506 3400 0 FreeSans 224 90 0 0 HI[64]
port 60 nsew signal output
flabel metal2 s 13634 3000 13690 3400 0 FreeSans 224 90 0 0 HI[65]
port 61 nsew signal output
flabel metal2 s 13818 3000 13874 3400 0 FreeSans 224 90 0 0 HI[66]
port 62 nsew signal output
flabel metal2 s 14002 3000 14058 3400 0 FreeSans 224 90 0 0 HI[67]
port 63 nsew signal output
flabel metal2 s 14186 3000 14242 3400 0 FreeSans 224 90 0 0 HI[68]
port 64 nsew signal output
flabel metal2 s 14370 3000 14426 3400 0 FreeSans 224 90 0 0 HI[69]
port 65 nsew signal output
flabel metal2 s 2778 3000 2834 3400 0 FreeSans 224 90 0 0 HI[6]
port 66 nsew signal output
flabel metal2 s 14554 3000 14610 3400 0 FreeSans 224 90 0 0 HI[70]
port 67 nsew signal output
flabel metal2 s 14738 3000 14794 3400 0 FreeSans 224 90 0 0 HI[71]
port 68 nsew signal output
flabel metal2 s 14922 3000 14978 3400 0 FreeSans 224 90 0 0 HI[72]
port 69 nsew signal output
flabel metal2 s 15106 3000 15162 3400 0 FreeSans 224 90 0 0 HI[73]
port 70 nsew signal output
flabel metal2 s 15290 3000 15346 3400 0 FreeSans 224 90 0 0 HI[74]
port 71 nsew signal output
flabel metal2 s 15474 3000 15530 3400 0 FreeSans 224 90 0 0 HI[75]
port 72 nsew signal output
flabel metal2 s 15658 3000 15714 3400 0 FreeSans 224 90 0 0 HI[76]
port 73 nsew signal output
flabel metal2 s 15842 3000 15898 3400 0 FreeSans 224 90 0 0 HI[77]
port 74 nsew signal output
flabel metal2 s 16026 3000 16082 3400 0 FreeSans 224 90 0 0 HI[78]
port 75 nsew signal output
flabel metal2 s 16210 3000 16266 3400 0 FreeSans 224 90 0 0 HI[79]
port 76 nsew signal output
flabel metal2 s 2962 3000 3018 3400 0 FreeSans 224 90 0 0 HI[7]
port 77 nsew signal output
flabel metal2 s 16394 3000 16450 3400 0 FreeSans 224 90 0 0 HI[80]
port 78 nsew signal output
flabel metal2 s 16578 3000 16634 3400 0 FreeSans 224 90 0 0 HI[81]
port 79 nsew signal output
flabel metal2 s 16762 3000 16818 3400 0 FreeSans 224 90 0 0 HI[82]
port 80 nsew signal output
flabel metal2 s 16946 3000 17002 3400 0 FreeSans 224 90 0 0 HI[83]
port 81 nsew signal output
flabel metal2 s 17130 3000 17186 3400 0 FreeSans 224 90 0 0 HI[84]
port 82 nsew signal output
flabel metal2 s 17314 3000 17370 3400 0 FreeSans 224 90 0 0 HI[85]
port 83 nsew signal output
flabel metal2 s 17498 3000 17554 3400 0 FreeSans 224 90 0 0 HI[86]
port 84 nsew signal output
flabel metal2 s 17682 3000 17738 3400 0 FreeSans 224 90 0 0 HI[87]
port 85 nsew signal output
flabel metal2 s 17866 3000 17922 3400 0 FreeSans 224 90 0 0 HI[88]
port 86 nsew signal output
flabel metal2 s 18050 3000 18106 3400 0 FreeSans 224 90 0 0 HI[89]
port 87 nsew signal output
flabel metal2 s 3146 3000 3202 3400 0 FreeSans 224 90 0 0 HI[8]
port 88 nsew signal output
flabel metal2 s 18234 3000 18290 3400 0 FreeSans 224 90 0 0 HI[90]
port 89 nsew signal output
flabel metal2 s 3330 3000 3386 3400 0 FreeSans 224 90 0 0 HI[9]
port 90 nsew signal output
flabel metal2 s 1116 496 1436 2224 0 FreeSans 1792 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal2 s 9116 496 9436 2224 0 FreeSans 1792 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal2 s 17116 496 17436 2224 0 FreeSans 1792 90 0 0 vccd1
port 91 nsew power bidirectional
flabel metal3 s 228 880 19828 1200 0 FreeSans 1920 0 0 0 vccd1
port 91 nsew power bidirectional
flabel metal2 s 1756 496 2076 2224 0 FreeSans 1792 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal2 s 9756 496 10076 2224 0 FreeSans 1792 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal2 s 17756 496 18076 2224 0 FreeSans 1792 90 0 0 vssd1
port 92 nsew ground bidirectional
flabel metal3 s 228 1520 19828 1840 0 FreeSans 1920 0 0 0 vssd1
port 92 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 20000 3400
<< end >>
