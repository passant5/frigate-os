magic
tech sky130A
magscale 1 2
timestamp 1750117369
<< viali >>
rect 5549 13957 5583 13991
rect 1685 13889 1719 13923
rect 2605 13889 2639 13923
rect 3341 13889 3375 13923
rect 3617 13889 3651 13923
rect 4445 13889 4479 13923
rect 6837 13889 6871 13923
rect 8125 13889 8159 13923
rect 8493 13889 8527 13923
rect 8677 13889 8711 13923
rect 1777 13821 1811 13855
rect 4261 13821 4295 13855
rect 6561 13821 6595 13855
rect 7849 13821 7883 13855
rect 3157 13753 3191 13787
rect 1041 13685 1075 13719
rect 2421 13685 2455 13719
rect 3525 13685 3559 13719
rect 5917 13685 5951 13719
rect 6653 13685 6687 13719
rect 8861 13685 8895 13719
rect 4721 13345 4755 13379
rect 5365 13345 5399 13379
rect 6377 13345 6411 13379
rect 949 13277 983 13311
rect 1225 13277 1259 13311
rect 1501 13277 1535 13311
rect 1869 13277 1903 13311
rect 2513 13277 2547 13311
rect 3157 13277 3191 13311
rect 3709 13277 3743 13311
rect 4629 13277 4663 13311
rect 6653 13277 6687 13311
rect 7113 13277 7147 13311
rect 8677 13277 8711 13311
rect 8861 13277 8895 13311
rect 3525 13209 3559 13243
rect 3893 13209 3927 13243
rect 8125 13209 8159 13243
rect 1133 13141 1167 13175
rect 1409 13141 1443 13175
rect 1685 13141 1719 13175
rect 2421 13141 2455 13175
rect 3985 13141 4019 13175
rect 8493 13141 8527 13175
rect 949 12801 983 12835
rect 3249 12801 3283 12835
rect 5089 12801 5123 12835
rect 6192 12801 6226 12835
rect 6285 12801 6319 12835
rect 8401 12801 8435 12835
rect 1409 12733 1443 12767
rect 2513 12733 2547 12767
rect 3157 12733 3191 12767
rect 3617 12733 3651 12767
rect 6561 12733 6595 12767
rect 6929 12733 6963 12767
rect 5653 12597 5687 12631
rect 6101 12597 6135 12631
rect 8961 12597 8995 12631
rect 1225 12393 1259 12427
rect 1409 12393 1443 12427
rect 7121 12393 7155 12427
rect 3893 12325 3927 12359
rect 7297 12325 7331 12359
rect 3157 12257 3191 12291
rect 4537 12257 4571 12291
rect 8125 12257 8159 12291
rect 1133 12189 1167 12223
rect 3525 12189 3559 12223
rect 3679 12189 3713 12223
rect 4721 12189 4755 12223
rect 5089 12189 5123 12223
rect 6561 12189 6595 12223
rect 7849 12189 7883 12223
rect 8033 12189 8067 12223
rect 8768 12189 8802 12223
rect 8861 12189 8895 12223
rect 2881 12121 2915 12155
rect 3985 12121 4019 12155
rect 8493 12053 8527 12087
rect 949 11849 983 11883
rect 6285 11849 6319 11883
rect 8777 11849 8811 11883
rect 3065 11781 3099 11815
rect 2697 11713 2731 11747
rect 2789 11713 2823 11747
rect 5549 11713 5583 11747
rect 5917 11713 5951 11747
rect 6010 11713 6044 11747
rect 6377 11713 6411 11747
rect 8217 11713 8251 11747
rect 2421 11645 2455 11679
rect 4537 11645 4571 11679
rect 4813 11645 4847 11679
rect 6745 11645 6779 11679
rect 5733 11577 5767 11611
rect 5457 11509 5491 11543
rect 3065 11305 3099 11339
rect 6837 11305 6871 11339
rect 2329 11237 2363 11271
rect 2789 11169 2823 11203
rect 3525 11169 3559 11203
rect 3893 11169 3927 11203
rect 2145 11101 2179 11135
rect 2421 11101 2455 11135
rect 2697 11101 2731 11135
rect 2973 11101 3007 11135
rect 5365 11101 5399 11135
rect 6285 11101 6319 11135
rect 6929 11101 6963 11135
rect 8861 11101 8895 11135
rect 1041 11033 1075 11067
rect 1869 11033 1903 11067
rect 5929 11033 5963 11067
rect 8125 11033 8159 11067
rect 8677 11033 8711 11067
rect 2605 10965 2639 10999
rect 8493 10965 8527 10999
rect 4537 10761 4571 10795
rect 5273 10761 5307 10795
rect 6469 10761 6503 10795
rect 1041 10693 1075 10727
rect 1869 10693 1903 10727
rect 5641 10693 5675 10727
rect 6101 10693 6135 10727
rect 5457 10625 5491 10659
rect 6285 10625 6319 10659
rect 8401 10625 8435 10659
rect 1961 10557 1995 10591
rect 2237 10557 2271 10591
rect 3801 10557 3835 10591
rect 5089 10557 5123 10591
rect 6561 10557 6595 10591
rect 6929 10557 6963 10591
rect 3709 10489 3743 10523
rect 4445 10421 4479 10455
rect 8961 10421 8995 10455
rect 2053 10217 2087 10251
rect 2513 10217 2547 10251
rect 3341 10217 3375 10251
rect 5733 10217 5767 10251
rect 5181 10149 5215 10183
rect 8493 10149 8527 10183
rect 1041 10081 1075 10115
rect 7849 10081 7883 10115
rect 2237 10013 2271 10047
rect 3065 10013 3099 10047
rect 5089 10013 5123 10047
rect 5456 10013 5490 10047
rect 5549 10013 5583 10047
rect 5641 10013 5675 10047
rect 5917 10013 5951 10047
rect 6837 10013 6871 10047
rect 8309 10013 8343 10047
rect 8768 10013 8802 10047
rect 8861 10013 8895 10047
rect 1869 9945 1903 9979
rect 4813 9945 4847 9979
rect 6745 9945 6779 9979
rect 6561 9877 6595 9911
rect 5733 9673 5767 9707
rect 4261 9605 4295 9639
rect 6009 9605 6043 9639
rect 6193 9605 6227 9639
rect 1041 9537 1075 9571
rect 2973 9537 3007 9571
rect 3433 9537 3467 9571
rect 3525 9537 3559 9571
rect 6377 9537 6411 9571
rect 8217 9537 8251 9571
rect 1317 9469 1351 9503
rect 3341 9469 3375 9503
rect 3985 9469 4019 9503
rect 6745 9469 6779 9503
rect 2789 9401 2823 9435
rect 3157 9333 3191 9367
rect 3709 9333 3743 9367
rect 8777 9333 8811 9367
rect 7389 9129 7423 9163
rect 2973 9061 3007 9095
rect 4997 9061 5031 9095
rect 8493 9061 8527 9095
rect 6745 8993 6779 9027
rect 2145 8925 2179 8959
rect 2727 8925 2761 8959
rect 2881 8925 2915 8959
rect 3157 8925 3191 8959
rect 3341 8925 3375 8959
rect 3617 8925 3651 8959
rect 6837 8925 6871 8959
rect 6991 8925 7025 8959
rect 7481 8925 7515 8959
rect 7665 8925 7699 8959
rect 8737 8925 8771 8959
rect 8861 8925 8895 8959
rect 1133 8857 1167 8891
rect 6469 8857 6503 8891
rect 2513 8789 2547 8823
rect 3525 8789 3559 8823
rect 3801 8789 3835 8823
rect 7205 8789 7239 8823
rect 8217 8789 8251 8823
rect 3893 8517 3927 8551
rect 1041 8449 1075 8483
rect 1685 8449 1719 8483
rect 3157 8449 3191 8483
rect 4077 8449 4111 8483
rect 6377 8449 6411 8483
rect 8953 8449 8987 8483
rect 1133 8381 1167 8415
rect 1317 8381 1351 8415
rect 4261 8381 4295 8415
rect 6745 8381 6779 8415
rect 8585 8381 8619 8415
rect 6193 8313 6227 8347
rect 3717 8245 3751 8279
rect 6653 8245 6687 8279
rect 7389 8245 7423 8279
rect 1777 8041 1811 8075
rect 8493 8041 8527 8075
rect 2605 7973 2639 8007
rect 1225 7905 1259 7939
rect 2053 7905 2087 7939
rect 7849 7905 7883 7939
rect 1409 7837 1443 7871
rect 4077 7837 4111 7871
rect 6101 7837 6135 7871
rect 8309 7837 8343 7871
rect 8861 7837 8895 7871
rect 2145 7769 2179 7803
rect 5641 7769 5675 7803
rect 5825 7769 5859 7803
rect 6745 7769 6779 7803
rect 8677 7769 8711 7803
rect 1317 7701 1351 7735
rect 2237 7701 2271 7735
rect 4721 7701 4755 7735
rect 6009 7701 6043 7735
rect 1133 7497 1167 7531
rect 1409 7497 1443 7531
rect 3157 7497 3191 7531
rect 8501 7497 8535 7531
rect 4629 7429 4663 7463
rect 8677 7429 8711 7463
rect 949 7361 983 7395
rect 1225 7361 1259 7395
rect 4905 7361 4939 7395
rect 5089 7361 5123 7395
rect 5640 7361 5674 7395
rect 5733 7361 5767 7395
rect 6469 7361 6503 7395
rect 7941 7361 7975 7395
rect 8861 7361 8895 7395
rect 2237 7293 2271 7327
rect 2789 7293 2823 7327
rect 5181 7293 5215 7327
rect 6101 7293 6135 7327
rect 9045 7293 9079 7327
rect 5549 7157 5583 7191
rect 7297 6953 7331 6987
rect 8309 6953 8343 6987
rect 6941 6885 6975 6919
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 4537 6749 4571 6783
rect 4905 6749 4939 6783
rect 6377 6749 6411 6783
rect 7849 6749 7883 6783
rect 8125 6749 8159 6783
rect 8707 6749 8741 6783
rect 8861 6749 8895 6783
rect 8493 6613 8527 6647
rect 1133 6409 1167 6443
rect 949 6273 983 6307
rect 6009 6273 6043 6307
rect 6285 6273 6319 6307
rect 8401 6273 8435 6307
rect 3893 6205 3927 6239
rect 4169 6205 4203 6239
rect 5641 6205 5675 6239
rect 6377 6205 6411 6239
rect 6561 6205 6595 6239
rect 6929 6205 6963 6239
rect 6193 6069 6227 6103
rect 8961 6069 8995 6103
rect 6561 5865 6595 5899
rect 8493 5865 8527 5899
rect 6653 5797 6687 5831
rect 1409 5729 1443 5763
rect 4813 5729 4847 5763
rect 5089 5729 5123 5763
rect 7849 5729 7883 5763
rect 1133 5661 1167 5695
rect 6837 5661 6871 5695
rect 8309 5661 8343 5695
rect 8861 5661 8895 5695
rect 8677 5593 8711 5627
rect 5733 5321 5767 5355
rect 8861 5253 8895 5287
rect 6377 5185 6411 5219
rect 7665 5185 7699 5219
rect 949 5117 983 5151
rect 1225 5117 1259 5151
rect 2697 5117 2731 5151
rect 5089 5117 5123 5151
rect 7389 5117 7423 5151
rect 1133 4777 1167 4811
rect 2145 4709 2179 4743
rect 4261 4641 4295 4675
rect 4905 4641 4939 4675
rect 6653 4641 6687 4675
rect 7849 4641 7883 4675
rect 949 4573 983 4607
rect 1409 4573 1443 4607
rect 8309 4573 8343 4607
rect 8707 4573 8741 4607
rect 8861 4573 8895 4607
rect 1961 4505 1995 4539
rect 6377 4505 6411 4539
rect 1225 4437 1259 4471
rect 4813 4437 4847 4471
rect 8493 4437 8527 4471
rect 6285 4233 6319 4267
rect 8961 4233 8995 4267
rect 3709 4097 3743 4131
rect 5549 4097 5583 4131
rect 6101 4097 6135 4131
rect 6929 4097 6963 4131
rect 8401 4097 8435 4131
rect 3985 4029 4019 4063
rect 5641 4029 5675 4063
rect 6561 4029 6595 4063
rect 5457 3893 5491 3927
rect 3985 3689 4019 3723
rect 8493 3689 8527 3723
rect 7665 3621 7699 3655
rect 5733 3553 5767 3587
rect 5917 3553 5951 3587
rect 6193 3553 6227 3587
rect 7849 3485 7883 3519
rect 7941 3485 7975 3519
rect 8861 3485 8895 3519
rect 5457 3417 5491 3451
rect 8677 3417 8711 3451
rect 8493 3077 8527 3111
rect 4997 3009 5031 3043
rect 5168 3009 5202 3043
rect 5733 3009 5767 3043
rect 7205 3009 7239 3043
rect 7573 3009 7607 3043
rect 8677 3009 8711 3043
rect 4537 2941 4571 2975
rect 7757 2941 7791 2975
rect 8309 2941 8343 2975
rect 8861 2805 8895 2839
rect 2789 2601 2823 2635
rect 5825 2601 5859 2635
rect 8769 2601 8803 2635
rect 4905 2465 4939 2499
rect 6009 2465 6043 2499
rect 6377 2465 6411 2499
rect 2973 2397 3007 2431
rect 3065 2397 3099 2431
rect 4813 2397 4847 2431
rect 5273 2397 5307 2431
rect 7849 2397 7883 2431
rect 8585 2397 8619 2431
rect 8739 2397 8773 2431
rect 8409 2261 8443 2295
rect 7205 2057 7239 2091
rect 5181 1989 5215 2023
rect 8677 1989 8711 2023
rect 4721 1921 4755 1955
rect 4905 1921 4939 1955
rect 6837 1921 6871 1955
rect 6930 1921 6964 1955
rect 8861 1921 8895 1955
rect 4353 1853 4387 1887
rect 6653 1785 6687 1819
rect 9045 1717 9079 1751
rect 8861 1513 8895 1547
rect 7389 1377 7423 1411
rect 6377 1309 6411 1343
rect 9045 1309 9079 1343
<< metal1 >>
rect 5350 14288 5356 14340
rect 5408 14328 5414 14340
rect 7098 14328 7104 14340
rect 5408 14300 7104 14328
rect 5408 14288 5414 14300
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 8018 14260 8024 14272
rect 3292 14232 8024 14260
rect 3292 14220 3298 14232
rect 8018 14220 8024 14232
rect 8076 14220 8082 14272
rect 644 14170 9384 14192
rect 644 14118 2954 14170
rect 3006 14118 3018 14170
rect 3070 14118 3082 14170
rect 3134 14118 6954 14170
rect 7006 14118 7018 14170
rect 7070 14118 7082 14170
rect 7134 14118 9384 14170
rect 644 14096 9384 14118
rect 6822 14056 6828 14068
rect 1596 14028 6828 14056
rect 1596 13852 1624 14028
rect 6822 14016 6828 14028
rect 6880 14016 6886 14068
rect 4798 13988 4804 14000
rect 1688 13960 4804 13988
rect 1688 13929 1716 13960
rect 4798 13948 4804 13960
rect 4856 13948 4862 14000
rect 5537 13991 5595 13997
rect 5537 13957 5549 13991
rect 5583 13988 5595 13991
rect 9582 13988 9588 14000
rect 5583 13960 9588 13988
rect 5583 13957 5595 13960
rect 5537 13951 5595 13957
rect 9582 13948 9588 13960
rect 9640 13948 9646 14000
rect 1673 13923 1731 13929
rect 1673 13889 1685 13923
rect 1719 13889 1731 13923
rect 1673 13883 1731 13889
rect 2593 13923 2651 13929
rect 2593 13889 2605 13923
rect 2639 13920 2651 13923
rect 3234 13920 3240 13932
rect 2639 13892 3240 13920
rect 2639 13889 2651 13892
rect 2593 13883 2651 13889
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 3329 13923 3387 13929
rect 3329 13889 3341 13923
rect 3375 13920 3387 13923
rect 3605 13923 3663 13929
rect 3605 13920 3617 13923
rect 3375 13892 3617 13920
rect 3375 13889 3387 13892
rect 3329 13883 3387 13889
rect 3605 13889 3617 13892
rect 3651 13889 3663 13923
rect 3605 13883 3663 13889
rect 4430 13880 4436 13932
rect 4488 13880 4494 13932
rect 6270 13880 6276 13932
rect 6328 13920 6334 13932
rect 6825 13923 6883 13929
rect 6825 13920 6837 13923
rect 6328 13892 6837 13920
rect 6328 13880 6334 13892
rect 6825 13889 6837 13892
rect 6871 13889 6883 13923
rect 6825 13883 6883 13889
rect 8110 13880 8116 13932
rect 8168 13880 8174 13932
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13920 8539 13923
rect 8570 13920 8576 13932
rect 8527 13892 8576 13920
rect 8527 13889 8539 13892
rect 8481 13883 8539 13889
rect 8570 13880 8576 13892
rect 8628 13880 8634 13932
rect 8665 13923 8723 13929
rect 8665 13889 8677 13923
rect 8711 13889 8723 13923
rect 8665 13883 8723 13889
rect 1765 13855 1823 13861
rect 1765 13852 1777 13855
rect 1596 13824 1777 13852
rect 1765 13821 1777 13824
rect 1811 13821 1823 13855
rect 1765 13815 1823 13821
rect 4249 13855 4307 13861
rect 4249 13821 4261 13855
rect 4295 13852 4307 13855
rect 6454 13852 6460 13864
rect 4295 13824 6460 13852
rect 4295 13821 4307 13824
rect 4249 13815 4307 13821
rect 6454 13812 6460 13824
rect 6512 13812 6518 13864
rect 6549 13855 6607 13861
rect 6549 13821 6561 13855
rect 6595 13821 6607 13855
rect 6549 13815 6607 13821
rect 7837 13855 7895 13861
rect 7837 13821 7849 13855
rect 7883 13852 7895 13855
rect 8680 13852 8708 13883
rect 7883 13824 8524 13852
rect 7883 13821 7895 13824
rect 7837 13815 7895 13821
rect 3145 13787 3203 13793
rect 3145 13753 3157 13787
rect 3191 13784 3203 13787
rect 3970 13784 3976 13796
rect 3191 13756 3976 13784
rect 3191 13753 3203 13756
rect 3145 13747 3203 13753
rect 3970 13744 3976 13756
rect 4028 13744 4034 13796
rect 5626 13744 5632 13796
rect 5684 13784 5690 13796
rect 6564 13784 6592 13815
rect 8496 13796 8524 13824
rect 8588 13824 8708 13852
rect 5684 13756 6040 13784
rect 6564 13756 7236 13784
rect 5684 13744 5690 13756
rect 934 13676 940 13728
rect 992 13716 998 13728
rect 1029 13719 1087 13725
rect 1029 13716 1041 13719
rect 992 13688 1041 13716
rect 992 13676 998 13688
rect 1029 13685 1041 13688
rect 1075 13685 1087 13719
rect 1029 13679 1087 13685
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 2409 13719 2467 13725
rect 2409 13716 2421 13719
rect 1728 13688 2421 13716
rect 1728 13676 1734 13688
rect 2409 13685 2421 13688
rect 2455 13685 2467 13719
rect 2409 13679 2467 13685
rect 3513 13719 3571 13725
rect 3513 13685 3525 13719
rect 3559 13716 3571 13719
rect 4890 13716 4896 13728
rect 3559 13688 4896 13716
rect 3559 13685 3571 13688
rect 3513 13679 3571 13685
rect 4890 13676 4896 13688
rect 4948 13676 4954 13728
rect 5902 13676 5908 13728
rect 5960 13676 5966 13728
rect 6012 13716 6040 13756
rect 7208 13728 7236 13756
rect 8478 13744 8484 13796
rect 8536 13744 8542 13796
rect 8588 13728 8616 13824
rect 6641 13719 6699 13725
rect 6641 13716 6653 13719
rect 6012 13688 6653 13716
rect 6641 13685 6653 13688
rect 6687 13685 6699 13719
rect 6641 13679 6699 13685
rect 7190 13676 7196 13728
rect 7248 13676 7254 13728
rect 8570 13676 8576 13728
rect 8628 13676 8634 13728
rect 8846 13676 8852 13728
rect 8904 13676 8910 13728
rect 644 13626 9384 13648
rect 644 13574 2554 13626
rect 2606 13574 2618 13626
rect 2670 13574 2682 13626
rect 2734 13574 6554 13626
rect 6606 13574 6618 13626
rect 6670 13574 6682 13626
rect 6734 13574 9384 13626
rect 644 13552 9384 13574
rect 1854 13472 1860 13524
rect 1912 13512 1918 13524
rect 5718 13512 5724 13524
rect 1912 13484 5724 13512
rect 1912 13472 1918 13484
rect 5718 13472 5724 13484
rect 5776 13472 5782 13524
rect 6178 13472 6184 13524
rect 6236 13512 6242 13524
rect 8846 13512 8852 13524
rect 6236 13484 8852 13512
rect 6236 13472 6242 13484
rect 8846 13472 8852 13484
rect 8904 13472 8910 13524
rect 5902 13444 5908 13456
rect 2746 13416 5908 13444
rect 2746 13376 2774 13416
rect 5902 13404 5908 13416
rect 5960 13404 5966 13456
rect 7650 13444 7656 13456
rect 6196 13416 7656 13444
rect 4709 13379 4767 13385
rect 4709 13376 4721 13379
rect 1228 13348 2774 13376
rect 3436 13348 4721 13376
rect 934 13268 940 13320
rect 992 13268 998 13320
rect 1228 13317 1256 13348
rect 1213 13311 1271 13317
rect 1213 13277 1225 13311
rect 1259 13277 1271 13311
rect 1213 13271 1271 13277
rect 1489 13311 1547 13317
rect 1489 13277 1501 13311
rect 1535 13277 1547 13311
rect 1489 13271 1547 13277
rect 1504 13240 1532 13271
rect 1854 13268 1860 13320
rect 1912 13268 1918 13320
rect 2406 13268 2412 13320
rect 2464 13308 2470 13320
rect 2501 13311 2559 13317
rect 2501 13308 2513 13311
rect 2464 13280 2513 13308
rect 2464 13268 2470 13280
rect 2501 13277 2513 13280
rect 2547 13277 2559 13311
rect 2501 13271 2559 13277
rect 3145 13311 3203 13317
rect 3145 13277 3157 13311
rect 3191 13308 3203 13311
rect 3234 13308 3240 13320
rect 3191 13280 3240 13308
rect 3191 13277 3203 13280
rect 3145 13271 3203 13277
rect 3234 13268 3240 13280
rect 3292 13268 3298 13320
rect 3436 13240 3464 13348
rect 4709 13345 4721 13348
rect 4755 13345 4767 13379
rect 4709 13339 4767 13345
rect 5350 13336 5356 13388
rect 5408 13336 5414 13388
rect 3697 13311 3755 13317
rect 3697 13277 3709 13311
rect 3743 13308 3755 13311
rect 4522 13308 4528 13320
rect 3743 13280 4528 13308
rect 3743 13277 3755 13280
rect 3697 13271 3755 13277
rect 4522 13268 4528 13280
rect 4580 13268 4586 13320
rect 4617 13311 4675 13317
rect 4617 13277 4629 13311
rect 4663 13308 4675 13311
rect 6196 13308 6224 13416
rect 7650 13404 7656 13416
rect 7708 13404 7714 13456
rect 9582 13444 9588 13456
rect 8496 13416 9588 13444
rect 6365 13379 6423 13385
rect 6365 13345 6377 13379
rect 6411 13376 6423 13379
rect 8496 13376 8524 13416
rect 9582 13404 9588 13416
rect 9640 13404 9646 13456
rect 6411 13348 8524 13376
rect 6411 13345 6423 13348
rect 6365 13339 6423 13345
rect 8570 13336 8576 13388
rect 8628 13336 8634 13388
rect 4663 13280 6224 13308
rect 4663 13277 4675 13280
rect 4617 13271 4675 13277
rect 6454 13268 6460 13320
rect 6512 13308 6518 13320
rect 6641 13311 6699 13317
rect 6641 13308 6653 13311
rect 6512 13280 6653 13308
rect 6512 13268 6518 13280
rect 6641 13277 6653 13280
rect 6687 13277 6699 13311
rect 6641 13271 6699 13277
rect 7101 13311 7159 13317
rect 7101 13277 7113 13311
rect 7147 13308 7159 13311
rect 7650 13308 7656 13320
rect 7147 13280 7656 13308
rect 7147 13277 7159 13280
rect 7101 13271 7159 13277
rect 7650 13268 7656 13280
rect 7708 13268 7714 13320
rect 8588 13308 8616 13336
rect 8665 13311 8723 13317
rect 8665 13308 8677 13311
rect 7760 13280 8677 13308
rect 1504 13212 3464 13240
rect 3513 13243 3571 13249
rect 3513 13209 3525 13243
rect 3559 13209 3571 13243
rect 3513 13203 3571 13209
rect 3881 13243 3939 13249
rect 3881 13209 3893 13243
rect 3927 13240 3939 13243
rect 5074 13240 5080 13252
rect 3927 13212 5080 13240
rect 3927 13209 3939 13212
rect 3881 13203 3939 13209
rect 1118 13132 1124 13184
rect 1176 13132 1182 13184
rect 1394 13132 1400 13184
rect 1452 13132 1458 13184
rect 1578 13132 1584 13184
rect 1636 13172 1642 13184
rect 1673 13175 1731 13181
rect 1673 13172 1685 13175
rect 1636 13144 1685 13172
rect 1636 13132 1642 13144
rect 1673 13141 1685 13144
rect 1719 13141 1731 13175
rect 1673 13135 1731 13141
rect 2038 13132 2044 13184
rect 2096 13172 2102 13184
rect 2409 13175 2467 13181
rect 2409 13172 2421 13175
rect 2096 13144 2421 13172
rect 2096 13132 2102 13144
rect 2409 13141 2421 13144
rect 2455 13141 2467 13175
rect 2409 13135 2467 13141
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 3528 13172 3556 13203
rect 5074 13200 5080 13212
rect 5132 13200 5138 13252
rect 6362 13200 6368 13252
rect 6420 13240 6426 13252
rect 7760 13240 7788 13280
rect 8665 13277 8677 13280
rect 8711 13277 8723 13311
rect 8665 13271 8723 13277
rect 6420 13212 7788 13240
rect 8113 13243 8171 13249
rect 6420 13200 6426 13212
rect 8113 13209 8125 13243
rect 8159 13240 8171 13243
rect 8570 13240 8576 13252
rect 8159 13212 8576 13240
rect 8159 13209 8171 13212
rect 8113 13203 8171 13209
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 8680 13240 8708 13271
rect 8846 13268 8852 13320
rect 8904 13268 8910 13320
rect 9122 13240 9128 13252
rect 8680 13212 9128 13240
rect 9122 13200 9128 13212
rect 9180 13200 9186 13252
rect 2832 13144 3556 13172
rect 3973 13175 4031 13181
rect 2832 13132 2838 13144
rect 3973 13141 3985 13175
rect 4019 13172 4031 13175
rect 4062 13172 4068 13184
rect 4019 13144 4068 13172
rect 4019 13141 4031 13144
rect 3973 13135 4031 13141
rect 4062 13132 4068 13144
rect 4120 13132 4126 13184
rect 8202 13132 8208 13184
rect 8260 13172 8266 13184
rect 8481 13175 8539 13181
rect 8481 13172 8493 13175
rect 8260 13144 8493 13172
rect 8260 13132 8266 13144
rect 8481 13141 8493 13144
rect 8527 13141 8539 13175
rect 8481 13135 8539 13141
rect 644 13082 9384 13104
rect 644 13030 2954 13082
rect 3006 13030 3018 13082
rect 3070 13030 3082 13082
rect 3134 13030 6954 13082
rect 7006 13030 7018 13082
rect 7070 13030 7082 13082
rect 7134 13030 9384 13082
rect 644 13008 9384 13030
rect 2884 12940 3188 12968
rect 934 12792 940 12844
rect 992 12792 998 12844
rect 1210 12792 1216 12844
rect 1268 12832 1274 12844
rect 1268 12828 2820 12832
rect 2884 12828 2912 12940
rect 1268 12804 2912 12828
rect 3160 12832 3188 12940
rect 3234 12928 3240 12980
rect 3292 12968 3298 12980
rect 8294 12968 8300 12980
rect 3292 12940 8300 12968
rect 3292 12928 3298 12940
rect 8294 12928 8300 12940
rect 8352 12928 8358 12980
rect 4154 12860 4160 12912
rect 4212 12860 4218 12912
rect 6362 12900 6368 12912
rect 5000 12872 6368 12900
rect 3237 12835 3295 12841
rect 3237 12832 3249 12835
rect 3160 12804 3249 12832
rect 1268 12792 1274 12804
rect 2792 12800 2912 12804
rect 3237 12801 3249 12804
rect 3283 12801 3295 12835
rect 3237 12795 3295 12801
rect 4522 12792 4528 12844
rect 4580 12832 4586 12844
rect 5000 12832 5028 12872
rect 4580 12804 5028 12832
rect 4580 12792 4586 12804
rect 5074 12792 5080 12844
rect 5132 12792 5138 12844
rect 6288 12841 6316 12872
rect 6362 12860 6368 12872
rect 6420 12860 6426 12912
rect 7650 12860 7656 12912
rect 7708 12860 7714 12912
rect 6180 12835 6238 12841
rect 6180 12801 6192 12835
rect 6226 12801 6238 12835
rect 6180 12795 6238 12801
rect 6273 12835 6331 12841
rect 6273 12801 6285 12835
rect 6319 12801 6331 12835
rect 6273 12795 6331 12801
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 1486 12724 1492 12776
rect 1544 12764 1550 12776
rect 2501 12767 2559 12773
rect 2501 12764 2513 12767
rect 1544 12736 2513 12764
rect 1544 12724 1550 12736
rect 2501 12733 2513 12736
rect 2547 12733 2559 12767
rect 2501 12727 2559 12733
rect 3145 12767 3203 12773
rect 3145 12733 3157 12767
rect 3191 12764 3203 12767
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 3191 12736 3617 12764
rect 3191 12733 3203 12736
rect 3145 12727 3203 12733
rect 3252 12708 3280 12736
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3234 12656 3240 12708
rect 3292 12656 3298 12708
rect 5641 12631 5699 12637
rect 5641 12597 5653 12631
rect 5687 12628 5699 12631
rect 5810 12628 5816 12640
rect 5687 12600 5816 12628
rect 5687 12597 5699 12600
rect 5641 12591 5699 12597
rect 5810 12588 5816 12600
rect 5868 12588 5874 12640
rect 6086 12588 6092 12640
rect 6144 12588 6150 12640
rect 6196 12628 6224 12795
rect 8386 12792 8392 12844
rect 8444 12792 8450 12844
rect 6549 12767 6607 12773
rect 6549 12733 6561 12767
rect 6595 12764 6607 12767
rect 6822 12764 6828 12776
rect 6595 12736 6828 12764
rect 6595 12733 6607 12736
rect 6549 12727 6607 12733
rect 6822 12724 6828 12736
rect 6880 12724 6886 12776
rect 6917 12767 6975 12773
rect 6917 12733 6929 12767
rect 6963 12764 6975 12767
rect 7190 12764 7196 12776
rect 6963 12736 7196 12764
rect 6963 12733 6975 12736
rect 6917 12727 6975 12733
rect 7190 12724 7196 12736
rect 7248 12724 7254 12776
rect 8662 12628 8668 12640
rect 6196 12600 8668 12628
rect 8662 12588 8668 12600
rect 8720 12588 8726 12640
rect 8938 12588 8944 12640
rect 8996 12637 9002 12640
rect 8996 12591 9007 12637
rect 8996 12588 9002 12591
rect 644 12538 9384 12560
rect 644 12486 2554 12538
rect 2606 12486 2618 12538
rect 2670 12486 2682 12538
rect 2734 12486 6554 12538
rect 6606 12486 6618 12538
rect 6670 12486 6682 12538
rect 6734 12486 9384 12538
rect 644 12464 9384 12486
rect 1210 12384 1216 12436
rect 1268 12384 1274 12436
rect 1397 12427 1455 12433
rect 1397 12393 1409 12427
rect 1443 12424 1455 12427
rect 1486 12424 1492 12436
rect 1443 12396 1492 12424
rect 1443 12393 1455 12396
rect 1397 12387 1455 12393
rect 1486 12384 1492 12396
rect 1544 12384 1550 12436
rect 2774 12384 2780 12436
rect 2832 12424 2838 12436
rect 5994 12424 6000 12436
rect 2832 12396 3740 12424
rect 2832 12384 2838 12396
rect 2406 12248 2412 12300
rect 2464 12288 2470 12300
rect 3145 12291 3203 12297
rect 3145 12288 3157 12291
rect 2464 12260 3157 12288
rect 2464 12248 2470 12260
rect 3145 12257 3157 12260
rect 3191 12257 3203 12291
rect 3145 12251 3203 12257
rect 1121 12223 1179 12229
rect 1121 12189 1133 12223
rect 1167 12220 1179 12223
rect 1394 12220 1400 12232
rect 1167 12192 1400 12220
rect 1167 12189 1179 12192
rect 1121 12183 1179 12189
rect 1394 12180 1400 12192
rect 1452 12180 1458 12232
rect 3712 12229 3740 12396
rect 4540 12396 6000 12424
rect 3881 12359 3939 12365
rect 3881 12325 3893 12359
rect 3927 12356 3939 12359
rect 4154 12356 4160 12368
rect 3927 12328 4160 12356
rect 3927 12325 3939 12328
rect 3881 12319 3939 12325
rect 4154 12316 4160 12328
rect 4212 12316 4218 12368
rect 4540 12297 4568 12396
rect 5994 12384 6000 12396
rect 6052 12384 6058 12436
rect 6270 12384 6276 12436
rect 6328 12384 6334 12436
rect 6454 12384 6460 12436
rect 6512 12424 6518 12436
rect 7109 12427 7167 12433
rect 7109 12424 7121 12427
rect 6512 12396 7121 12424
rect 6512 12384 6518 12396
rect 7109 12393 7121 12396
rect 7155 12393 7167 12427
rect 7109 12387 7167 12393
rect 6288 12356 6316 12384
rect 7285 12359 7343 12365
rect 7285 12356 7297 12359
rect 6288 12328 7297 12356
rect 7285 12325 7297 12328
rect 7331 12325 7343 12359
rect 7285 12319 7343 12325
rect 4525 12291 4583 12297
rect 4525 12257 4537 12291
rect 4571 12257 4583 12291
rect 8113 12291 8171 12297
rect 8113 12288 8125 12291
rect 4525 12251 4583 12257
rect 6656 12260 8125 12288
rect 3513 12223 3571 12229
rect 3513 12189 3525 12223
rect 3559 12189 3571 12223
rect 3513 12183 3571 12189
rect 3667 12223 3740 12229
rect 3667 12189 3679 12223
rect 3713 12220 3740 12223
rect 4246 12220 4252 12232
rect 3713 12192 4252 12220
rect 3713 12189 3725 12192
rect 3667 12183 3725 12189
rect 2314 12112 2320 12164
rect 2372 12112 2378 12164
rect 2774 12112 2780 12164
rect 2832 12152 2838 12164
rect 2869 12155 2927 12161
rect 2869 12152 2881 12155
rect 2832 12124 2881 12152
rect 2832 12112 2838 12124
rect 2869 12121 2881 12124
rect 2915 12121 2927 12155
rect 2869 12115 2927 12121
rect 3528 12084 3556 12183
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 4614 12180 4620 12232
rect 4672 12220 4678 12232
rect 4709 12223 4767 12229
rect 4709 12220 4721 12223
rect 4672 12192 4721 12220
rect 4672 12180 4678 12192
rect 4709 12189 4721 12192
rect 4755 12189 4767 12223
rect 4709 12183 4767 12189
rect 5074 12180 5080 12232
rect 5132 12180 5138 12232
rect 6270 12180 6276 12232
rect 6328 12220 6334 12232
rect 6549 12223 6607 12229
rect 6549 12220 6561 12223
rect 6328 12192 6561 12220
rect 6328 12180 6334 12192
rect 6549 12189 6561 12192
rect 6595 12189 6607 12223
rect 6549 12183 6607 12189
rect 3973 12155 4031 12161
rect 3973 12121 3985 12155
rect 4019 12152 4031 12155
rect 4154 12152 4160 12164
rect 4019 12124 4160 12152
rect 4019 12121 4031 12124
rect 3973 12115 4031 12121
rect 4154 12112 4160 12124
rect 4212 12112 4218 12164
rect 6086 12112 6092 12164
rect 6144 12112 6150 12164
rect 6362 12112 6368 12164
rect 6420 12152 6426 12164
rect 6656 12152 6684 12260
rect 8113 12257 8125 12260
rect 8159 12257 8171 12291
rect 8113 12251 8171 12257
rect 7837 12223 7895 12229
rect 7837 12189 7849 12223
rect 7883 12189 7895 12223
rect 7837 12183 7895 12189
rect 6420 12124 6684 12152
rect 6420 12112 6426 12124
rect 3602 12084 3608 12096
rect 3528 12056 3608 12084
rect 3602 12044 3608 12056
rect 3660 12084 3666 12096
rect 4522 12084 4528 12096
rect 3660 12056 4528 12084
rect 3660 12044 3666 12056
rect 4522 12044 4528 12056
rect 4580 12044 4586 12096
rect 5534 12044 5540 12096
rect 5592 12084 5598 12096
rect 7852 12084 7880 12183
rect 8018 12180 8024 12232
rect 8076 12180 8082 12232
rect 8754 12220 8760 12232
rect 8715 12192 8760 12220
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 8849 12223 8907 12229
rect 8849 12189 8861 12223
rect 8895 12220 8907 12223
rect 9122 12220 9128 12232
rect 8895 12192 9128 12220
rect 8895 12189 8907 12192
rect 8849 12183 8907 12189
rect 9122 12180 9128 12192
rect 9180 12180 9186 12232
rect 5592 12056 7880 12084
rect 5592 12044 5598 12056
rect 8478 12044 8484 12096
rect 8536 12044 8542 12096
rect 644 11994 9384 12016
rect 644 11942 2954 11994
rect 3006 11942 3018 11994
rect 3070 11942 3082 11994
rect 3134 11942 6954 11994
rect 7006 11942 7018 11994
rect 7070 11942 7082 11994
rect 7134 11942 9384 11994
rect 644 11920 9384 11942
rect 934 11840 940 11892
rect 992 11840 998 11892
rect 1670 11840 1676 11892
rect 1728 11880 1734 11892
rect 2406 11880 2412 11892
rect 1728 11852 2412 11880
rect 1728 11840 1734 11852
rect 2406 11840 2412 11852
rect 2464 11880 2470 11892
rect 2464 11852 2820 11880
rect 2464 11840 2470 11852
rect 2314 11812 2320 11824
rect 1978 11784 2320 11812
rect 2314 11772 2320 11784
rect 2372 11772 2378 11824
rect 2792 11753 2820 11852
rect 3234 11840 3240 11892
rect 3292 11840 3298 11892
rect 6273 11883 6331 11889
rect 6273 11849 6285 11883
rect 6319 11880 6331 11883
rect 7650 11880 7656 11892
rect 6319 11852 7656 11880
rect 6319 11849 6331 11852
rect 6273 11843 6331 11849
rect 7650 11840 7656 11852
rect 7708 11840 7714 11892
rect 8110 11840 8116 11892
rect 8168 11880 8174 11892
rect 8765 11883 8823 11889
rect 8765 11880 8777 11883
rect 8168 11852 8777 11880
rect 8168 11840 8174 11852
rect 8765 11849 8777 11852
rect 8811 11849 8823 11883
rect 8765 11843 8823 11849
rect 3053 11815 3111 11821
rect 3053 11781 3065 11815
rect 3099 11812 3111 11815
rect 3252 11812 3280 11840
rect 4522 11812 4528 11824
rect 3099 11784 3280 11812
rect 4278 11784 4528 11812
rect 3099 11781 3111 11784
rect 3053 11775 3111 11781
rect 4522 11772 4528 11784
rect 4580 11772 4586 11824
rect 8478 11812 8484 11824
rect 7866 11784 8484 11812
rect 8478 11772 8484 11784
rect 8536 11772 8542 11824
rect 2685 11747 2743 11753
rect 2685 11713 2697 11747
rect 2731 11713 2743 11747
rect 2685 11707 2743 11713
rect 2777 11747 2835 11753
rect 2777 11713 2789 11747
rect 2823 11713 2835 11747
rect 2777 11707 2835 11713
rect 5537 11747 5595 11753
rect 5537 11713 5549 11747
rect 5583 11713 5595 11747
rect 5537 11707 5595 11713
rect 5905 11747 5963 11753
rect 5905 11713 5917 11747
rect 5951 11713 5963 11747
rect 5905 11707 5963 11713
rect 2406 11636 2412 11688
rect 2464 11636 2470 11688
rect 2314 11500 2320 11552
rect 2372 11540 2378 11552
rect 2700 11540 2728 11707
rect 4525 11679 4583 11685
rect 4525 11645 4537 11679
rect 4571 11676 4583 11679
rect 4801 11679 4859 11685
rect 4801 11676 4813 11679
rect 4571 11648 4813 11676
rect 4571 11645 4583 11648
rect 4525 11639 4583 11645
rect 4801 11645 4813 11648
rect 4847 11645 4859 11679
rect 4801 11639 4859 11645
rect 2372 11512 2728 11540
rect 2372 11500 2378 11512
rect 3234 11500 3240 11552
rect 3292 11540 3298 11552
rect 4062 11540 4068 11552
rect 3292 11512 4068 11540
rect 3292 11500 3298 11512
rect 4062 11500 4068 11512
rect 4120 11500 4126 11552
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 5074 11540 5080 11552
rect 4764 11512 5080 11540
rect 4764 11500 4770 11512
rect 5074 11500 5080 11512
rect 5132 11540 5138 11552
rect 5445 11543 5503 11549
rect 5445 11540 5457 11543
rect 5132 11512 5457 11540
rect 5132 11500 5138 11512
rect 5445 11509 5457 11512
rect 5491 11509 5503 11543
rect 5552 11540 5580 11707
rect 5920 11676 5948 11707
rect 5994 11704 6000 11756
rect 6052 11744 6058 11756
rect 6052 11716 6097 11744
rect 6052 11704 6058 11716
rect 6362 11704 6368 11756
rect 6420 11704 6426 11756
rect 8202 11704 8208 11756
rect 8260 11704 8266 11756
rect 6086 11676 6092 11688
rect 5920 11648 6092 11676
rect 6086 11636 6092 11648
rect 6144 11636 6150 11688
rect 6454 11636 6460 11688
rect 6512 11676 6518 11688
rect 6733 11679 6791 11685
rect 6733 11676 6745 11679
rect 6512 11648 6745 11676
rect 6512 11636 6518 11648
rect 6733 11645 6745 11648
rect 6779 11645 6791 11679
rect 6733 11639 6791 11645
rect 5721 11611 5779 11617
rect 5721 11577 5733 11611
rect 5767 11608 5779 11611
rect 5994 11608 6000 11620
rect 5767 11580 6000 11608
rect 5767 11577 5779 11580
rect 5721 11571 5779 11577
rect 5994 11568 6000 11580
rect 6052 11568 6058 11620
rect 9030 11540 9036 11552
rect 5552 11512 9036 11540
rect 5445 11503 5503 11509
rect 9030 11500 9036 11512
rect 9088 11500 9094 11552
rect 644 11450 9384 11472
rect 644 11398 2554 11450
rect 2606 11398 2618 11450
rect 2670 11398 2682 11450
rect 2734 11398 6554 11450
rect 6606 11398 6618 11450
rect 6670 11398 6682 11450
rect 6734 11398 9384 11450
rect 644 11376 9384 11398
rect 2774 11296 2780 11348
rect 2832 11296 2838 11348
rect 3053 11339 3111 11345
rect 3053 11305 3065 11339
rect 3099 11336 3111 11339
rect 4614 11336 4620 11348
rect 3099 11308 4620 11336
rect 3099 11305 3111 11308
rect 3053 11299 3111 11305
rect 4614 11296 4620 11308
rect 4672 11296 4678 11348
rect 6825 11339 6883 11345
rect 6825 11305 6837 11339
rect 6871 11336 6883 11339
rect 7190 11336 7196 11348
rect 6871 11308 7196 11336
rect 6871 11305 6883 11308
rect 6825 11299 6883 11305
rect 7190 11296 7196 11308
rect 7248 11296 7254 11348
rect 2317 11271 2375 11277
rect 2317 11237 2329 11271
rect 2363 11268 2375 11271
rect 2406 11268 2412 11280
rect 2363 11240 2412 11268
rect 2363 11237 2375 11240
rect 2317 11231 2375 11237
rect 2406 11228 2412 11240
rect 2464 11228 2470 11280
rect 2792 11268 2820 11296
rect 2792 11240 3648 11268
rect 1394 11160 1400 11212
rect 1452 11200 1458 11212
rect 2777 11203 2835 11209
rect 1452 11172 2728 11200
rect 1452 11160 1458 11172
rect 2130 11092 2136 11144
rect 2188 11092 2194 11144
rect 2222 11092 2228 11144
rect 2280 11132 2286 11144
rect 2700 11141 2728 11172
rect 2777 11169 2789 11203
rect 2823 11200 2835 11203
rect 3513 11203 3571 11209
rect 3513 11200 3525 11203
rect 2823 11172 3525 11200
rect 2823 11169 2835 11172
rect 2777 11163 2835 11169
rect 3513 11169 3525 11172
rect 3559 11169 3571 11203
rect 3620 11200 3648 11240
rect 3881 11203 3939 11209
rect 3881 11200 3893 11203
rect 3620 11172 3893 11200
rect 3513 11163 3571 11169
rect 3881 11169 3893 11172
rect 3927 11200 3939 11203
rect 4062 11200 4068 11212
rect 3927 11172 4068 11200
rect 3927 11169 3939 11172
rect 3881 11163 3939 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 8754 11200 8760 11212
rect 5828 11172 8760 11200
rect 2409 11135 2467 11141
rect 2409 11132 2421 11135
rect 2280 11104 2421 11132
rect 2280 11092 2286 11104
rect 2409 11101 2421 11104
rect 2455 11101 2467 11135
rect 2409 11095 2467 11101
rect 2685 11135 2743 11141
rect 2685 11101 2697 11135
rect 2731 11132 2743 11135
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2731 11104 2973 11132
rect 2731 11101 2743 11104
rect 2685 11095 2743 11101
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 5350 11092 5356 11144
rect 5408 11092 5414 11144
rect 1026 11024 1032 11076
rect 1084 11024 1090 11076
rect 1670 11024 1676 11076
rect 1728 11064 1734 11076
rect 1857 11067 1915 11073
rect 1857 11064 1869 11067
rect 1728 11036 1869 11064
rect 1728 11024 1734 11036
rect 1857 11033 1869 11036
rect 1903 11033 1915 11067
rect 5166 11064 5172 11076
rect 1857 11027 1915 11033
rect 2746 11036 3556 11064
rect 5014 11036 5172 11064
rect 2593 10999 2651 11005
rect 2593 10965 2605 10999
rect 2639 10996 2651 10999
rect 2746 10996 2774 11036
rect 2639 10968 2774 10996
rect 3528 10996 3556 11036
rect 5166 11024 5172 11036
rect 5224 11024 5230 11076
rect 5828 11064 5856 11172
rect 8754 11160 8760 11172
rect 8812 11200 8818 11212
rect 8812 11172 8892 11200
rect 8812 11160 8818 11172
rect 6270 11092 6276 11144
rect 6328 11092 6334 11144
rect 8864 11141 8892 11172
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11101 6975 11135
rect 6917 11095 6975 11101
rect 8849 11135 8907 11141
rect 8849 11101 8861 11135
rect 8895 11101 8907 11135
rect 8849 11095 8907 11101
rect 5276 11036 5856 11064
rect 5917 11067 5975 11073
rect 5276 10996 5304 11036
rect 5917 11033 5929 11067
rect 5963 11064 5975 11067
rect 6932 11064 6960 11095
rect 5963 11036 6960 11064
rect 5963 11033 5975 11036
rect 5917 11027 5975 11033
rect 8110 11024 8116 11076
rect 8168 11024 8174 11076
rect 8665 11067 8723 11073
rect 8665 11033 8677 11067
rect 8711 11064 8723 11067
rect 9122 11064 9128 11076
rect 8711 11036 9128 11064
rect 8711 11033 8723 11036
rect 8665 11027 8723 11033
rect 9122 11024 9128 11036
rect 9180 11024 9186 11076
rect 3528 10968 5304 10996
rect 2639 10965 2651 10968
rect 2593 10959 2651 10965
rect 8478 10956 8484 11008
rect 8536 10956 8542 11008
rect 644 10906 9384 10928
rect 644 10854 2954 10906
rect 3006 10854 3018 10906
rect 3070 10854 3082 10906
rect 3134 10854 6954 10906
rect 7006 10854 7018 10906
rect 7070 10854 7082 10906
rect 7134 10854 9384 10906
rect 644 10832 9384 10854
rect 4062 10752 4068 10804
rect 4120 10792 4126 10804
rect 4525 10795 4583 10801
rect 4525 10792 4537 10795
rect 4120 10764 4537 10792
rect 4120 10752 4126 10764
rect 4525 10761 4537 10764
rect 4571 10761 4583 10795
rect 4525 10755 4583 10761
rect 5261 10795 5319 10801
rect 5261 10761 5273 10795
rect 5307 10792 5319 10795
rect 5350 10792 5356 10804
rect 5307 10764 5356 10792
rect 5307 10761 5319 10764
rect 5261 10755 5319 10761
rect 5350 10752 5356 10764
rect 5408 10752 5414 10804
rect 6457 10795 6515 10801
rect 6457 10761 6469 10795
rect 6503 10792 6515 10795
rect 8294 10792 8300 10804
rect 6503 10764 8300 10792
rect 6503 10761 6515 10764
rect 6457 10755 6515 10761
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 474 10684 480 10736
rect 532 10724 538 10736
rect 1029 10727 1087 10733
rect 1029 10724 1041 10727
rect 532 10696 1041 10724
rect 532 10684 538 10696
rect 1029 10693 1041 10696
rect 1075 10693 1087 10727
rect 1029 10687 1087 10693
rect 1394 10684 1400 10736
rect 1452 10724 1458 10736
rect 1762 10724 1768 10736
rect 1452 10696 1768 10724
rect 1452 10684 1458 10696
rect 1762 10684 1768 10696
rect 1820 10724 1826 10736
rect 1857 10727 1915 10733
rect 1857 10724 1869 10727
rect 1820 10696 1869 10724
rect 1820 10684 1826 10696
rect 1857 10693 1869 10696
rect 1903 10693 1915 10727
rect 1857 10687 1915 10693
rect 5626 10684 5632 10736
rect 5684 10684 5690 10736
rect 5994 10684 6000 10736
rect 6052 10724 6058 10736
rect 6089 10727 6147 10733
rect 6089 10724 6101 10727
rect 6052 10696 6101 10724
rect 6052 10684 6058 10696
rect 6089 10693 6101 10696
rect 6135 10693 6147 10727
rect 8202 10724 8208 10736
rect 8050 10696 8208 10724
rect 6089 10687 6147 10693
rect 8202 10684 8208 10696
rect 8260 10684 8266 10736
rect 4154 10656 4160 10668
rect 3358 10642 4160 10656
rect 3344 10628 4160 10642
rect 1670 10548 1676 10600
rect 1728 10588 1734 10600
rect 1949 10591 2007 10597
rect 1949 10588 1961 10591
rect 1728 10560 1961 10588
rect 1728 10548 1734 10560
rect 1949 10557 1961 10560
rect 1995 10557 2007 10591
rect 1949 10551 2007 10557
rect 2222 10548 2228 10600
rect 2280 10548 2286 10600
rect 2038 10412 2044 10464
rect 2096 10452 2102 10464
rect 3344 10452 3372 10628
rect 4154 10616 4160 10628
rect 4212 10656 4218 10668
rect 4522 10656 4528 10668
rect 4212 10628 4528 10656
rect 4212 10616 4218 10628
rect 4522 10616 4528 10628
rect 4580 10616 4586 10668
rect 5350 10616 5356 10668
rect 5408 10656 5414 10668
rect 5445 10659 5503 10665
rect 5445 10656 5457 10659
rect 5408 10628 5457 10656
rect 5408 10616 5414 10628
rect 5445 10625 5457 10628
rect 5491 10625 5503 10659
rect 5445 10619 5503 10625
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 6178 10656 6184 10668
rect 5592 10628 6184 10656
rect 5592 10616 5598 10628
rect 6178 10616 6184 10628
rect 6236 10656 6242 10668
rect 6273 10659 6331 10665
rect 6273 10656 6285 10659
rect 6236 10628 6285 10656
rect 6236 10616 6242 10628
rect 6273 10625 6285 10628
rect 6319 10625 6331 10659
rect 6273 10619 6331 10625
rect 8389 10659 8447 10665
rect 8389 10625 8401 10659
rect 8435 10656 8447 10659
rect 8478 10656 8484 10668
rect 8435 10628 8484 10656
rect 8435 10625 8447 10628
rect 8389 10619 8447 10625
rect 8478 10616 8484 10628
rect 8536 10616 8542 10668
rect 3602 10548 3608 10600
rect 3660 10588 3666 10600
rect 3789 10591 3847 10597
rect 3789 10588 3801 10591
rect 3660 10560 3801 10588
rect 3660 10548 3666 10560
rect 3789 10557 3801 10560
rect 3835 10557 3847 10591
rect 5077 10591 5135 10597
rect 5077 10588 5089 10591
rect 3789 10551 3847 10557
rect 4126 10560 5089 10588
rect 3697 10523 3755 10529
rect 3697 10489 3709 10523
rect 3743 10520 3755 10523
rect 4126 10520 4154 10560
rect 5077 10557 5089 10560
rect 5123 10557 5135 10591
rect 5077 10551 5135 10557
rect 5718 10548 5724 10600
rect 5776 10588 5782 10600
rect 6549 10591 6607 10597
rect 6549 10588 6561 10591
rect 5776 10560 6561 10588
rect 5776 10548 5782 10560
rect 6549 10557 6561 10560
rect 6595 10557 6607 10591
rect 6917 10591 6975 10597
rect 6917 10588 6929 10591
rect 6549 10551 6607 10557
rect 6656 10560 6929 10588
rect 3743 10492 4154 10520
rect 3743 10489 3755 10492
rect 3697 10483 3755 10489
rect 6178 10480 6184 10532
rect 6236 10520 6242 10532
rect 6656 10520 6684 10560
rect 6917 10557 6929 10560
rect 6963 10557 6975 10591
rect 6917 10551 6975 10557
rect 8662 10520 8668 10532
rect 6236 10492 6684 10520
rect 7852 10492 8668 10520
rect 6236 10480 6242 10492
rect 2096 10424 3372 10452
rect 2096 10412 2102 10424
rect 4338 10412 4344 10464
rect 4396 10452 4402 10464
rect 4433 10455 4491 10461
rect 4433 10452 4445 10455
rect 4396 10424 4445 10452
rect 4396 10412 4402 10424
rect 4433 10421 4445 10424
rect 4479 10421 4491 10455
rect 4433 10415 4491 10421
rect 4982 10412 4988 10464
rect 5040 10452 5046 10464
rect 7852 10452 7880 10492
rect 8662 10480 8668 10492
rect 8720 10480 8726 10532
rect 5040 10424 7880 10452
rect 5040 10412 5046 10424
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 8949 10455 9007 10461
rect 8949 10452 8961 10455
rect 8352 10424 8961 10452
rect 8352 10412 8358 10424
rect 8949 10421 8961 10424
rect 8995 10421 9007 10455
rect 8949 10415 9007 10421
rect 644 10362 9384 10384
rect 644 10310 2554 10362
rect 2606 10310 2618 10362
rect 2670 10310 2682 10362
rect 2734 10310 6554 10362
rect 6606 10310 6618 10362
rect 6670 10310 6682 10362
rect 6734 10310 9384 10362
rect 644 10288 9384 10310
rect 2038 10208 2044 10260
rect 2096 10208 2102 10260
rect 2222 10208 2228 10260
rect 2280 10248 2286 10260
rect 2501 10251 2559 10257
rect 2501 10248 2513 10251
rect 2280 10220 2513 10248
rect 2280 10208 2286 10220
rect 2501 10217 2513 10220
rect 2547 10217 2559 10251
rect 2501 10211 2559 10217
rect 3329 10251 3387 10257
rect 3329 10217 3341 10251
rect 3375 10248 3387 10251
rect 3602 10248 3608 10260
rect 3375 10220 3608 10248
rect 3375 10217 3387 10220
rect 3329 10211 3387 10217
rect 3602 10208 3608 10220
rect 3660 10208 3666 10260
rect 5718 10208 5724 10260
rect 5776 10208 5782 10260
rect 5166 10140 5172 10192
rect 5224 10140 5230 10192
rect 5626 10180 5632 10192
rect 5460 10152 5632 10180
rect 474 10072 480 10124
rect 532 10112 538 10124
rect 1029 10115 1087 10121
rect 1029 10112 1041 10115
rect 532 10084 1041 10112
rect 532 10072 538 10084
rect 1029 10081 1041 10084
rect 1075 10081 1087 10115
rect 1029 10075 1087 10081
rect 2222 10004 2228 10056
rect 2280 10004 2286 10056
rect 2774 10004 2780 10056
rect 2832 10044 2838 10056
rect 3053 10047 3111 10053
rect 3053 10044 3065 10047
rect 2832 10016 3065 10044
rect 2832 10004 2838 10016
rect 3053 10013 3065 10016
rect 3099 10013 3111 10047
rect 3053 10007 3111 10013
rect 5074 10004 5080 10056
rect 5132 10004 5138 10056
rect 5460 10053 5488 10152
rect 5626 10140 5632 10152
rect 5684 10140 5690 10192
rect 5902 10140 5908 10192
rect 5960 10180 5966 10192
rect 7650 10180 7656 10192
rect 5960 10152 7656 10180
rect 5960 10140 5966 10152
rect 7650 10140 7656 10152
rect 7708 10140 7714 10192
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8481 10183 8539 10189
rect 8481 10180 8493 10183
rect 8260 10152 8493 10180
rect 8260 10140 8266 10152
rect 8481 10149 8493 10152
rect 8527 10149 8539 10183
rect 8481 10143 8539 10149
rect 7837 10115 7895 10121
rect 5644 10084 6868 10112
rect 5644 10056 5672 10084
rect 5444 10047 5502 10053
rect 5444 10013 5456 10047
rect 5490 10013 5502 10047
rect 5444 10007 5502 10013
rect 5534 10004 5540 10056
rect 5592 10004 5598 10056
rect 5626 10004 5632 10056
rect 5684 10004 5690 10056
rect 5905 10047 5963 10053
rect 5905 10013 5917 10047
rect 5951 10013 5963 10047
rect 5905 10007 5963 10013
rect 1857 9979 1915 9985
rect 1857 9945 1869 9979
rect 1903 9976 1915 9979
rect 1946 9976 1952 9988
rect 1903 9948 1952 9976
rect 1903 9945 1915 9948
rect 1857 9939 1915 9945
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 4154 9936 4160 9988
rect 4212 9936 4218 9988
rect 4801 9979 4859 9985
rect 4801 9945 4813 9979
rect 4847 9945 4859 9979
rect 4801 9939 4859 9945
rect 4816 9908 4844 9939
rect 5166 9936 5172 9988
rect 5224 9976 5230 9988
rect 5920 9976 5948 10007
rect 5994 10004 6000 10056
rect 6052 10044 6058 10056
rect 6454 10044 6460 10056
rect 6052 10016 6460 10044
rect 6052 10004 6058 10016
rect 6454 10004 6460 10016
rect 6512 10004 6518 10056
rect 6840 10053 6868 10084
rect 7837 10081 7849 10115
rect 7883 10112 7895 10115
rect 9582 10112 9588 10124
rect 7883 10084 9588 10112
rect 7883 10081 7895 10084
rect 7837 10075 7895 10081
rect 9582 10072 9588 10084
rect 9640 10072 9646 10124
rect 6825 10047 6883 10053
rect 6825 10013 6837 10047
rect 6871 10044 6883 10047
rect 8018 10044 8024 10056
rect 6871 10016 8024 10044
rect 6871 10013 6883 10016
rect 6825 10007 6883 10013
rect 8018 10004 8024 10016
rect 8076 10004 8082 10056
rect 8294 10004 8300 10056
rect 8352 10004 8358 10056
rect 8754 10004 8760 10056
rect 8812 10004 8818 10056
rect 8849 10047 8907 10053
rect 8849 10013 8861 10047
rect 8895 10044 8907 10047
rect 9122 10044 9128 10056
rect 8895 10016 9128 10044
rect 8895 10013 8907 10016
rect 8849 10007 8907 10013
rect 9122 10004 9128 10016
rect 9180 10004 9186 10056
rect 5224 9948 5948 9976
rect 5224 9936 5230 9948
rect 6362 9936 6368 9988
rect 6420 9976 6426 9988
rect 6733 9979 6791 9985
rect 6733 9976 6745 9979
rect 6420 9948 6745 9976
rect 6420 9936 6426 9948
rect 6733 9945 6745 9948
rect 6779 9945 6791 9979
rect 6733 9939 6791 9945
rect 6454 9908 6460 9920
rect 4816 9880 6460 9908
rect 6454 9868 6460 9880
rect 6512 9908 6518 9920
rect 6549 9911 6607 9917
rect 6549 9908 6561 9911
rect 6512 9880 6561 9908
rect 6512 9868 6518 9880
rect 6549 9877 6561 9880
rect 6595 9877 6607 9911
rect 6549 9871 6607 9877
rect 644 9818 9384 9840
rect 644 9766 2954 9818
rect 3006 9766 3018 9818
rect 3070 9766 3082 9818
rect 3134 9766 6954 9818
rect 7006 9766 7018 9818
rect 7070 9766 7082 9818
rect 7134 9766 9384 9818
rect 644 9744 9384 9766
rect 1670 9664 1676 9716
rect 1728 9704 1734 9716
rect 1728 9676 3464 9704
rect 1728 9664 1734 9676
rect 1688 9636 1716 9664
rect 1044 9608 1716 9636
rect 1044 9577 1072 9608
rect 2038 9596 2044 9648
rect 2096 9596 2102 9648
rect 3436 9636 3464 9676
rect 3602 9664 3608 9716
rect 3660 9704 3666 9716
rect 4154 9704 4160 9716
rect 3660 9676 4160 9704
rect 3660 9664 3666 9676
rect 4154 9664 4160 9676
rect 4212 9704 4218 9716
rect 5721 9707 5779 9713
rect 4212 9676 5580 9704
rect 4212 9664 4218 9676
rect 5552 9648 5580 9676
rect 5721 9673 5733 9707
rect 5767 9704 5779 9707
rect 6270 9704 6276 9716
rect 5767 9676 6276 9704
rect 5767 9673 5779 9676
rect 5721 9667 5779 9673
rect 6270 9664 6276 9676
rect 6328 9664 6334 9716
rect 9122 9704 9128 9716
rect 6380 9676 9128 9704
rect 4249 9639 4307 9645
rect 3436 9608 4016 9636
rect 1029 9571 1087 9577
rect 1029 9537 1041 9571
rect 1075 9537 1087 9571
rect 1029 9531 1087 9537
rect 2961 9571 3019 9577
rect 2961 9537 2973 9571
rect 3007 9568 3019 9571
rect 3234 9568 3240 9580
rect 3007 9540 3240 9568
rect 3007 9537 3019 9540
rect 2961 9531 3019 9537
rect 3234 9528 3240 9540
rect 3292 9528 3298 9580
rect 3436 9577 3464 9608
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3513 9571 3571 9577
rect 3513 9537 3525 9571
rect 3559 9537 3571 9571
rect 3513 9531 3571 9537
rect 1305 9503 1363 9509
rect 1305 9469 1317 9503
rect 1351 9500 1363 9503
rect 1670 9500 1676 9512
rect 1351 9472 1676 9500
rect 1351 9469 1363 9472
rect 1305 9463 1363 9469
rect 1670 9460 1676 9472
rect 1728 9460 1734 9512
rect 2314 9460 2320 9512
rect 2372 9500 2378 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 2372 9472 3341 9500
rect 2372 9460 2378 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 2774 9392 2780 9444
rect 2832 9392 2838 9444
rect 3528 9432 3556 9531
rect 3988 9512 4016 9608
rect 4249 9605 4261 9639
rect 4295 9636 4307 9639
rect 4338 9636 4344 9648
rect 4295 9608 4344 9636
rect 4295 9605 4307 9608
rect 4249 9599 4307 9605
rect 4338 9596 4344 9608
rect 4396 9596 4402 9648
rect 5534 9596 5540 9648
rect 5592 9636 5598 9648
rect 5997 9639 6055 9645
rect 5997 9636 6009 9639
rect 5592 9608 6009 9636
rect 5592 9596 5598 9608
rect 5997 9605 6009 9608
rect 6043 9605 6055 9639
rect 5997 9599 6055 9605
rect 6181 9639 6239 9645
rect 6181 9605 6193 9639
rect 6227 9636 6239 9639
rect 6380 9636 6408 9676
rect 9122 9664 9128 9676
rect 9180 9664 9186 9716
rect 8478 9636 8484 9648
rect 6227 9608 6408 9636
rect 7866 9608 8484 9636
rect 6227 9605 6239 9608
rect 6181 9599 6239 9605
rect 5350 9528 5356 9580
rect 5408 9568 5414 9580
rect 6196 9568 6224 9599
rect 8478 9596 8484 9608
rect 8536 9596 8542 9648
rect 5408 9540 6224 9568
rect 5408 9528 5414 9540
rect 6362 9528 6368 9580
rect 6420 9528 6426 9580
rect 8202 9528 8208 9580
rect 8260 9528 8266 9580
rect 3970 9460 3976 9512
rect 4028 9460 4034 9512
rect 4614 9500 4620 9512
rect 4080 9472 4620 9500
rect 4080 9432 4108 9472
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 6454 9460 6460 9512
rect 6512 9500 6518 9512
rect 6733 9503 6791 9509
rect 6733 9500 6745 9503
rect 6512 9472 6745 9500
rect 6512 9460 6518 9472
rect 6733 9469 6745 9472
rect 6779 9469 6791 9503
rect 6733 9463 6791 9469
rect 3068 9404 3556 9432
rect 3620 9404 4108 9432
rect 1854 9324 1860 9376
rect 1912 9364 1918 9376
rect 3068 9364 3096 9404
rect 1912 9336 3096 9364
rect 3145 9367 3203 9373
rect 1912 9324 1918 9336
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3620 9364 3648 9404
rect 3191 9336 3648 9364
rect 3697 9367 3755 9373
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3697 9333 3709 9367
rect 3743 9364 3755 9367
rect 4246 9364 4252 9376
rect 3743 9336 4252 9364
rect 3743 9333 3755 9336
rect 3697 9327 3755 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4890 9324 4896 9376
rect 4948 9364 4954 9376
rect 7190 9364 7196 9376
rect 4948 9336 7196 9364
rect 4948 9324 4954 9336
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 8110 9324 8116 9376
rect 8168 9364 8174 9376
rect 8765 9367 8823 9373
rect 8765 9364 8777 9367
rect 8168 9336 8777 9364
rect 8168 9324 8174 9336
rect 8765 9333 8777 9336
rect 8811 9333 8823 9367
rect 8765 9327 8823 9333
rect 644 9274 9384 9296
rect 644 9222 2554 9274
rect 2606 9222 2618 9274
rect 2670 9222 2682 9274
rect 2734 9222 6554 9274
rect 6606 9222 6618 9274
rect 6670 9222 6682 9274
rect 6734 9222 9384 9274
rect 644 9200 9384 9222
rect 2130 9120 2136 9172
rect 2188 9160 2194 9172
rect 6362 9160 6368 9172
rect 2188 9132 6368 9160
rect 2188 9120 2194 9132
rect 6362 9120 6368 9132
rect 6420 9120 6426 9172
rect 6454 9120 6460 9172
rect 6512 9160 6518 9172
rect 6512 9132 6776 9160
rect 6512 9120 6518 9132
rect 2038 9052 2044 9104
rect 2096 9092 2102 9104
rect 2096 9064 2544 9092
rect 2096 9052 2102 9064
rect 2516 9024 2544 9064
rect 2774 9052 2780 9104
rect 2832 9092 2838 9104
rect 2961 9095 3019 9101
rect 2961 9092 2973 9095
rect 2832 9064 2973 9092
rect 2832 9052 2838 9064
rect 2961 9061 2973 9064
rect 3007 9061 3019 9095
rect 4062 9092 4068 9104
rect 2961 9055 3019 9061
rect 3344 9064 4068 9092
rect 2516 8996 2912 9024
rect 2130 8916 2136 8968
rect 2188 8916 2194 8968
rect 2884 8965 2912 8996
rect 2715 8959 2773 8965
rect 2715 8925 2727 8959
rect 2761 8925 2773 8959
rect 2715 8919 2773 8925
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8925 2927 8959
rect 2869 8919 2927 8925
rect 3145 8959 3203 8965
rect 3145 8925 3157 8959
rect 3191 8956 3203 8959
rect 3234 8956 3240 8968
rect 3191 8928 3240 8956
rect 3191 8925 3203 8928
rect 3145 8919 3203 8925
rect 382 8848 388 8900
rect 440 8888 446 8900
rect 1121 8891 1179 8897
rect 1121 8888 1133 8891
rect 440 8860 1133 8888
rect 440 8848 446 8860
rect 1121 8857 1133 8860
rect 1167 8857 1179 8891
rect 1121 8851 1179 8857
rect 1210 8848 1216 8900
rect 1268 8888 1274 8900
rect 2038 8888 2044 8900
rect 1268 8860 2044 8888
rect 1268 8848 1274 8860
rect 2038 8848 2044 8860
rect 2096 8888 2102 8900
rect 2730 8888 2758 8919
rect 3234 8916 3240 8928
rect 3292 8916 3298 8968
rect 3344 8965 3372 9064
rect 4062 9052 4068 9064
rect 4120 9052 4126 9104
rect 4985 9095 5043 9101
rect 4985 9061 4997 9095
rect 5031 9092 5043 9095
rect 5166 9092 5172 9104
rect 5031 9064 5172 9092
rect 5031 9061 5043 9064
rect 4985 9055 5043 9061
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 6748 9092 6776 9132
rect 6822 9120 6828 9172
rect 6880 9160 6886 9172
rect 7377 9163 7435 9169
rect 7377 9160 7389 9163
rect 6880 9132 7389 9160
rect 6880 9120 6886 9132
rect 7377 9129 7389 9132
rect 7423 9129 7435 9163
rect 7377 9123 7435 9129
rect 6748 9064 6868 9092
rect 3970 8984 3976 9036
rect 4028 9024 4034 9036
rect 4890 9024 4896 9036
rect 4028 8996 4896 9024
rect 4028 8984 4034 8996
rect 4890 8984 4896 8996
rect 4948 9024 4954 9036
rect 5074 9024 5080 9036
rect 4948 8996 5080 9024
rect 4948 8984 4954 8996
rect 5074 8984 5080 8996
rect 5132 9024 5138 9036
rect 6733 9027 6791 9033
rect 6733 9024 6745 9027
rect 5132 8996 6745 9024
rect 5132 8984 5138 8996
rect 6733 8993 6745 8996
rect 6779 8993 6791 9027
rect 6733 8987 6791 8993
rect 3329 8959 3387 8965
rect 3329 8925 3341 8959
rect 3375 8925 3387 8959
rect 3329 8919 3387 8925
rect 3605 8959 3663 8965
rect 3605 8925 3617 8959
rect 3651 8956 3663 8959
rect 4982 8956 4988 8968
rect 3651 8928 4988 8956
rect 3651 8925 3663 8928
rect 3605 8919 3663 8925
rect 4982 8916 4988 8928
rect 5040 8916 5046 8968
rect 5350 8916 5356 8968
rect 5408 8916 5414 8968
rect 6840 8965 6868 9064
rect 8478 9052 8484 9104
rect 8536 9052 8542 9104
rect 8018 9024 8024 9036
rect 7484 8996 8024 9024
rect 6825 8959 6883 8965
rect 6825 8925 6837 8959
rect 6871 8925 6883 8959
rect 6825 8919 6883 8925
rect 6979 8959 7037 8965
rect 6979 8925 6991 8959
rect 7025 8956 7037 8959
rect 7190 8956 7196 8968
rect 7025 8928 7196 8956
rect 7025 8925 7037 8928
rect 6979 8919 7037 8925
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 7484 8965 7512 8996
rect 8018 8984 8024 8996
rect 8076 8984 8082 9036
rect 7469 8959 7527 8965
rect 7469 8925 7481 8959
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7650 8916 7656 8968
rect 7708 8916 7714 8968
rect 8754 8965 8760 8968
rect 8725 8959 8760 8965
rect 8725 8958 8737 8959
rect 8588 8930 8737 8958
rect 5166 8888 5172 8900
rect 2096 8860 2758 8888
rect 3528 8860 5172 8888
rect 2096 8848 2102 8860
rect 2406 8780 2412 8832
rect 2464 8820 2470 8832
rect 3528 8829 3556 8860
rect 5166 8848 5172 8860
rect 5224 8848 5230 8900
rect 6178 8848 6184 8900
rect 6236 8888 6242 8900
rect 6457 8891 6515 8897
rect 6457 8888 6469 8891
rect 6236 8860 6469 8888
rect 6236 8848 6242 8860
rect 6457 8857 6469 8860
rect 6503 8857 6515 8891
rect 8588 8888 8616 8930
rect 8725 8925 8737 8930
rect 8725 8919 8760 8925
rect 8754 8916 8760 8919
rect 8812 8916 8818 8968
rect 8849 8959 8907 8965
rect 8849 8925 8861 8959
rect 8895 8956 8907 8959
rect 9122 8956 9128 8968
rect 8895 8928 9128 8956
rect 8895 8925 8907 8928
rect 8849 8919 8907 8925
rect 9122 8916 9128 8928
rect 9180 8916 9186 8968
rect 6457 8851 6515 8857
rect 6748 8860 8616 8888
rect 2501 8823 2559 8829
rect 2501 8820 2513 8823
rect 2464 8792 2513 8820
rect 2464 8780 2470 8792
rect 2501 8789 2513 8792
rect 2547 8789 2559 8823
rect 2501 8783 2559 8789
rect 3513 8823 3571 8829
rect 3513 8789 3525 8823
rect 3559 8789 3571 8823
rect 3513 8783 3571 8789
rect 3789 8823 3847 8829
rect 3789 8789 3801 8823
rect 3835 8820 3847 8823
rect 6748 8820 6776 8860
rect 3835 8792 6776 8820
rect 3835 8789 3847 8792
rect 3789 8783 3847 8789
rect 6822 8780 6828 8832
rect 6880 8820 6886 8832
rect 7193 8823 7251 8829
rect 7193 8820 7205 8823
rect 6880 8792 7205 8820
rect 6880 8780 6886 8792
rect 7193 8789 7205 8792
rect 7239 8789 7251 8823
rect 7193 8783 7251 8789
rect 8110 8780 8116 8832
rect 8168 8820 8174 8832
rect 8205 8823 8263 8829
rect 8205 8820 8217 8823
rect 8168 8792 8217 8820
rect 8168 8780 8174 8792
rect 8205 8789 8217 8792
rect 8251 8789 8263 8823
rect 8205 8783 8263 8789
rect 644 8730 9384 8752
rect 644 8678 2954 8730
rect 3006 8678 3018 8730
rect 3070 8678 3082 8730
rect 3134 8678 6954 8730
rect 7006 8678 7018 8730
rect 7070 8678 7082 8730
rect 7134 8678 9384 8730
rect 644 8656 9384 8678
rect 1762 8616 1768 8628
rect 1044 8588 1768 8616
rect 1044 8492 1072 8588
rect 1762 8576 1768 8588
rect 1820 8616 1826 8628
rect 5074 8616 5080 8628
rect 1820 8588 5080 8616
rect 1820 8576 1826 8588
rect 5074 8576 5080 8588
rect 5132 8616 5138 8628
rect 5626 8616 5632 8628
rect 5132 8588 5632 8616
rect 5132 8576 5138 8588
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5718 8576 5724 8628
rect 5776 8616 5782 8628
rect 6454 8616 6460 8628
rect 5776 8588 6460 8616
rect 5776 8576 5782 8588
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 2406 8508 2412 8560
rect 2464 8508 2470 8560
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3881 8551 3939 8557
rect 3881 8548 3893 8551
rect 3292 8520 3893 8548
rect 3292 8508 3298 8520
rect 3881 8517 3893 8520
rect 3927 8517 3939 8551
rect 3881 8511 3939 8517
rect 5902 8508 5908 8560
rect 5960 8548 5966 8560
rect 7650 8548 7656 8560
rect 5960 8520 7656 8548
rect 5960 8508 5966 8520
rect 7650 8508 7656 8520
rect 7708 8508 7714 8560
rect 1026 8440 1032 8492
rect 1084 8440 1090 8492
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 3145 8483 3203 8489
rect 3145 8449 3157 8483
rect 3191 8449 3203 8483
rect 3145 8443 3203 8449
rect 1121 8415 1179 8421
rect 1121 8381 1133 8415
rect 1167 8412 1179 8415
rect 1305 8415 1363 8421
rect 1305 8412 1317 8415
rect 1167 8384 1317 8412
rect 1167 8381 1179 8384
rect 1121 8375 1179 8381
rect 1305 8381 1317 8384
rect 1351 8381 1363 8415
rect 3160 8412 3188 8443
rect 3602 8440 3608 8492
rect 3660 8480 3666 8492
rect 4065 8483 4123 8489
rect 4065 8480 4077 8483
rect 3660 8452 4077 8480
rect 3660 8440 3666 8452
rect 4065 8449 4077 8452
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 6362 8440 6368 8492
rect 6420 8440 6426 8492
rect 7190 8440 7196 8492
rect 7248 8480 7254 8492
rect 8662 8480 8668 8492
rect 7248 8452 8668 8480
rect 7248 8440 7254 8452
rect 8662 8440 8668 8452
rect 8720 8440 8726 8492
rect 8938 8440 8944 8492
rect 8996 8440 9002 8492
rect 4249 8415 4307 8421
rect 4249 8412 4261 8415
rect 3160 8384 4261 8412
rect 1305 8375 1363 8381
rect 4249 8381 4261 8384
rect 4295 8381 4307 8415
rect 4249 8375 4307 8381
rect 6454 8372 6460 8424
rect 6512 8412 6518 8424
rect 6733 8415 6791 8421
rect 6733 8412 6745 8415
rect 6512 8384 6745 8412
rect 6512 8372 6518 8384
rect 6733 8381 6745 8384
rect 6779 8381 6791 8415
rect 6733 8375 6791 8381
rect 8573 8415 8631 8421
rect 8573 8381 8585 8415
rect 8619 8412 8631 8415
rect 9582 8412 9588 8424
rect 8619 8384 9588 8412
rect 8619 8381 8631 8384
rect 8573 8375 8631 8381
rect 9582 8372 9588 8384
rect 9640 8372 9646 8424
rect 4338 8304 4344 8356
rect 4396 8344 4402 8356
rect 6181 8347 6239 8353
rect 6181 8344 6193 8347
rect 4396 8316 6193 8344
rect 4396 8304 4402 8316
rect 6181 8313 6193 8316
rect 6227 8313 6239 8347
rect 6181 8307 6239 8313
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 2222 8276 2228 8288
rect 2096 8248 2228 8276
rect 2096 8236 2102 8248
rect 2222 8236 2228 8248
rect 2280 8236 2286 8288
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 3705 8279 3763 8285
rect 3705 8276 3717 8279
rect 3660 8248 3717 8276
rect 3660 8236 3666 8248
rect 3705 8245 3717 8248
rect 3751 8245 3763 8279
rect 3705 8239 3763 8245
rect 6641 8279 6699 8285
rect 6641 8245 6653 8279
rect 6687 8276 6699 8279
rect 7190 8276 7196 8288
rect 6687 8248 7196 8276
rect 6687 8245 6699 8248
rect 6641 8239 6699 8245
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7377 8279 7435 8285
rect 7377 8245 7389 8279
rect 7423 8276 7435 8279
rect 7650 8276 7656 8288
rect 7423 8248 7656 8276
rect 7423 8245 7435 8248
rect 7377 8239 7435 8245
rect 7650 8236 7656 8248
rect 7708 8236 7714 8288
rect 644 8186 9384 8208
rect 644 8134 2554 8186
rect 2606 8134 2618 8186
rect 2670 8134 2682 8186
rect 2734 8134 6554 8186
rect 6606 8134 6618 8186
rect 6670 8134 6682 8186
rect 6734 8134 9384 8186
rect 644 8112 9384 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 4430 8072 4436 8084
rect 1811 8044 4436 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 4430 8032 4436 8044
rect 4488 8032 4494 8084
rect 8202 8032 8208 8084
rect 8260 8072 8266 8084
rect 8481 8075 8539 8081
rect 8481 8072 8493 8075
rect 8260 8044 8493 8072
rect 8260 8032 8266 8044
rect 8481 8041 8493 8044
rect 8527 8041 8539 8075
rect 8481 8035 8539 8041
rect 2593 8007 2651 8013
rect 2593 7973 2605 8007
rect 2639 8004 2651 8007
rect 5902 8004 5908 8016
rect 2639 7976 5908 8004
rect 2639 7973 2651 7976
rect 2593 7967 2651 7973
rect 5902 7964 5908 7976
rect 5960 7964 5966 8016
rect 1213 7939 1271 7945
rect 1213 7905 1225 7939
rect 1259 7936 1271 7939
rect 2041 7939 2099 7945
rect 2041 7936 2053 7939
rect 1259 7908 2053 7936
rect 1259 7905 1271 7908
rect 1213 7899 1271 7905
rect 2041 7905 2053 7908
rect 2087 7936 2099 7939
rect 3602 7936 3608 7948
rect 2087 7908 3608 7936
rect 2087 7905 2099 7908
rect 2041 7899 2099 7905
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8386 7936 8392 7948
rect 7883 7908 8392 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8386 7896 8392 7908
rect 8444 7896 8450 7948
rect 1397 7871 1455 7877
rect 1397 7837 1409 7871
rect 1443 7868 1455 7871
rect 2774 7868 2780 7880
rect 1443 7840 2780 7868
rect 1443 7837 1455 7840
rect 1397 7831 1455 7837
rect 2774 7828 2780 7840
rect 2832 7828 2838 7880
rect 3234 7828 3240 7880
rect 3292 7868 3298 7880
rect 4065 7871 4123 7877
rect 4065 7868 4077 7871
rect 3292 7840 4077 7868
rect 3292 7828 3298 7840
rect 4065 7837 4077 7840
rect 4111 7837 4123 7871
rect 4065 7831 4123 7837
rect 6086 7828 6092 7880
rect 6144 7828 6150 7880
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 8849 7871 8907 7877
rect 8849 7868 8861 7871
rect 8812 7840 8861 7868
rect 8812 7828 8818 7840
rect 8849 7837 8861 7840
rect 8895 7837 8907 7871
rect 8849 7831 8907 7837
rect 1118 7760 1124 7812
rect 1176 7800 1182 7812
rect 2133 7803 2191 7809
rect 2133 7800 2145 7803
rect 1176 7772 2145 7800
rect 1176 7760 1182 7772
rect 2133 7769 2145 7772
rect 2179 7769 2191 7803
rect 5626 7800 5632 7812
rect 2133 7763 2191 7769
rect 2746 7772 5632 7800
rect 1302 7692 1308 7744
rect 1360 7692 1366 7744
rect 2222 7692 2228 7744
rect 2280 7692 2286 7744
rect 2314 7692 2320 7744
rect 2372 7732 2378 7744
rect 2746 7732 2774 7772
rect 5626 7760 5632 7772
rect 5684 7760 5690 7812
rect 5718 7760 5724 7812
rect 5776 7800 5782 7812
rect 5813 7803 5871 7809
rect 5813 7800 5825 7803
rect 5776 7772 5825 7800
rect 5776 7760 5782 7772
rect 5813 7769 5825 7772
rect 5859 7769 5871 7803
rect 5813 7763 5871 7769
rect 6270 7760 6276 7812
rect 6328 7800 6334 7812
rect 6733 7803 6791 7809
rect 6733 7800 6745 7803
rect 6328 7772 6745 7800
rect 6328 7760 6334 7772
rect 6733 7769 6745 7772
rect 6779 7769 6791 7803
rect 6733 7763 6791 7769
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 9122 7800 9128 7812
rect 8711 7772 9128 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 9122 7760 9128 7772
rect 9180 7760 9186 7812
rect 2372 7704 2774 7732
rect 4709 7735 4767 7741
rect 2372 7692 2378 7704
rect 4709 7701 4721 7735
rect 4755 7732 4767 7735
rect 4798 7732 4804 7744
rect 4755 7704 4804 7732
rect 4755 7701 4767 7704
rect 4709 7695 4767 7701
rect 4798 7692 4804 7704
rect 4856 7692 4862 7744
rect 5997 7735 6055 7741
rect 5997 7701 6009 7735
rect 6043 7732 6055 7735
rect 6362 7732 6368 7744
rect 6043 7704 6368 7732
rect 6043 7701 6055 7704
rect 5997 7695 6055 7701
rect 6362 7692 6368 7704
rect 6420 7692 6426 7744
rect 644 7642 9384 7664
rect 644 7590 2954 7642
rect 3006 7590 3018 7642
rect 3070 7590 3082 7642
rect 3134 7590 6954 7642
rect 7006 7590 7018 7642
rect 7070 7590 7082 7642
rect 7134 7590 9384 7642
rect 644 7568 9384 7590
rect 1121 7531 1179 7537
rect 1121 7497 1133 7531
rect 1167 7497 1179 7531
rect 1121 7491 1179 7497
rect 1136 7460 1164 7491
rect 1394 7488 1400 7540
rect 1452 7488 1458 7540
rect 3145 7531 3203 7537
rect 3145 7497 3157 7531
rect 3191 7528 3203 7531
rect 3234 7528 3240 7540
rect 3191 7500 3240 7528
rect 3191 7497 3203 7500
rect 3145 7491 3203 7497
rect 3234 7488 3240 7500
rect 3292 7488 3298 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 8489 7531 8547 7537
rect 8489 7528 8501 7531
rect 8352 7500 8501 7528
rect 8352 7488 8358 7500
rect 8489 7497 8501 7500
rect 8535 7497 8547 7531
rect 8489 7491 8547 7497
rect 2222 7460 2228 7472
rect 1136 7432 2228 7460
rect 2222 7420 2228 7432
rect 2280 7420 2286 7472
rect 4617 7463 4675 7469
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 4706 7460 4712 7472
rect 4663 7432 4712 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 4706 7420 4712 7432
rect 4764 7420 4770 7472
rect 6822 7420 6828 7472
rect 6880 7420 6886 7472
rect 8662 7420 8668 7472
rect 8720 7420 8726 7472
rect 934 7352 940 7404
rect 992 7352 998 7404
rect 1210 7352 1216 7404
rect 1268 7352 1274 7404
rect 1670 7284 1676 7336
rect 1728 7324 1734 7336
rect 2225 7327 2283 7333
rect 2225 7324 2237 7327
rect 1728 7296 2237 7324
rect 1728 7284 1734 7296
rect 2225 7293 2237 7296
rect 2271 7293 2283 7327
rect 2225 7287 2283 7293
rect 2406 7284 2412 7336
rect 2464 7324 2470 7336
rect 2777 7327 2835 7333
rect 2777 7324 2789 7327
rect 2464 7296 2789 7324
rect 2464 7284 2470 7296
rect 2777 7293 2789 7296
rect 2823 7293 2835 7327
rect 2777 7287 2835 7293
rect 2038 7216 2044 7268
rect 2096 7256 2102 7268
rect 2314 7256 2320 7268
rect 2096 7228 2320 7256
rect 2096 7216 2102 7228
rect 2314 7216 2320 7228
rect 2372 7256 2378 7268
rect 3528 7256 3556 7378
rect 4890 7352 4896 7404
rect 4948 7352 4954 7404
rect 5074 7352 5080 7404
rect 5132 7352 5138 7404
rect 5626 7392 5632 7404
rect 5587 7364 5632 7392
rect 5626 7352 5632 7364
rect 5684 7352 5690 7404
rect 5718 7352 5724 7404
rect 5776 7352 5782 7404
rect 6270 7352 6276 7404
rect 6328 7392 6334 7404
rect 6457 7395 6515 7401
rect 6457 7392 6469 7395
rect 6328 7364 6469 7392
rect 6328 7352 6334 7364
rect 6457 7361 6469 7364
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 7929 7395 7987 7401
rect 7929 7361 7941 7395
rect 7975 7361 7987 7395
rect 7929 7355 7987 7361
rect 8849 7395 8907 7401
rect 8849 7361 8861 7395
rect 8895 7392 8907 7395
rect 8938 7392 8944 7404
rect 8895 7364 8944 7392
rect 8895 7361 8907 7364
rect 8849 7355 8907 7361
rect 5169 7327 5227 7333
rect 5169 7293 5181 7327
rect 5215 7324 5227 7327
rect 6089 7327 6147 7333
rect 6089 7324 6101 7327
rect 5215 7296 6101 7324
rect 5215 7293 5227 7296
rect 5169 7287 5227 7293
rect 6089 7293 6101 7296
rect 6135 7293 6147 7327
rect 7944 7324 7972 7355
rect 8938 7352 8944 7364
rect 8996 7352 9002 7404
rect 9033 7327 9091 7333
rect 9033 7324 9045 7327
rect 7944 7296 9045 7324
rect 6089 7287 6147 7293
rect 9033 7293 9045 7296
rect 9079 7293 9091 7327
rect 9033 7287 9091 7293
rect 2372 7228 3556 7256
rect 2372 7216 2378 7228
rect 3528 7188 3556 7228
rect 5442 7216 5448 7268
rect 5500 7256 5506 7268
rect 5902 7256 5908 7268
rect 5500 7228 5908 7256
rect 5500 7216 5506 7228
rect 5902 7216 5908 7228
rect 5960 7216 5966 7268
rect 5460 7188 5488 7216
rect 3528 7160 5488 7188
rect 5534 7148 5540 7200
rect 5592 7148 5598 7200
rect 7190 7148 7196 7200
rect 7248 7188 7254 7200
rect 7650 7188 7656 7200
rect 7248 7160 7656 7188
rect 7248 7148 7254 7160
rect 7650 7148 7656 7160
rect 7708 7148 7714 7200
rect 644 7098 9384 7120
rect 644 7046 2554 7098
rect 2606 7046 2618 7098
rect 2670 7046 2682 7098
rect 2734 7046 6554 7098
rect 6606 7046 6618 7098
rect 6670 7046 6682 7098
rect 6734 7046 9384 7098
rect 644 7024 9384 7046
rect 4062 6944 4068 6996
rect 4120 6984 4126 6996
rect 4120 6956 6132 6984
rect 4120 6944 4126 6956
rect 6104 6916 6132 6956
rect 6178 6944 6184 6996
rect 6236 6984 6242 6996
rect 7285 6987 7343 6993
rect 7285 6984 7297 6987
rect 6236 6956 7297 6984
rect 6236 6944 6242 6956
rect 7285 6953 7297 6956
rect 7331 6953 7343 6987
rect 7285 6947 7343 6953
rect 8297 6987 8355 6993
rect 8297 6953 8309 6987
rect 8343 6984 8355 6987
rect 8570 6984 8576 6996
rect 8343 6956 8576 6984
rect 8343 6953 8355 6956
rect 8297 6947 8355 6953
rect 8570 6944 8576 6956
rect 8628 6944 8634 6996
rect 6929 6919 6987 6925
rect 6104 6888 6868 6916
rect 5074 6848 5080 6860
rect 4264 6820 5080 6848
rect 4264 6789 4292 6820
rect 5074 6808 5080 6820
rect 5132 6808 5138 6860
rect 6840 6848 6868 6888
rect 6929 6885 6941 6919
rect 6975 6916 6987 6919
rect 7650 6916 7656 6928
rect 6975 6888 7656 6916
rect 6975 6885 6987 6888
rect 6929 6879 6987 6885
rect 7650 6876 7656 6888
rect 7708 6876 7714 6928
rect 6840 6820 8248 6848
rect 4249 6783 4307 6789
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4525 6783 4583 6789
rect 4525 6780 4537 6783
rect 4387 6752 4537 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4525 6749 4537 6752
rect 4571 6749 4583 6783
rect 4525 6743 4583 6749
rect 4798 6740 4804 6792
rect 4856 6780 4862 6792
rect 4893 6783 4951 6789
rect 4893 6780 4905 6783
rect 4856 6752 4905 6780
rect 4856 6740 4862 6752
rect 4893 6749 4905 6752
rect 4939 6749 4951 6783
rect 4893 6743 4951 6749
rect 6362 6740 6368 6792
rect 6420 6740 6426 6792
rect 7650 6740 7656 6792
rect 7708 6780 7714 6792
rect 7837 6783 7895 6789
rect 7837 6780 7849 6783
rect 7708 6752 7849 6780
rect 7708 6740 7714 6752
rect 7837 6749 7849 6752
rect 7883 6749 7895 6783
rect 7837 6743 7895 6749
rect 8110 6740 8116 6792
rect 8168 6740 8174 6792
rect 8220 6780 8248 6820
rect 8570 6780 8576 6792
rect 8220 6752 8576 6780
rect 8570 6740 8576 6752
rect 8628 6780 8634 6792
rect 8695 6783 8753 6789
rect 8695 6780 8707 6783
rect 8628 6752 8707 6780
rect 8628 6740 8634 6752
rect 8695 6749 8707 6752
rect 8741 6749 8753 6783
rect 8695 6743 8753 6749
rect 8849 6783 8907 6789
rect 8849 6749 8861 6783
rect 8895 6780 8907 6783
rect 8938 6780 8944 6792
rect 8895 6752 8944 6780
rect 8895 6749 8907 6752
rect 8849 6743 8907 6749
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 5534 6672 5540 6724
rect 5592 6672 5598 6724
rect 8478 6604 8484 6656
rect 8536 6604 8542 6656
rect 644 6554 9384 6576
rect 644 6502 2954 6554
rect 3006 6502 3018 6554
rect 3070 6502 3082 6554
rect 3134 6502 6954 6554
rect 7006 6502 7018 6554
rect 7070 6502 7082 6554
rect 7134 6502 9384 6554
rect 644 6480 9384 6502
rect 1118 6400 1124 6452
rect 1176 6400 1182 6452
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 5442 6440 5448 6452
rect 5132 6412 5448 6440
rect 5132 6400 5138 6412
rect 5442 6400 5448 6412
rect 5500 6440 5506 6452
rect 5500 6412 6316 6440
rect 5500 6400 5506 6412
rect 474 6264 480 6316
rect 532 6304 538 6316
rect 937 6307 995 6313
rect 937 6304 949 6307
rect 532 6276 949 6304
rect 532 6264 538 6276
rect 937 6273 949 6276
rect 983 6273 995 6307
rect 937 6267 995 6273
rect 5258 6264 5264 6316
rect 5316 6264 5322 6316
rect 5902 6264 5908 6316
rect 5960 6304 5966 6316
rect 6288 6313 6316 6412
rect 8478 6372 8484 6384
rect 8050 6344 8484 6372
rect 8478 6332 8484 6344
rect 8536 6332 8542 6384
rect 5997 6307 6055 6313
rect 5997 6304 6009 6307
rect 5960 6276 6009 6304
rect 5960 6264 5966 6276
rect 5997 6273 6009 6276
rect 6043 6273 6055 6307
rect 5997 6267 6055 6273
rect 6273 6307 6331 6313
rect 6273 6273 6285 6307
rect 6319 6273 6331 6307
rect 6273 6267 6331 6273
rect 8386 6264 8392 6316
rect 8444 6264 8450 6316
rect 3602 6196 3608 6248
rect 3660 6236 3666 6248
rect 3881 6239 3939 6245
rect 3881 6236 3893 6239
rect 3660 6208 3893 6236
rect 3660 6196 3666 6208
rect 3881 6205 3893 6208
rect 3927 6205 3939 6239
rect 3881 6199 3939 6205
rect 4157 6239 4215 6245
rect 4157 6205 4169 6239
rect 4203 6236 4215 6239
rect 4798 6236 4804 6248
rect 4203 6208 4804 6236
rect 4203 6205 4215 6208
rect 4157 6199 4215 6205
rect 4798 6196 4804 6208
rect 4856 6196 4862 6248
rect 5629 6239 5687 6245
rect 5629 6205 5641 6239
rect 5675 6236 5687 6239
rect 6086 6236 6092 6248
rect 5675 6208 6092 6236
rect 5675 6205 5687 6208
rect 5629 6199 5687 6205
rect 6086 6196 6092 6208
rect 6144 6196 6150 6248
rect 6365 6239 6423 6245
rect 6365 6205 6377 6239
rect 6411 6236 6423 6239
rect 6549 6239 6607 6245
rect 6549 6236 6561 6239
rect 6411 6208 6561 6236
rect 6411 6205 6423 6208
rect 6365 6199 6423 6205
rect 6549 6205 6561 6208
rect 6595 6205 6607 6239
rect 6549 6199 6607 6205
rect 6917 6239 6975 6245
rect 6917 6205 6929 6239
rect 6963 6236 6975 6239
rect 7190 6236 7196 6248
rect 6963 6208 7196 6236
rect 6963 6205 6975 6208
rect 6917 6199 6975 6205
rect 7190 6196 7196 6208
rect 7248 6196 7254 6248
rect 5718 6060 5724 6112
rect 5776 6100 5782 6112
rect 6178 6100 6184 6112
rect 5776 6072 6184 6100
rect 5776 6060 5782 6072
rect 6178 6060 6184 6072
rect 6236 6060 6242 6112
rect 8294 6060 8300 6112
rect 8352 6100 8358 6112
rect 8949 6103 9007 6109
rect 8949 6100 8961 6103
rect 8352 6072 8961 6100
rect 8352 6060 8358 6072
rect 8949 6069 8961 6072
rect 8995 6069 9007 6103
rect 8949 6063 9007 6069
rect 644 6010 9384 6032
rect 644 5958 2554 6010
rect 2606 5958 2618 6010
rect 2670 5958 2682 6010
rect 2734 5958 6554 6010
rect 6606 5958 6618 6010
rect 6670 5958 6682 6010
rect 6734 5958 9384 6010
rect 644 5936 9384 5958
rect 6454 5856 6460 5908
rect 6512 5896 6518 5908
rect 6549 5899 6607 5905
rect 6549 5896 6561 5899
rect 6512 5868 6561 5896
rect 6512 5856 6518 5868
rect 6549 5865 6561 5868
rect 6595 5865 6607 5899
rect 6549 5859 6607 5865
rect 8386 5856 8392 5908
rect 8444 5896 8450 5908
rect 8481 5899 8539 5905
rect 8481 5896 8493 5899
rect 8444 5868 8493 5896
rect 8444 5856 8450 5868
rect 8481 5865 8493 5868
rect 8527 5865 8539 5899
rect 8481 5859 8539 5865
rect 6362 5788 6368 5840
rect 6420 5828 6426 5840
rect 6641 5831 6699 5837
rect 6641 5828 6653 5831
rect 6420 5800 6653 5828
rect 6420 5788 6426 5800
rect 6641 5797 6653 5800
rect 6687 5797 6699 5831
rect 6641 5791 6699 5797
rect 382 5720 388 5772
rect 440 5760 446 5772
rect 1397 5763 1455 5769
rect 1397 5760 1409 5763
rect 440 5732 1409 5760
rect 440 5720 446 5732
rect 1397 5729 1409 5732
rect 1443 5729 1455 5763
rect 1397 5723 1455 5729
rect 3602 5720 3608 5772
rect 3660 5760 3666 5772
rect 4798 5760 4804 5772
rect 3660 5732 4804 5760
rect 3660 5720 3666 5732
rect 4798 5720 4804 5732
rect 4856 5720 4862 5772
rect 5077 5763 5135 5769
rect 5077 5729 5089 5763
rect 5123 5760 5135 5763
rect 6270 5760 6276 5772
rect 5123 5732 6276 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 6270 5720 6276 5732
rect 6328 5720 6334 5772
rect 7837 5763 7895 5769
rect 7837 5729 7849 5763
rect 7883 5760 7895 5763
rect 9582 5760 9588 5772
rect 7883 5732 9588 5760
rect 7883 5729 7895 5732
rect 7837 5723 7895 5729
rect 9582 5720 9588 5732
rect 9640 5720 9646 5772
rect 1118 5652 1124 5704
rect 1176 5652 1182 5704
rect 6178 5652 6184 5704
rect 6236 5692 6242 5704
rect 6825 5695 6883 5701
rect 6236 5664 6776 5692
rect 6236 5652 6242 5664
rect 6748 5624 6776 5664
rect 6825 5661 6837 5695
rect 6871 5692 6883 5695
rect 8018 5692 8024 5704
rect 6871 5664 8024 5692
rect 6871 5661 6883 5664
rect 6825 5655 6883 5661
rect 8018 5652 8024 5664
rect 8076 5652 8082 5704
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 8570 5652 8576 5704
rect 8628 5692 8634 5704
rect 8849 5695 8907 5701
rect 8849 5692 8861 5695
rect 8628 5664 8861 5692
rect 8628 5652 8634 5664
rect 8849 5661 8861 5664
rect 8895 5661 8907 5695
rect 8849 5655 8907 5661
rect 8665 5627 8723 5633
rect 8665 5624 8677 5627
rect 6748 5596 8677 5624
rect 8665 5593 8677 5596
rect 8711 5624 8723 5627
rect 8938 5624 8944 5636
rect 8711 5596 8944 5624
rect 8711 5593 8723 5596
rect 8665 5587 8723 5593
rect 8938 5584 8944 5596
rect 8996 5584 9002 5636
rect 5166 5516 5172 5568
rect 5224 5556 5230 5568
rect 9030 5556 9036 5568
rect 5224 5528 9036 5556
rect 5224 5516 5230 5528
rect 9030 5516 9036 5528
rect 9088 5516 9094 5568
rect 644 5466 9384 5488
rect 644 5414 2954 5466
rect 3006 5414 3018 5466
rect 3070 5414 3082 5466
rect 3134 5414 6954 5466
rect 7006 5414 7018 5466
rect 7070 5414 7082 5466
rect 7134 5414 9384 5466
rect 644 5392 9384 5414
rect 5721 5355 5779 5361
rect 5721 5321 5733 5355
rect 5767 5352 5779 5355
rect 5994 5352 6000 5364
rect 5767 5324 6000 5352
rect 5767 5321 5779 5324
rect 5721 5315 5779 5321
rect 5994 5312 6000 5324
rect 6052 5312 6058 5364
rect 5810 5244 5816 5296
rect 5868 5284 5874 5296
rect 5868 5256 7696 5284
rect 5868 5244 5874 5256
rect 2314 5176 2320 5228
rect 2372 5176 2378 5228
rect 6362 5176 6368 5228
rect 6420 5176 6426 5228
rect 7668 5225 7696 5256
rect 8846 5244 8852 5296
rect 8904 5244 8910 5296
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5185 7711 5219
rect 7653 5179 7711 5185
rect 934 5108 940 5160
rect 992 5108 998 5160
rect 1210 5108 1216 5160
rect 1268 5108 1274 5160
rect 2406 5108 2412 5160
rect 2464 5148 2470 5160
rect 2685 5151 2743 5157
rect 2685 5148 2697 5151
rect 2464 5120 2697 5148
rect 2464 5108 2470 5120
rect 2685 5117 2697 5120
rect 2731 5117 2743 5151
rect 2685 5111 2743 5117
rect 4154 5108 4160 5160
rect 4212 5148 4218 5160
rect 5077 5151 5135 5157
rect 5077 5148 5089 5151
rect 4212 5120 5089 5148
rect 4212 5108 4218 5120
rect 5077 5117 5089 5120
rect 5123 5117 5135 5151
rect 5077 5111 5135 5117
rect 7377 5151 7435 5157
rect 7377 5117 7389 5151
rect 7423 5148 7435 5151
rect 9582 5148 9588 5160
rect 7423 5120 9588 5148
rect 7423 5117 7435 5120
rect 7377 5111 7435 5117
rect 9582 5108 9588 5120
rect 9640 5108 9646 5160
rect 644 4922 9384 4944
rect 644 4870 2554 4922
rect 2606 4870 2618 4922
rect 2670 4870 2682 4922
rect 2734 4870 6554 4922
rect 6606 4870 6618 4922
rect 6670 4870 6682 4922
rect 6734 4870 9384 4922
rect 644 4848 9384 4870
rect 1121 4811 1179 4817
rect 1121 4777 1133 4811
rect 1167 4808 1179 4811
rect 1210 4808 1216 4820
rect 1167 4780 1216 4808
rect 1167 4777 1179 4780
rect 1121 4771 1179 4777
rect 1210 4768 1216 4780
rect 1268 4768 1274 4820
rect 4614 4768 4620 4820
rect 4672 4808 4678 4820
rect 4672 4780 8432 4808
rect 4672 4768 4678 4780
rect 2133 4743 2191 4749
rect 2133 4709 2145 4743
rect 2179 4740 2191 4743
rect 2314 4740 2320 4752
rect 2179 4712 2320 4740
rect 2179 4709 2191 4712
rect 2133 4703 2191 4709
rect 2314 4700 2320 4712
rect 2372 4700 2378 4752
rect 4249 4675 4307 4681
rect 4249 4641 4261 4675
rect 4295 4672 4307 4675
rect 4893 4675 4951 4681
rect 4893 4672 4905 4675
rect 4295 4644 4905 4672
rect 4295 4641 4307 4644
rect 4249 4635 4307 4641
rect 4893 4641 4905 4644
rect 4939 4641 4951 4675
rect 4893 4635 4951 4641
rect 6270 4632 6276 4684
rect 6328 4672 6334 4684
rect 6641 4675 6699 4681
rect 6641 4672 6653 4675
rect 6328 4644 6653 4672
rect 6328 4632 6334 4644
rect 6641 4641 6653 4644
rect 6687 4641 6699 4675
rect 6641 4635 6699 4641
rect 7837 4675 7895 4681
rect 7837 4641 7849 4675
rect 7883 4672 7895 4675
rect 8202 4672 8208 4684
rect 7883 4644 8208 4672
rect 7883 4641 7895 4644
rect 7837 4635 7895 4641
rect 8202 4632 8208 4644
rect 8260 4632 8266 4684
rect 382 4564 388 4616
rect 440 4604 446 4616
rect 937 4607 995 4613
rect 937 4604 949 4607
rect 440 4576 949 4604
rect 440 4564 446 4576
rect 937 4573 949 4576
rect 983 4573 995 4607
rect 937 4567 995 4573
rect 1397 4607 1455 4613
rect 1397 4573 1409 4607
rect 1443 4604 1455 4607
rect 2774 4604 2780 4616
rect 1443 4576 2780 4604
rect 1443 4573 1455 4576
rect 1397 4567 1455 4573
rect 2774 4564 2780 4576
rect 2832 4564 2838 4616
rect 5258 4564 5264 4616
rect 5316 4564 5322 4616
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 8404 4604 8432 4780
rect 8938 4672 8944 4684
rect 8680 4644 8944 4672
rect 8680 4613 8708 4644
rect 8938 4632 8944 4644
rect 8996 4632 9002 4684
rect 8680 4607 8753 4613
rect 8680 4604 8707 4607
rect 8404 4576 8707 4604
rect 8695 4573 8707 4576
rect 8741 4573 8753 4607
rect 8695 4567 8753 4573
rect 8849 4607 8907 4613
rect 8849 4573 8861 4607
rect 8895 4573 8907 4607
rect 8849 4567 8907 4573
rect 1946 4496 1952 4548
rect 2004 4496 2010 4548
rect 6086 4496 6092 4548
rect 6144 4536 6150 4548
rect 6365 4539 6423 4545
rect 6365 4536 6377 4539
rect 6144 4508 6377 4536
rect 6144 4496 6150 4508
rect 6365 4505 6377 4508
rect 6411 4505 6423 4539
rect 6365 4499 6423 4505
rect 8570 4496 8576 4548
rect 8628 4536 8634 4548
rect 8864 4536 8892 4567
rect 8628 4508 8892 4536
rect 8628 4496 8634 4508
rect 1118 4428 1124 4480
rect 1176 4468 1182 4480
rect 1213 4471 1271 4477
rect 1213 4468 1225 4471
rect 1176 4440 1225 4468
rect 1176 4428 1182 4440
rect 1213 4437 1225 4440
rect 1259 4437 1271 4471
rect 1213 4431 1271 4437
rect 4801 4471 4859 4477
rect 4801 4437 4813 4471
rect 4847 4468 4859 4471
rect 5350 4468 5356 4480
rect 4847 4440 5356 4468
rect 4847 4437 4859 4440
rect 4801 4431 4859 4437
rect 5350 4428 5356 4440
rect 5408 4428 5414 4480
rect 8478 4428 8484 4480
rect 8536 4428 8542 4480
rect 644 4378 9384 4400
rect 644 4326 2954 4378
rect 3006 4326 3018 4378
rect 3070 4326 3082 4378
rect 3134 4326 6954 4378
rect 7006 4326 7018 4378
rect 7070 4326 7082 4378
rect 7134 4326 9384 4378
rect 644 4304 9384 4326
rect 6273 4267 6331 4273
rect 6273 4264 6285 4267
rect 5276 4236 6285 4264
rect 5276 4208 5304 4236
rect 6273 4233 6285 4236
rect 6319 4233 6331 4267
rect 6273 4227 6331 4233
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8949 4267 9007 4273
rect 8949 4264 8961 4267
rect 8352 4236 8961 4264
rect 8352 4224 8358 4236
rect 8949 4233 8961 4236
rect 8995 4233 9007 4267
rect 8949 4227 9007 4233
rect 5258 4196 5264 4208
rect 5198 4168 5264 4196
rect 5258 4156 5264 4168
rect 5316 4156 5322 4208
rect 5350 4156 5356 4208
rect 5408 4196 5414 4208
rect 8478 4196 8484 4208
rect 5408 4168 6224 4196
rect 8050 4168 8484 4196
rect 5408 4156 5414 4168
rect 934 4088 940 4140
rect 992 4128 998 4140
rect 3602 4128 3608 4140
rect 992 4100 3608 4128
rect 992 4088 998 4100
rect 3602 4088 3608 4100
rect 3660 4128 3666 4140
rect 3697 4131 3755 4137
rect 3697 4128 3709 4131
rect 3660 4100 3709 4128
rect 3660 4088 3666 4100
rect 3697 4097 3709 4100
rect 3743 4097 3755 4131
rect 3697 4091 3755 4097
rect 5442 4088 5448 4140
rect 5500 4128 5506 4140
rect 5537 4131 5595 4137
rect 5537 4128 5549 4131
rect 5500 4100 5549 4128
rect 5500 4088 5506 4100
rect 5537 4097 5549 4100
rect 5583 4097 5595 4131
rect 5537 4091 5595 4097
rect 5994 4088 6000 4140
rect 6052 4128 6058 4140
rect 6089 4131 6147 4137
rect 6089 4128 6101 4131
rect 6052 4100 6101 4128
rect 6052 4088 6058 4100
rect 6089 4097 6101 4100
rect 6135 4097 6147 4131
rect 6196 4128 6224 4168
rect 8478 4156 8484 4168
rect 8536 4156 8542 4208
rect 6917 4131 6975 4137
rect 6917 4128 6929 4131
rect 6196 4100 6929 4128
rect 6089 4091 6147 4097
rect 6917 4097 6929 4100
rect 6963 4097 6975 4131
rect 6917 4091 6975 4097
rect 8386 4088 8392 4140
rect 8444 4088 8450 4140
rect 3973 4063 4031 4069
rect 3973 4029 3985 4063
rect 4019 4060 4031 4063
rect 5629 4063 5687 4069
rect 4019 4032 5534 4060
rect 4019 4029 4031 4032
rect 3973 4023 4031 4029
rect 5506 3992 5534 4032
rect 5629 4029 5641 4063
rect 5675 4060 5687 4063
rect 6549 4063 6607 4069
rect 6549 4060 6561 4063
rect 5675 4032 6561 4060
rect 5675 4029 5687 4032
rect 5629 4023 5687 4029
rect 6549 4029 6561 4032
rect 6595 4029 6607 4063
rect 7190 4060 7196 4072
rect 6549 4023 6607 4029
rect 6656 4032 7196 4060
rect 6656 3992 6684 4032
rect 7190 4020 7196 4032
rect 7248 4020 7254 4072
rect 5506 3964 6684 3992
rect 5258 3884 5264 3936
rect 5316 3924 5322 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 5316 3896 5457 3924
rect 5316 3884 5322 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 5445 3887 5503 3893
rect 644 3834 9384 3856
rect 644 3782 6554 3834
rect 6606 3782 6618 3834
rect 6670 3782 6682 3834
rect 6734 3782 9384 3834
rect 644 3760 9384 3782
rect 3973 3723 4031 3729
rect 3973 3689 3985 3723
rect 4019 3720 4031 3723
rect 4154 3720 4160 3732
rect 4019 3692 4160 3720
rect 4019 3689 4031 3692
rect 3973 3683 4031 3689
rect 4154 3680 4160 3692
rect 4212 3680 4218 3732
rect 4982 3680 4988 3732
rect 5040 3720 5046 3732
rect 5442 3720 5448 3732
rect 5040 3692 5448 3720
rect 5040 3680 5046 3692
rect 5442 3680 5448 3692
rect 5500 3720 5506 3732
rect 5500 3692 7972 3720
rect 5500 3680 5506 3692
rect 7650 3612 7656 3664
rect 7708 3612 7714 3664
rect 3602 3544 3608 3596
rect 3660 3584 3666 3596
rect 4890 3584 4896 3596
rect 3660 3556 4896 3584
rect 3660 3544 3666 3556
rect 4890 3544 4896 3556
rect 4948 3584 4954 3596
rect 5721 3587 5779 3593
rect 5721 3584 5733 3587
rect 4948 3556 5733 3584
rect 4948 3544 4954 3556
rect 5721 3553 5733 3556
rect 5767 3584 5779 3587
rect 5902 3584 5908 3596
rect 5767 3556 5908 3584
rect 5767 3553 5779 3556
rect 5721 3547 5779 3553
rect 5902 3544 5908 3556
rect 5960 3544 5966 3596
rect 6181 3587 6239 3593
rect 6181 3553 6193 3587
rect 6227 3584 6239 3587
rect 7190 3584 7196 3596
rect 6227 3556 7196 3584
rect 6227 3553 6239 3556
rect 6181 3547 6239 3553
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 7650 3476 7656 3528
rect 7708 3516 7714 3528
rect 7944 3525 7972 3692
rect 8386 3680 8392 3732
rect 8444 3720 8450 3732
rect 8481 3723 8539 3729
rect 8481 3720 8493 3723
rect 8444 3692 8493 3720
rect 8444 3680 8450 3692
rect 8481 3689 8493 3692
rect 8527 3689 8539 3723
rect 8481 3683 8539 3689
rect 7837 3519 7895 3525
rect 7837 3516 7849 3519
rect 7708 3488 7849 3516
rect 7708 3476 7714 3488
rect 7837 3485 7849 3488
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 7929 3519 7987 3525
rect 7929 3485 7941 3519
rect 7975 3485 7987 3519
rect 7929 3479 7987 3485
rect 8849 3519 8907 3525
rect 8849 3485 8861 3519
rect 8895 3516 8907 3519
rect 8938 3516 8944 3528
rect 8895 3488 8944 3516
rect 8895 3485 8907 3488
rect 8849 3479 8907 3485
rect 8938 3476 8944 3488
rect 8996 3476 9002 3528
rect 5014 3420 5120 3448
rect 5092 3392 5120 3420
rect 5442 3408 5448 3460
rect 5500 3408 5506 3460
rect 6270 3408 6276 3460
rect 6328 3448 6334 3460
rect 8665 3451 8723 3457
rect 6328 3420 6670 3448
rect 6328 3408 6334 3420
rect 5074 3340 5080 3392
rect 5132 3380 5138 3392
rect 6288 3380 6316 3408
rect 5132 3352 6316 3380
rect 6564 3380 6592 3420
rect 8665 3417 8677 3451
rect 8711 3417 8723 3451
rect 8665 3411 8723 3417
rect 8570 3380 8576 3392
rect 6564 3352 8576 3380
rect 5132 3340 5138 3352
rect 8570 3340 8576 3352
rect 8628 3380 8634 3392
rect 8680 3380 8708 3411
rect 8628 3352 8708 3380
rect 8628 3340 8634 3352
rect 644 3290 9384 3312
rect 644 3238 6954 3290
rect 7006 3238 7018 3290
rect 7070 3238 7082 3290
rect 7134 3238 9384 3290
rect 644 3216 9384 3238
rect 6454 3136 6460 3188
rect 6512 3176 6518 3188
rect 6512 3148 8524 3176
rect 6512 3136 6518 3148
rect 6822 3068 6828 3120
rect 6880 3068 6886 3120
rect 8496 3117 8524 3148
rect 8481 3111 8539 3117
rect 8481 3077 8493 3111
rect 8527 3077 8539 3111
rect 8481 3071 8539 3077
rect 4985 3043 5043 3049
rect 4985 3009 4997 3043
rect 5031 3040 5043 3043
rect 5156 3043 5214 3049
rect 5156 3040 5168 3043
rect 5031 3012 5168 3040
rect 5031 3009 5043 3012
rect 4985 3003 5043 3009
rect 5156 3009 5168 3012
rect 5202 3009 5214 3043
rect 5156 3003 5214 3009
rect 5718 3000 5724 3052
rect 5776 3000 5782 3052
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7561 3043 7619 3049
rect 7561 3009 7573 3043
rect 7607 3040 7619 3043
rect 7650 3040 7656 3052
rect 7607 3012 7656 3040
rect 7607 3009 7619 3012
rect 7561 3003 7619 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 8570 3000 8576 3052
rect 8628 3040 8634 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8628 3012 8677 3040
rect 8628 3000 8634 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 4525 2975 4583 2981
rect 4525 2941 4537 2975
rect 4571 2972 4583 2975
rect 5626 2972 5632 2984
rect 4571 2944 5632 2972
rect 4571 2941 4583 2944
rect 4525 2935 4583 2941
rect 5626 2932 5632 2944
rect 5684 2932 5690 2984
rect 7208 2972 7236 3000
rect 7745 2975 7803 2981
rect 7745 2972 7757 2975
rect 7208 2944 7757 2972
rect 7745 2941 7757 2944
rect 7791 2941 7803 2975
rect 7745 2935 7803 2941
rect 8294 2932 8300 2984
rect 8352 2932 8358 2984
rect 8018 2796 8024 2848
rect 8076 2836 8082 2848
rect 8849 2839 8907 2845
rect 8849 2836 8861 2839
rect 8076 2808 8861 2836
rect 8076 2796 8082 2808
rect 8849 2805 8861 2808
rect 8895 2805 8907 2839
rect 8849 2799 8907 2805
rect 2484 2746 9384 2768
rect 2484 2694 6554 2746
rect 6606 2694 6618 2746
rect 6670 2694 6682 2746
rect 6734 2694 9384 2746
rect 2484 2672 9384 2694
rect 2130 2592 2136 2644
rect 2188 2632 2194 2644
rect 2777 2635 2835 2641
rect 2777 2632 2789 2635
rect 2188 2604 2789 2632
rect 2188 2592 2194 2604
rect 2777 2601 2789 2604
rect 2823 2601 2835 2635
rect 2777 2595 2835 2601
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 5813 2635 5871 2641
rect 5813 2632 5825 2635
rect 5500 2604 5825 2632
rect 5500 2592 5506 2604
rect 5813 2601 5825 2604
rect 5859 2601 5871 2635
rect 5813 2595 5871 2601
rect 5828 2564 5856 2595
rect 6822 2592 6828 2644
rect 6880 2632 6886 2644
rect 8757 2635 8815 2641
rect 8757 2632 8769 2635
rect 6880 2604 8769 2632
rect 6880 2592 6886 2604
rect 8757 2601 8769 2604
rect 8803 2601 8815 2635
rect 8757 2595 8815 2601
rect 5828 2536 6132 2564
rect 4893 2499 4951 2505
rect 4893 2465 4905 2499
rect 4939 2496 4951 2499
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 4939 2468 6009 2496
rect 4939 2465 4951 2468
rect 4893 2459 4951 2465
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 6104 2496 6132 2536
rect 6365 2499 6423 2505
rect 6365 2496 6377 2499
rect 6104 2468 6377 2496
rect 5997 2459 6055 2465
rect 6365 2465 6377 2468
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 2958 2388 2964 2440
rect 3016 2388 3022 2440
rect 3053 2431 3111 2437
rect 3053 2397 3065 2431
rect 3099 2397 3111 2431
rect 3053 2391 3111 2397
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2428 4859 2431
rect 4982 2428 4988 2440
rect 4847 2400 4988 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 3068 2360 3096 2391
rect 4982 2388 4988 2400
rect 5040 2388 5046 2440
rect 5258 2388 5264 2440
rect 5316 2388 5322 2440
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2428 7895 2431
rect 8018 2428 8024 2440
rect 7883 2400 8024 2428
rect 7883 2397 7895 2400
rect 7837 2391 7895 2397
rect 8018 2388 8024 2400
rect 8076 2388 8082 2440
rect 8570 2388 8576 2440
rect 8628 2388 8634 2440
rect 8727 2431 8785 2437
rect 8727 2397 8739 2431
rect 8773 2428 8785 2431
rect 9030 2428 9036 2440
rect 8773 2400 9036 2428
rect 8773 2397 8785 2400
rect 8727 2391 8785 2397
rect 9030 2388 9036 2400
rect 9088 2388 9094 2440
rect 7650 2360 7656 2372
rect 2332 2332 3096 2360
rect 7498 2332 7656 2360
rect 2332 1544 2360 2332
rect 7650 2320 7656 2332
rect 7708 2320 7714 2372
rect 6822 2252 6828 2304
rect 6880 2292 6886 2304
rect 8397 2295 8455 2301
rect 8397 2292 8409 2295
rect 6880 2264 8409 2292
rect 6880 2252 6886 2264
rect 8397 2261 8409 2264
rect 8443 2261 8455 2295
rect 8397 2255 8455 2261
rect 2484 2202 9384 2224
rect 2484 2150 6954 2202
rect 7006 2150 7018 2202
rect 7070 2150 7082 2202
rect 7134 2150 9384 2202
rect 2484 2128 9384 2150
rect 6822 2088 6828 2100
rect 4816 2060 6828 2088
rect 4816 2020 4844 2060
rect 6822 2048 6828 2060
rect 6880 2048 6886 2100
rect 7193 2091 7251 2097
rect 7193 2057 7205 2091
rect 7239 2088 7251 2091
rect 7650 2088 7656 2100
rect 7239 2060 7656 2088
rect 7239 2057 7251 2060
rect 7193 2051 7251 2057
rect 7650 2048 7656 2060
rect 7708 2048 7714 2100
rect 4724 1992 4844 2020
rect 4724 1961 4752 1992
rect 5166 1980 5172 2032
rect 5224 1980 5230 2032
rect 6454 1980 6460 2032
rect 6512 2020 6518 2032
rect 8665 2023 8723 2029
rect 6512 1992 6960 2020
rect 6512 1980 6518 1992
rect 4709 1955 4767 1961
rect 4709 1921 4721 1955
rect 4755 1921 4767 1955
rect 4709 1915 4767 1921
rect 4890 1912 4896 1964
rect 4948 1912 4954 1964
rect 6270 1912 6276 1964
rect 6328 1952 6334 1964
rect 6932 1961 6960 1992
rect 8665 1989 8677 2023
rect 8711 2020 8723 2023
rect 9030 2020 9036 2032
rect 8711 1992 9036 2020
rect 8711 1989 8723 1992
rect 8665 1983 8723 1989
rect 9030 1980 9036 1992
rect 9088 1980 9094 2032
rect 6825 1955 6883 1961
rect 6825 1952 6837 1955
rect 6328 1924 6837 1952
rect 6328 1912 6334 1924
rect 6825 1921 6837 1924
rect 6871 1921 6883 1955
rect 6825 1915 6883 1921
rect 6918 1955 6976 1961
rect 6918 1921 6930 1955
rect 6964 1921 6976 1955
rect 6918 1915 6976 1921
rect 8570 1912 8576 1964
rect 8628 1952 8634 1964
rect 8849 1955 8907 1961
rect 8849 1952 8861 1955
rect 8628 1924 8861 1952
rect 8628 1912 8634 1924
rect 8849 1921 8861 1924
rect 8895 1921 8907 1955
rect 8849 1915 8907 1921
rect 4341 1887 4399 1893
rect 4341 1853 4353 1887
rect 4387 1884 4399 1887
rect 9582 1884 9588 1896
rect 4387 1856 9588 1884
rect 4387 1853 4399 1856
rect 4341 1847 4399 1853
rect 9582 1844 9588 1856
rect 9640 1844 9646 1896
rect 6641 1819 6699 1825
rect 6641 1785 6653 1819
rect 6687 1816 6699 1819
rect 8294 1816 8300 1828
rect 6687 1788 8300 1816
rect 6687 1785 6699 1788
rect 6641 1779 6699 1785
rect 8294 1776 8300 1788
rect 8352 1776 8358 1828
rect 5718 1708 5724 1760
rect 5776 1748 5782 1760
rect 9033 1751 9091 1757
rect 9033 1748 9045 1751
rect 5776 1720 9045 1748
rect 5776 1708 5782 1720
rect 9033 1717 9045 1720
rect 9079 1717 9091 1751
rect 9033 1711 9091 1717
rect 2484 1658 9384 1680
rect 2484 1606 6554 1658
rect 6606 1606 6618 1658
rect 6670 1606 6682 1658
rect 6734 1606 9384 1658
rect 2484 1584 9384 1606
rect 1702 1516 2360 1544
rect 2958 1504 2964 1556
rect 3016 1544 3022 1556
rect 8849 1547 8907 1553
rect 8849 1544 8861 1547
rect 3016 1516 8861 1544
rect 3016 1504 3022 1516
rect 8849 1513 8861 1516
rect 8895 1513 8907 1547
rect 8849 1507 8907 1513
rect 7377 1411 7435 1417
rect 7377 1377 7389 1411
rect 7423 1408 7435 1411
rect 9122 1408 9128 1420
rect 7423 1380 9128 1408
rect 7423 1377 7435 1380
rect 7377 1371 7435 1377
rect 9122 1368 9128 1380
rect 9180 1368 9186 1420
rect 6365 1343 6423 1349
rect 6365 1309 6377 1343
rect 6411 1340 6423 1343
rect 7650 1340 7656 1352
rect 6411 1312 7656 1340
rect 6411 1309 6423 1312
rect 6365 1303 6423 1309
rect 7650 1300 7656 1312
rect 7708 1300 7714 1352
rect 9030 1300 9036 1352
rect 9088 1300 9094 1352
rect 2484 1114 9384 1136
rect 2484 1062 6954 1114
rect 7006 1062 7018 1114
rect 7070 1062 7082 1114
rect 7134 1062 9384 1114
rect 2484 1040 9384 1062
<< via1 >>
rect 5356 14288 5408 14340
rect 7104 14288 7156 14340
rect 3240 14220 3292 14272
rect 8024 14220 8076 14272
rect 2954 14118 3006 14170
rect 3018 14118 3070 14170
rect 3082 14118 3134 14170
rect 6954 14118 7006 14170
rect 7018 14118 7070 14170
rect 7082 14118 7134 14170
rect 6828 14016 6880 14068
rect 4804 13948 4856 14000
rect 9588 13948 9640 14000
rect 3240 13880 3292 13932
rect 4436 13923 4488 13932
rect 4436 13889 4445 13923
rect 4445 13889 4479 13923
rect 4479 13889 4488 13923
rect 4436 13880 4488 13889
rect 6276 13880 6328 13932
rect 8116 13923 8168 13932
rect 8116 13889 8125 13923
rect 8125 13889 8159 13923
rect 8159 13889 8168 13923
rect 8116 13880 8168 13889
rect 8576 13880 8628 13932
rect 6460 13812 6512 13864
rect 3976 13744 4028 13796
rect 5632 13744 5684 13796
rect 940 13676 992 13728
rect 1676 13676 1728 13728
rect 4896 13676 4948 13728
rect 5908 13719 5960 13728
rect 5908 13685 5917 13719
rect 5917 13685 5951 13719
rect 5951 13685 5960 13719
rect 5908 13676 5960 13685
rect 8484 13744 8536 13796
rect 7196 13676 7248 13728
rect 8576 13676 8628 13728
rect 8852 13719 8904 13728
rect 8852 13685 8861 13719
rect 8861 13685 8895 13719
rect 8895 13685 8904 13719
rect 8852 13676 8904 13685
rect 2554 13574 2606 13626
rect 2618 13574 2670 13626
rect 2682 13574 2734 13626
rect 6554 13574 6606 13626
rect 6618 13574 6670 13626
rect 6682 13574 6734 13626
rect 1860 13472 1912 13524
rect 5724 13472 5776 13524
rect 6184 13472 6236 13524
rect 8852 13472 8904 13524
rect 5908 13404 5960 13456
rect 940 13311 992 13320
rect 940 13277 949 13311
rect 949 13277 983 13311
rect 983 13277 992 13311
rect 940 13268 992 13277
rect 1860 13311 1912 13320
rect 1860 13277 1869 13311
rect 1869 13277 1903 13311
rect 1903 13277 1912 13311
rect 1860 13268 1912 13277
rect 2412 13268 2464 13320
rect 3240 13268 3292 13320
rect 5356 13379 5408 13388
rect 5356 13345 5365 13379
rect 5365 13345 5399 13379
rect 5399 13345 5408 13379
rect 5356 13336 5408 13345
rect 4528 13268 4580 13320
rect 7656 13404 7708 13456
rect 9588 13404 9640 13456
rect 8576 13336 8628 13388
rect 6460 13268 6512 13320
rect 7656 13268 7708 13320
rect 1124 13175 1176 13184
rect 1124 13141 1133 13175
rect 1133 13141 1167 13175
rect 1167 13141 1176 13175
rect 1124 13132 1176 13141
rect 1400 13175 1452 13184
rect 1400 13141 1409 13175
rect 1409 13141 1443 13175
rect 1443 13141 1452 13175
rect 1400 13132 1452 13141
rect 1584 13132 1636 13184
rect 2044 13132 2096 13184
rect 2780 13132 2832 13184
rect 5080 13200 5132 13252
rect 6368 13200 6420 13252
rect 8576 13200 8628 13252
rect 8852 13311 8904 13320
rect 8852 13277 8861 13311
rect 8861 13277 8895 13311
rect 8895 13277 8904 13311
rect 8852 13268 8904 13277
rect 9128 13200 9180 13252
rect 4068 13132 4120 13184
rect 8208 13132 8260 13184
rect 2954 13030 3006 13082
rect 3018 13030 3070 13082
rect 3082 13030 3134 13082
rect 6954 13030 7006 13082
rect 7018 13030 7070 13082
rect 7082 13030 7134 13082
rect 940 12835 992 12844
rect 940 12801 949 12835
rect 949 12801 983 12835
rect 983 12801 992 12835
rect 940 12792 992 12801
rect 1216 12792 1268 12844
rect 3240 12928 3292 12980
rect 8300 12928 8352 12980
rect 4160 12860 4212 12912
rect 4528 12792 4580 12844
rect 5080 12835 5132 12844
rect 5080 12801 5089 12835
rect 5089 12801 5123 12835
rect 5123 12801 5132 12835
rect 5080 12792 5132 12801
rect 6368 12860 6420 12912
rect 7656 12860 7708 12912
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 1492 12724 1544 12776
rect 3240 12656 3292 12708
rect 5816 12588 5868 12640
rect 6092 12631 6144 12640
rect 6092 12597 6101 12631
rect 6101 12597 6135 12631
rect 6135 12597 6144 12631
rect 6092 12588 6144 12597
rect 8392 12835 8444 12844
rect 8392 12801 8401 12835
rect 8401 12801 8435 12835
rect 8435 12801 8444 12835
rect 8392 12792 8444 12801
rect 6828 12724 6880 12776
rect 7196 12724 7248 12776
rect 8668 12588 8720 12640
rect 8944 12631 8996 12640
rect 8944 12597 8961 12631
rect 8961 12597 8995 12631
rect 8995 12597 8996 12631
rect 8944 12588 8996 12597
rect 2554 12486 2606 12538
rect 2618 12486 2670 12538
rect 2682 12486 2734 12538
rect 6554 12486 6606 12538
rect 6618 12486 6670 12538
rect 6682 12486 6734 12538
rect 1216 12427 1268 12436
rect 1216 12393 1225 12427
rect 1225 12393 1259 12427
rect 1259 12393 1268 12427
rect 1216 12384 1268 12393
rect 1492 12384 1544 12436
rect 2780 12384 2832 12436
rect 2412 12248 2464 12300
rect 1400 12180 1452 12232
rect 4160 12316 4212 12368
rect 6000 12384 6052 12436
rect 6276 12384 6328 12436
rect 6460 12384 6512 12436
rect 2320 12112 2372 12164
rect 2780 12112 2832 12164
rect 4252 12180 4304 12232
rect 4620 12180 4672 12232
rect 5080 12223 5132 12232
rect 5080 12189 5089 12223
rect 5089 12189 5123 12223
rect 5123 12189 5132 12223
rect 5080 12180 5132 12189
rect 6276 12180 6328 12232
rect 4160 12112 4212 12164
rect 6092 12112 6144 12164
rect 6368 12112 6420 12164
rect 3608 12044 3660 12096
rect 4528 12044 4580 12096
rect 5540 12044 5592 12096
rect 8024 12223 8076 12232
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8760 12223 8812 12232
rect 8760 12189 8768 12223
rect 8768 12189 8802 12223
rect 8802 12189 8812 12223
rect 8760 12180 8812 12189
rect 9128 12180 9180 12232
rect 8484 12087 8536 12096
rect 8484 12053 8493 12087
rect 8493 12053 8527 12087
rect 8527 12053 8536 12087
rect 8484 12044 8536 12053
rect 2954 11942 3006 11994
rect 3018 11942 3070 11994
rect 3082 11942 3134 11994
rect 6954 11942 7006 11994
rect 7018 11942 7070 11994
rect 7082 11942 7134 11994
rect 940 11883 992 11892
rect 940 11849 949 11883
rect 949 11849 983 11883
rect 983 11849 992 11883
rect 940 11840 992 11849
rect 1676 11840 1728 11892
rect 2412 11840 2464 11892
rect 2320 11772 2372 11824
rect 3240 11840 3292 11892
rect 7656 11840 7708 11892
rect 8116 11840 8168 11892
rect 4528 11772 4580 11824
rect 8484 11772 8536 11824
rect 2412 11679 2464 11688
rect 2412 11645 2421 11679
rect 2421 11645 2455 11679
rect 2455 11645 2464 11679
rect 2412 11636 2464 11645
rect 2320 11500 2372 11552
rect 3240 11500 3292 11552
rect 4068 11500 4120 11552
rect 4712 11500 4764 11552
rect 5080 11500 5132 11552
rect 6000 11747 6052 11756
rect 6000 11713 6010 11747
rect 6010 11713 6044 11747
rect 6044 11713 6052 11747
rect 6000 11704 6052 11713
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 8208 11747 8260 11756
rect 8208 11713 8217 11747
rect 8217 11713 8251 11747
rect 8251 11713 8260 11747
rect 8208 11704 8260 11713
rect 6092 11636 6144 11688
rect 6460 11636 6512 11688
rect 6000 11568 6052 11620
rect 9036 11500 9088 11552
rect 2554 11398 2606 11450
rect 2618 11398 2670 11450
rect 2682 11398 2734 11450
rect 6554 11398 6606 11450
rect 6618 11398 6670 11450
rect 6682 11398 6734 11450
rect 2780 11296 2832 11348
rect 4620 11296 4672 11348
rect 7196 11296 7248 11348
rect 2412 11228 2464 11280
rect 1400 11160 1452 11212
rect 2136 11135 2188 11144
rect 2136 11101 2145 11135
rect 2145 11101 2179 11135
rect 2179 11101 2188 11135
rect 2136 11092 2188 11101
rect 2228 11092 2280 11144
rect 4068 11160 4120 11212
rect 5356 11135 5408 11144
rect 5356 11101 5365 11135
rect 5365 11101 5399 11135
rect 5399 11101 5408 11135
rect 5356 11092 5408 11101
rect 1032 11067 1084 11076
rect 1032 11033 1041 11067
rect 1041 11033 1075 11067
rect 1075 11033 1084 11067
rect 1032 11024 1084 11033
rect 1676 11024 1728 11076
rect 5172 11024 5224 11076
rect 8760 11160 8812 11212
rect 6276 11135 6328 11144
rect 6276 11101 6285 11135
rect 6285 11101 6319 11135
rect 6319 11101 6328 11135
rect 6276 11092 6328 11101
rect 8116 11067 8168 11076
rect 8116 11033 8125 11067
rect 8125 11033 8159 11067
rect 8159 11033 8168 11067
rect 8116 11024 8168 11033
rect 9128 11024 9180 11076
rect 8484 10999 8536 11008
rect 8484 10965 8493 10999
rect 8493 10965 8527 10999
rect 8527 10965 8536 10999
rect 8484 10956 8536 10965
rect 2954 10854 3006 10906
rect 3018 10854 3070 10906
rect 3082 10854 3134 10906
rect 6954 10854 7006 10906
rect 7018 10854 7070 10906
rect 7082 10854 7134 10906
rect 4068 10752 4120 10804
rect 5356 10752 5408 10804
rect 8300 10752 8352 10804
rect 480 10684 532 10736
rect 1400 10684 1452 10736
rect 1768 10684 1820 10736
rect 5632 10727 5684 10736
rect 5632 10693 5641 10727
rect 5641 10693 5675 10727
rect 5675 10693 5684 10727
rect 5632 10684 5684 10693
rect 6000 10684 6052 10736
rect 8208 10684 8260 10736
rect 1676 10548 1728 10600
rect 2228 10591 2280 10600
rect 2228 10557 2237 10591
rect 2237 10557 2271 10591
rect 2271 10557 2280 10591
rect 2228 10548 2280 10557
rect 2044 10412 2096 10464
rect 4160 10616 4212 10668
rect 4528 10616 4580 10668
rect 5356 10616 5408 10668
rect 5540 10616 5592 10668
rect 6184 10616 6236 10668
rect 8484 10616 8536 10668
rect 3608 10548 3660 10600
rect 5724 10548 5776 10600
rect 6184 10480 6236 10532
rect 4344 10412 4396 10464
rect 4988 10412 5040 10464
rect 8668 10480 8720 10532
rect 8300 10412 8352 10464
rect 2554 10310 2606 10362
rect 2618 10310 2670 10362
rect 2682 10310 2734 10362
rect 6554 10310 6606 10362
rect 6618 10310 6670 10362
rect 6682 10310 6734 10362
rect 2044 10251 2096 10260
rect 2044 10217 2053 10251
rect 2053 10217 2087 10251
rect 2087 10217 2096 10251
rect 2044 10208 2096 10217
rect 2228 10208 2280 10260
rect 3608 10208 3660 10260
rect 5724 10251 5776 10260
rect 5724 10217 5733 10251
rect 5733 10217 5767 10251
rect 5767 10217 5776 10251
rect 5724 10208 5776 10217
rect 5172 10183 5224 10192
rect 5172 10149 5181 10183
rect 5181 10149 5215 10183
rect 5215 10149 5224 10183
rect 5172 10140 5224 10149
rect 480 10072 532 10124
rect 2228 10047 2280 10056
rect 2228 10013 2237 10047
rect 2237 10013 2271 10047
rect 2271 10013 2280 10047
rect 2228 10004 2280 10013
rect 2780 10004 2832 10056
rect 5080 10047 5132 10056
rect 5080 10013 5089 10047
rect 5089 10013 5123 10047
rect 5123 10013 5132 10047
rect 5080 10004 5132 10013
rect 5632 10140 5684 10192
rect 5908 10140 5960 10192
rect 7656 10140 7708 10192
rect 8208 10140 8260 10192
rect 5540 10047 5592 10056
rect 5540 10013 5549 10047
rect 5549 10013 5583 10047
rect 5583 10013 5592 10047
rect 5540 10004 5592 10013
rect 5632 10047 5684 10056
rect 5632 10013 5641 10047
rect 5641 10013 5675 10047
rect 5675 10013 5684 10047
rect 5632 10004 5684 10013
rect 1952 9936 2004 9988
rect 4160 9936 4212 9988
rect 5172 9936 5224 9988
rect 6000 10004 6052 10056
rect 6460 10004 6512 10056
rect 9588 10072 9640 10124
rect 8024 10004 8076 10056
rect 8300 10047 8352 10056
rect 8300 10013 8309 10047
rect 8309 10013 8343 10047
rect 8343 10013 8352 10047
rect 8300 10004 8352 10013
rect 8760 10047 8812 10056
rect 8760 10013 8768 10047
rect 8768 10013 8802 10047
rect 8802 10013 8812 10047
rect 8760 10004 8812 10013
rect 9128 10004 9180 10056
rect 6368 9936 6420 9988
rect 6460 9868 6512 9920
rect 2954 9766 3006 9818
rect 3018 9766 3070 9818
rect 3082 9766 3134 9818
rect 6954 9766 7006 9818
rect 7018 9766 7070 9818
rect 7082 9766 7134 9818
rect 1676 9664 1728 9716
rect 2044 9596 2096 9648
rect 3608 9664 3660 9716
rect 4160 9664 4212 9716
rect 6276 9664 6328 9716
rect 3240 9528 3292 9580
rect 1676 9460 1728 9512
rect 2320 9460 2372 9512
rect 2780 9435 2832 9444
rect 2780 9401 2789 9435
rect 2789 9401 2823 9435
rect 2823 9401 2832 9435
rect 2780 9392 2832 9401
rect 4344 9596 4396 9648
rect 5540 9596 5592 9648
rect 9128 9664 9180 9716
rect 5356 9528 5408 9580
rect 8484 9596 8536 9648
rect 6368 9571 6420 9580
rect 6368 9537 6377 9571
rect 6377 9537 6411 9571
rect 6411 9537 6420 9571
rect 6368 9528 6420 9537
rect 8208 9571 8260 9580
rect 8208 9537 8217 9571
rect 8217 9537 8251 9571
rect 8251 9537 8260 9571
rect 8208 9528 8260 9537
rect 3976 9503 4028 9512
rect 3976 9469 3985 9503
rect 3985 9469 4019 9503
rect 4019 9469 4028 9503
rect 3976 9460 4028 9469
rect 4620 9460 4672 9512
rect 6460 9460 6512 9512
rect 1860 9324 1912 9376
rect 4252 9324 4304 9376
rect 4896 9324 4948 9376
rect 7196 9324 7248 9376
rect 8116 9324 8168 9376
rect 2554 9222 2606 9274
rect 2618 9222 2670 9274
rect 2682 9222 2734 9274
rect 6554 9222 6606 9274
rect 6618 9222 6670 9274
rect 6682 9222 6734 9274
rect 2136 9120 2188 9172
rect 6368 9120 6420 9172
rect 6460 9120 6512 9172
rect 2044 9052 2096 9104
rect 2780 9052 2832 9104
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 388 8848 440 8900
rect 1216 8848 1268 8900
rect 2044 8848 2096 8900
rect 3240 8916 3292 8968
rect 4068 9052 4120 9104
rect 5172 9052 5224 9104
rect 6828 9120 6880 9172
rect 3976 8984 4028 9036
rect 4896 8984 4948 9036
rect 5080 8984 5132 9036
rect 4988 8916 5040 8968
rect 5356 8916 5408 8968
rect 8484 9095 8536 9104
rect 8484 9061 8493 9095
rect 8493 9061 8527 9095
rect 8527 9061 8536 9095
rect 8484 9052 8536 9061
rect 7196 8916 7248 8968
rect 8024 8984 8076 9036
rect 7656 8959 7708 8968
rect 7656 8925 7665 8959
rect 7665 8925 7699 8959
rect 7699 8925 7708 8959
rect 7656 8916 7708 8925
rect 8760 8959 8812 8968
rect 2412 8780 2464 8832
rect 5172 8848 5224 8900
rect 6184 8848 6236 8900
rect 8760 8925 8771 8959
rect 8771 8925 8812 8959
rect 8760 8916 8812 8925
rect 9128 8916 9180 8968
rect 6828 8780 6880 8832
rect 8116 8780 8168 8832
rect 2954 8678 3006 8730
rect 3018 8678 3070 8730
rect 3082 8678 3134 8730
rect 6954 8678 7006 8730
rect 7018 8678 7070 8730
rect 7082 8678 7134 8730
rect 1768 8576 1820 8628
rect 5080 8576 5132 8628
rect 5632 8576 5684 8628
rect 5724 8576 5776 8628
rect 6460 8576 6512 8628
rect 2412 8508 2464 8560
rect 3240 8508 3292 8560
rect 5908 8508 5960 8560
rect 7656 8508 7708 8560
rect 1032 8483 1084 8492
rect 1032 8449 1041 8483
rect 1041 8449 1075 8483
rect 1075 8449 1084 8483
rect 1032 8440 1084 8449
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 3608 8440 3660 8492
rect 6368 8483 6420 8492
rect 6368 8449 6377 8483
rect 6377 8449 6411 8483
rect 6411 8449 6420 8483
rect 6368 8440 6420 8449
rect 7196 8440 7248 8492
rect 8668 8440 8720 8492
rect 8944 8483 8996 8492
rect 8944 8449 8953 8483
rect 8953 8449 8987 8483
rect 8987 8449 8996 8483
rect 8944 8440 8996 8449
rect 6460 8372 6512 8424
rect 9588 8372 9640 8424
rect 4344 8304 4396 8356
rect 2044 8236 2096 8288
rect 2228 8236 2280 8288
rect 3608 8236 3660 8288
rect 7196 8236 7248 8288
rect 7656 8236 7708 8288
rect 2554 8134 2606 8186
rect 2618 8134 2670 8186
rect 2682 8134 2734 8186
rect 6554 8134 6606 8186
rect 6618 8134 6670 8186
rect 6682 8134 6734 8186
rect 4436 8032 4488 8084
rect 8208 8032 8260 8084
rect 5908 7964 5960 8016
rect 3608 7896 3660 7948
rect 8392 7896 8444 7948
rect 2780 7828 2832 7880
rect 3240 7828 3292 7880
rect 6092 7871 6144 7880
rect 6092 7837 6101 7871
rect 6101 7837 6135 7871
rect 6135 7837 6144 7871
rect 6092 7828 6144 7837
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 8760 7828 8812 7880
rect 1124 7760 1176 7812
rect 5632 7803 5684 7812
rect 1308 7735 1360 7744
rect 1308 7701 1317 7735
rect 1317 7701 1351 7735
rect 1351 7701 1360 7735
rect 1308 7692 1360 7701
rect 2228 7735 2280 7744
rect 2228 7701 2237 7735
rect 2237 7701 2271 7735
rect 2271 7701 2280 7735
rect 2228 7692 2280 7701
rect 2320 7692 2372 7744
rect 5632 7769 5641 7803
rect 5641 7769 5675 7803
rect 5675 7769 5684 7803
rect 5632 7760 5684 7769
rect 5724 7760 5776 7812
rect 6276 7760 6328 7812
rect 9128 7760 9180 7812
rect 4804 7692 4856 7744
rect 6368 7692 6420 7744
rect 2954 7590 3006 7642
rect 3018 7590 3070 7642
rect 3082 7590 3134 7642
rect 6954 7590 7006 7642
rect 7018 7590 7070 7642
rect 7082 7590 7134 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 3240 7488 3292 7540
rect 8300 7488 8352 7540
rect 2228 7420 2280 7472
rect 4712 7420 4764 7472
rect 6828 7420 6880 7472
rect 8668 7463 8720 7472
rect 8668 7429 8677 7463
rect 8677 7429 8711 7463
rect 8711 7429 8720 7463
rect 8668 7420 8720 7429
rect 940 7395 992 7404
rect 940 7361 949 7395
rect 949 7361 983 7395
rect 983 7361 992 7395
rect 940 7352 992 7361
rect 1216 7395 1268 7404
rect 1216 7361 1225 7395
rect 1225 7361 1259 7395
rect 1259 7361 1268 7395
rect 1216 7352 1268 7361
rect 1676 7284 1728 7336
rect 2412 7284 2464 7336
rect 2044 7216 2096 7268
rect 2320 7216 2372 7268
rect 4896 7395 4948 7404
rect 4896 7361 4905 7395
rect 4905 7361 4939 7395
rect 4939 7361 4948 7395
rect 4896 7352 4948 7361
rect 5080 7395 5132 7404
rect 5080 7361 5089 7395
rect 5089 7361 5123 7395
rect 5123 7361 5132 7395
rect 5080 7352 5132 7361
rect 5632 7395 5684 7404
rect 5632 7361 5640 7395
rect 5640 7361 5674 7395
rect 5674 7361 5684 7395
rect 5632 7352 5684 7361
rect 5724 7395 5776 7404
rect 5724 7361 5733 7395
rect 5733 7361 5767 7395
rect 5767 7361 5776 7395
rect 5724 7352 5776 7361
rect 6276 7352 6328 7404
rect 8944 7352 8996 7404
rect 5448 7216 5500 7268
rect 5908 7216 5960 7268
rect 5540 7191 5592 7200
rect 5540 7157 5549 7191
rect 5549 7157 5583 7191
rect 5583 7157 5592 7191
rect 5540 7148 5592 7157
rect 7196 7148 7248 7200
rect 7656 7148 7708 7200
rect 2554 7046 2606 7098
rect 2618 7046 2670 7098
rect 2682 7046 2734 7098
rect 6554 7046 6606 7098
rect 6618 7046 6670 7098
rect 6682 7046 6734 7098
rect 4068 6944 4120 6996
rect 6184 6944 6236 6996
rect 8576 6944 8628 6996
rect 5080 6808 5132 6860
rect 7656 6876 7708 6928
rect 4804 6740 4856 6792
rect 6368 6783 6420 6792
rect 6368 6749 6377 6783
rect 6377 6749 6411 6783
rect 6411 6749 6420 6783
rect 6368 6740 6420 6749
rect 7656 6740 7708 6792
rect 8116 6783 8168 6792
rect 8116 6749 8125 6783
rect 8125 6749 8159 6783
rect 8159 6749 8168 6783
rect 8116 6740 8168 6749
rect 8576 6740 8628 6792
rect 8944 6740 8996 6792
rect 5540 6672 5592 6724
rect 8484 6647 8536 6656
rect 8484 6613 8493 6647
rect 8493 6613 8527 6647
rect 8527 6613 8536 6647
rect 8484 6604 8536 6613
rect 2954 6502 3006 6554
rect 3018 6502 3070 6554
rect 3082 6502 3134 6554
rect 6954 6502 7006 6554
rect 7018 6502 7070 6554
rect 7082 6502 7134 6554
rect 1124 6443 1176 6452
rect 1124 6409 1133 6443
rect 1133 6409 1167 6443
rect 1167 6409 1176 6443
rect 1124 6400 1176 6409
rect 5080 6400 5132 6452
rect 5448 6400 5500 6452
rect 480 6264 532 6316
rect 5264 6264 5316 6316
rect 5908 6264 5960 6316
rect 8484 6332 8536 6384
rect 8392 6307 8444 6316
rect 8392 6273 8401 6307
rect 8401 6273 8435 6307
rect 8435 6273 8444 6307
rect 8392 6264 8444 6273
rect 3608 6196 3660 6248
rect 4804 6196 4856 6248
rect 6092 6196 6144 6248
rect 7196 6196 7248 6248
rect 5724 6060 5776 6112
rect 6184 6103 6236 6112
rect 6184 6069 6193 6103
rect 6193 6069 6227 6103
rect 6227 6069 6236 6103
rect 6184 6060 6236 6069
rect 8300 6060 8352 6112
rect 2554 5958 2606 6010
rect 2618 5958 2670 6010
rect 2682 5958 2734 6010
rect 6554 5958 6606 6010
rect 6618 5958 6670 6010
rect 6682 5958 6734 6010
rect 6460 5856 6512 5908
rect 8392 5856 8444 5908
rect 6368 5788 6420 5840
rect 388 5720 440 5772
rect 3608 5720 3660 5772
rect 4804 5763 4856 5772
rect 4804 5729 4813 5763
rect 4813 5729 4847 5763
rect 4847 5729 4856 5763
rect 4804 5720 4856 5729
rect 6276 5720 6328 5772
rect 9588 5720 9640 5772
rect 1124 5695 1176 5704
rect 1124 5661 1133 5695
rect 1133 5661 1167 5695
rect 1167 5661 1176 5695
rect 1124 5652 1176 5661
rect 6184 5652 6236 5704
rect 8024 5652 8076 5704
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 8576 5652 8628 5704
rect 8944 5584 8996 5636
rect 5172 5516 5224 5568
rect 9036 5516 9088 5568
rect 2954 5414 3006 5466
rect 3018 5414 3070 5466
rect 3082 5414 3134 5466
rect 6954 5414 7006 5466
rect 7018 5414 7070 5466
rect 7082 5414 7134 5466
rect 6000 5312 6052 5364
rect 5816 5244 5868 5296
rect 2320 5176 2372 5228
rect 6368 5219 6420 5228
rect 6368 5185 6377 5219
rect 6377 5185 6411 5219
rect 6411 5185 6420 5219
rect 6368 5176 6420 5185
rect 8852 5287 8904 5296
rect 8852 5253 8861 5287
rect 8861 5253 8895 5287
rect 8895 5253 8904 5287
rect 8852 5244 8904 5253
rect 940 5151 992 5160
rect 940 5117 949 5151
rect 949 5117 983 5151
rect 983 5117 992 5151
rect 940 5108 992 5117
rect 1216 5151 1268 5160
rect 1216 5117 1225 5151
rect 1225 5117 1259 5151
rect 1259 5117 1268 5151
rect 1216 5108 1268 5117
rect 2412 5108 2464 5160
rect 4160 5108 4212 5160
rect 9588 5108 9640 5160
rect 2554 4870 2606 4922
rect 2618 4870 2670 4922
rect 2682 4870 2734 4922
rect 6554 4870 6606 4922
rect 6618 4870 6670 4922
rect 6682 4870 6734 4922
rect 1216 4768 1268 4820
rect 4620 4768 4672 4820
rect 2320 4700 2372 4752
rect 6276 4632 6328 4684
rect 8208 4632 8260 4684
rect 388 4564 440 4616
rect 2780 4564 2832 4616
rect 5264 4564 5316 4616
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 8944 4632 8996 4684
rect 1952 4539 2004 4548
rect 1952 4505 1961 4539
rect 1961 4505 1995 4539
rect 1995 4505 2004 4539
rect 1952 4496 2004 4505
rect 6092 4496 6144 4548
rect 8576 4496 8628 4548
rect 1124 4428 1176 4480
rect 5356 4428 5408 4480
rect 8484 4471 8536 4480
rect 8484 4437 8493 4471
rect 8493 4437 8527 4471
rect 8527 4437 8536 4471
rect 8484 4428 8536 4437
rect 2954 4326 3006 4378
rect 3018 4326 3070 4378
rect 3082 4326 3134 4378
rect 6954 4326 7006 4378
rect 7018 4326 7070 4378
rect 7082 4326 7134 4378
rect 8300 4224 8352 4276
rect 5264 4156 5316 4208
rect 5356 4156 5408 4208
rect 940 4088 992 4140
rect 3608 4088 3660 4140
rect 5448 4088 5500 4140
rect 6000 4088 6052 4140
rect 8484 4156 8536 4208
rect 8392 4131 8444 4140
rect 8392 4097 8401 4131
rect 8401 4097 8435 4131
rect 8435 4097 8444 4131
rect 8392 4088 8444 4097
rect 7196 4020 7248 4072
rect 5264 3884 5316 3936
rect 6554 3782 6606 3834
rect 6618 3782 6670 3834
rect 6682 3782 6734 3834
rect 4160 3680 4212 3732
rect 4988 3680 5040 3732
rect 5448 3680 5500 3732
rect 7656 3655 7708 3664
rect 7656 3621 7665 3655
rect 7665 3621 7699 3655
rect 7699 3621 7708 3655
rect 7656 3612 7708 3621
rect 3608 3544 3660 3596
rect 4896 3544 4948 3596
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 7196 3544 7248 3596
rect 7656 3476 7708 3528
rect 8392 3680 8444 3732
rect 8944 3476 8996 3528
rect 5448 3451 5500 3460
rect 5448 3417 5457 3451
rect 5457 3417 5491 3451
rect 5491 3417 5500 3451
rect 5448 3408 5500 3417
rect 6276 3408 6328 3460
rect 5080 3340 5132 3392
rect 8576 3340 8628 3392
rect 6954 3238 7006 3290
rect 7018 3238 7070 3290
rect 7082 3238 7134 3290
rect 6460 3136 6512 3188
rect 6828 3068 6880 3120
rect 5724 3043 5776 3052
rect 5724 3009 5733 3043
rect 5733 3009 5767 3043
rect 5767 3009 5776 3043
rect 5724 3000 5776 3009
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7656 3000 7708 3052
rect 8576 3000 8628 3052
rect 5632 2932 5684 2984
rect 8300 2975 8352 2984
rect 8300 2941 8309 2975
rect 8309 2941 8343 2975
rect 8343 2941 8352 2975
rect 8300 2932 8352 2941
rect 8024 2796 8076 2848
rect 6554 2694 6606 2746
rect 6618 2694 6670 2746
rect 6682 2694 6734 2746
rect 2136 2592 2188 2644
rect 5448 2592 5500 2644
rect 6828 2592 6880 2644
rect 2964 2431 3016 2440
rect 2964 2397 2973 2431
rect 2973 2397 3007 2431
rect 3007 2397 3016 2431
rect 2964 2388 3016 2397
rect 4988 2388 5040 2440
rect 5264 2431 5316 2440
rect 5264 2397 5273 2431
rect 5273 2397 5307 2431
rect 5307 2397 5316 2431
rect 5264 2388 5316 2397
rect 8024 2388 8076 2440
rect 8576 2431 8628 2440
rect 8576 2397 8585 2431
rect 8585 2397 8619 2431
rect 8619 2397 8628 2431
rect 8576 2388 8628 2397
rect 9036 2388 9088 2440
rect 7656 2320 7708 2372
rect 6828 2252 6880 2304
rect 6954 2150 7006 2202
rect 7018 2150 7070 2202
rect 7082 2150 7134 2202
rect 6828 2048 6880 2100
rect 7656 2048 7708 2100
rect 5172 2023 5224 2032
rect 5172 1989 5181 2023
rect 5181 1989 5215 2023
rect 5215 1989 5224 2023
rect 5172 1980 5224 1989
rect 6460 1980 6512 2032
rect 4896 1955 4948 1964
rect 4896 1921 4905 1955
rect 4905 1921 4939 1955
rect 4939 1921 4948 1955
rect 4896 1912 4948 1921
rect 6276 1912 6328 1964
rect 9036 1980 9088 2032
rect 8576 1912 8628 1964
rect 9588 1844 9640 1896
rect 8300 1776 8352 1828
rect 5724 1708 5776 1760
rect 6554 1606 6606 1658
rect 6618 1606 6670 1658
rect 6682 1606 6734 1658
rect 2964 1504 3016 1556
rect 9128 1368 9180 1420
rect 7656 1300 7708 1352
rect 9036 1343 9088 1352
rect 9036 1309 9045 1343
rect 9045 1309 9079 1343
rect 9079 1309 9088 1343
rect 9036 1300 9088 1309
rect 6954 1062 7006 1114
rect 7018 1062 7070 1114
rect 7082 1062 7134 1114
<< metal2 >>
rect 5078 14498 5134 15000
rect 4816 14470 5134 14498
rect 3240 14272 3292 14278
rect 3240 14214 3292 14220
rect 940 13728 992 13734
rect 940 13670 992 13676
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 952 13326 980 13670
rect 940 13320 992 13326
rect 940 13262 992 13268
rect 1124 13184 1176 13190
rect 1124 13126 1176 13132
rect 1400 13184 1452 13190
rect 1400 13126 1452 13132
rect 1584 13184 1636 13190
rect 1584 13126 1636 13132
rect 940 12844 992 12850
rect 940 12786 992 12792
rect 952 11898 980 12786
rect 940 11892 992 11898
rect 940 11834 992 11840
rect 478 11792 534 11801
rect 478 11727 534 11736
rect 492 10742 520 11727
rect 1032 11076 1084 11082
rect 1032 11018 1084 11024
rect 1044 10985 1072 11018
rect 1030 10976 1086 10985
rect 1030 10911 1086 10920
rect 480 10736 532 10742
rect 480 10678 532 10684
rect 478 10160 534 10169
rect 478 10095 480 10104
rect 532 10095 534 10104
rect 480 10066 532 10072
rect 386 9344 442 9353
rect 386 9279 442 9288
rect 400 8906 428 9279
rect 388 8900 440 8906
rect 1136 8888 1164 13126
rect 1412 12889 1440 13126
rect 1398 12880 1454 12889
rect 1216 12844 1268 12850
rect 1398 12815 1454 12824
rect 1216 12786 1268 12792
rect 1228 12442 1256 12786
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1492 12776 1544 12782
rect 1492 12718 1544 12724
rect 1412 12617 1440 12718
rect 1398 12608 1454 12617
rect 1398 12543 1454 12552
rect 1504 12442 1532 12718
rect 1216 12436 1268 12442
rect 1216 12378 1268 12384
rect 1492 12436 1544 12442
rect 1492 12378 1544 12384
rect 1400 12232 1452 12238
rect 1400 12174 1452 12180
rect 1412 11218 1440 12174
rect 1596 12050 1624 13126
rect 1688 12434 1716 13670
rect 2544 13626 2744 14192
rect 2544 13574 2554 13626
rect 2606 13574 2618 13626
rect 2670 13574 2682 13626
rect 2734 13574 2744 13626
rect 1860 13524 1912 13530
rect 1860 13466 1912 13472
rect 1872 13326 1900 13466
rect 1860 13320 1912 13326
rect 1860 13262 1912 13268
rect 2412 13320 2464 13326
rect 2412 13262 2464 13268
rect 2044 13184 2096 13190
rect 2044 13126 2096 13132
rect 1688 12406 1900 12434
rect 1504 12022 1624 12050
rect 1400 11212 1452 11218
rect 1400 11154 1452 11160
rect 1412 10742 1440 11154
rect 1400 10736 1452 10742
rect 1400 10678 1452 10684
rect 1504 9466 1532 12022
rect 1676 11892 1728 11898
rect 1676 11834 1728 11840
rect 1688 11082 1716 11834
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1688 10606 1716 11018
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1676 10600 1728 10606
rect 1676 10542 1728 10548
rect 1688 9722 1716 10542
rect 1676 9716 1728 9722
rect 1676 9658 1728 9664
rect 1676 9512 1728 9518
rect 1504 9438 1624 9466
rect 1676 9454 1728 9460
rect 1216 8900 1268 8906
rect 1136 8860 1216 8888
rect 388 8842 440 8848
rect 1216 8842 1268 8848
rect 1032 8492 1084 8498
rect 1032 8434 1084 8440
rect 938 7712 994 7721
rect 938 7647 994 7656
rect 952 7410 980 7647
rect 940 7404 992 7410
rect 940 7346 992 7352
rect 480 6316 532 6322
rect 480 6258 532 6264
rect 492 6089 520 6258
rect 478 6080 534 6089
rect 478 6015 534 6024
rect 388 5772 440 5778
rect 388 5714 440 5720
rect 400 5273 428 5714
rect 386 5264 442 5273
rect 386 5199 442 5208
rect 940 5160 992 5166
rect 940 5102 992 5108
rect 388 4616 440 4622
rect 388 4558 440 4564
rect 400 4457 428 4558
rect 386 4448 442 4457
rect 386 4383 442 4392
rect 952 4146 980 5102
rect 940 4140 992 4146
rect 940 4082 992 4088
rect 952 2825 980 4082
rect 1044 3641 1072 8434
rect 1124 7812 1176 7818
rect 1124 7754 1176 7760
rect 1136 6458 1164 7754
rect 1308 7744 1360 7750
rect 1308 7686 1360 7692
rect 1320 7562 1348 7686
rect 1320 7546 1440 7562
rect 1320 7540 1452 7546
rect 1320 7534 1400 7540
rect 1400 7482 1452 7488
rect 1216 7404 1268 7410
rect 1216 7346 1268 7352
rect 1228 6905 1256 7346
rect 1214 6896 1270 6905
rect 1214 6831 1270 6840
rect 1124 6452 1176 6458
rect 1124 6394 1176 6400
rect 1124 5704 1176 5710
rect 1124 5646 1176 5652
rect 1136 4486 1164 5646
rect 1216 5160 1268 5166
rect 1216 5102 1268 5108
rect 1228 4826 1256 5102
rect 1216 4820 1268 4826
rect 1216 4762 1268 4768
rect 1124 4480 1176 4486
rect 1124 4422 1176 4428
rect 1030 3632 1086 3641
rect 1030 3567 1086 3576
rect 1596 3233 1624 9438
rect 1688 8498 1716 9454
rect 1780 8634 1808 10678
rect 1872 9382 1900 12406
rect 2056 10826 2084 13126
rect 2424 12434 2452 13262
rect 2240 12406 2452 12434
rect 2544 13156 2744 13574
rect 2944 14170 3144 14192
rect 2944 14118 2954 14170
rect 3006 14118 3018 14170
rect 3070 14118 3082 14170
rect 3134 14118 3144 14170
rect 2944 13556 3144 14118
rect 3252 13938 3280 14214
rect 3344 13956 3544 14192
rect 3240 13932 3292 13938
rect 3240 13874 3292 13880
rect 3344 13900 3376 13956
rect 3432 13900 3456 13956
rect 3512 13900 3544 13956
rect 3344 13876 3544 13900
rect 2944 13500 2976 13556
rect 3032 13500 3056 13556
rect 3112 13500 3144 13556
rect 2944 13476 3144 13500
rect 2944 13420 2976 13476
rect 3032 13420 3056 13476
rect 3112 13420 3144 13476
rect 2544 13100 2576 13156
rect 2632 13100 2656 13156
rect 2712 13100 2744 13156
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2544 13076 2744 13100
rect 2544 13020 2576 13076
rect 2632 13020 2656 13076
rect 2712 13020 2744 13076
rect 2544 12538 2744 13020
rect 2544 12486 2554 12538
rect 2606 12486 2618 12538
rect 2670 12486 2682 12538
rect 2734 12486 2744 12538
rect 2134 11248 2190 11257
rect 2134 11183 2190 11192
rect 2148 11150 2176 11183
rect 2240 11150 2268 12406
rect 2412 12300 2464 12306
rect 2412 12242 2464 12248
rect 2318 12200 2374 12209
rect 2318 12135 2320 12144
rect 2372 12135 2374 12144
rect 2320 12106 2372 12112
rect 2332 11830 2360 12106
rect 2424 11898 2452 12242
rect 2412 11892 2464 11898
rect 2412 11834 2464 11840
rect 2320 11824 2372 11830
rect 2320 11766 2372 11772
rect 2412 11688 2464 11694
rect 2412 11630 2464 11636
rect 2320 11552 2372 11558
rect 2320 11494 2372 11500
rect 2136 11144 2188 11150
rect 2136 11086 2188 11092
rect 2228 11144 2280 11150
rect 2228 11086 2280 11092
rect 2056 10798 2176 10826
rect 2044 10464 2096 10470
rect 2044 10406 2096 10412
rect 2056 10266 2084 10406
rect 2044 10260 2096 10266
rect 2044 10202 2096 10208
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1860 9376 1912 9382
rect 1860 9318 1912 9324
rect 1768 8628 1820 8634
rect 1768 8570 1820 8576
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 7342 1716 8434
rect 1676 7336 1728 7342
rect 1676 7278 1728 7284
rect 1964 4554 1992 9930
rect 2056 9654 2084 10202
rect 2044 9648 2096 9654
rect 2044 9590 2096 9596
rect 2056 9110 2084 9590
rect 2148 9178 2176 10798
rect 2228 10600 2280 10606
rect 2228 10542 2280 10548
rect 2240 10266 2268 10542
rect 2228 10260 2280 10266
rect 2228 10202 2280 10208
rect 2228 10056 2280 10062
rect 2228 9998 2280 10004
rect 2136 9172 2188 9178
rect 2136 9114 2188 9120
rect 2044 9104 2096 9110
rect 2044 9046 2096 9052
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 2044 8900 2096 8906
rect 2044 8842 2096 8848
rect 2056 8673 2084 8842
rect 2042 8664 2098 8673
rect 2042 8599 2098 8608
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 2056 7274 2084 8230
rect 2044 7268 2096 7274
rect 2044 7210 2096 7216
rect 1952 4548 2004 4554
rect 1952 4490 2004 4496
rect 1582 3224 1638 3233
rect 1582 3159 1638 3168
rect 938 2816 994 2825
rect 938 2751 994 2760
rect 1964 2553 1992 4490
rect 2148 2650 2176 8910
rect 2240 8294 2268 9998
rect 2332 9518 2360 11494
rect 2424 11393 2452 11630
rect 2544 11450 2744 12486
rect 2792 12442 2820 13126
rect 2944 13082 3144 13420
rect 3344 13820 3376 13876
rect 3432 13820 3456 13876
rect 3512 13820 3544 13876
rect 3240 13320 3292 13326
rect 3240 13262 3292 13268
rect 2944 13030 2954 13082
rect 3006 13030 3018 13082
rect 3070 13030 3082 13082
rect 3134 13030 3144 13082
rect 2780 12436 2832 12442
rect 2780 12378 2832 12384
rect 2780 12164 2832 12170
rect 2780 12106 2832 12112
rect 2544 11398 2554 11450
rect 2606 11398 2618 11450
rect 2670 11398 2682 11450
rect 2734 11398 2744 11450
rect 2410 11384 2466 11393
rect 2410 11319 2466 11328
rect 2412 11280 2464 11286
rect 2412 11222 2464 11228
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2424 8922 2452 11222
rect 2332 8894 2452 8922
rect 2544 10362 2744 11398
rect 2792 11354 2820 12106
rect 2944 11994 3144 13030
rect 3252 12986 3280 13262
rect 3240 12980 3292 12986
rect 3240 12922 3292 12928
rect 3240 12708 3292 12714
rect 3240 12650 3292 12656
rect 2944 11942 2954 11994
rect 3006 11942 3018 11994
rect 3070 11942 3082 11994
rect 3134 11942 3144 11994
rect 2780 11348 2832 11354
rect 2780 11290 2832 11296
rect 2544 10310 2554 10362
rect 2606 10310 2618 10362
rect 2670 10310 2682 10362
rect 2734 10310 2744 10362
rect 2544 9274 2744 10310
rect 2944 10906 3144 11942
rect 3252 11898 3280 12650
rect 3240 11892 3292 11898
rect 3240 11834 3292 11840
rect 3240 11552 3292 11558
rect 3240 11494 3292 11500
rect 2944 10854 2954 10906
rect 3006 10854 3018 10906
rect 3070 10854 3082 10906
rect 3134 10854 3144 10906
rect 2780 10056 2832 10062
rect 2780 9998 2832 10004
rect 2792 9450 2820 9998
rect 2944 9818 3144 10854
rect 2944 9766 2954 9818
rect 3006 9766 3018 9818
rect 3070 9766 3082 9818
rect 3134 9766 3144 9818
rect 2944 9556 3144 9766
rect 3252 9586 3280 11494
rect 3344 9956 3544 13820
rect 3606 12200 3662 12209
rect 3606 12135 3662 12144
rect 3620 12102 3648 12135
rect 3608 12096 3660 12102
rect 3608 12038 3660 12044
rect 3608 10600 3660 10606
rect 3608 10542 3660 10548
rect 3620 10266 3648 10542
rect 3744 10356 3944 14192
rect 4816 14006 4844 14470
rect 5078 14400 5134 14470
rect 5354 14400 5410 15000
rect 5630 14498 5686 15000
rect 5906 14498 5962 15000
rect 6182 14498 6238 15000
rect 6458 14498 6514 15000
rect 6734 14498 6790 15000
rect 7010 14498 7066 15000
rect 7286 14498 7342 15000
rect 7562 14498 7618 15000
rect 7838 14498 7894 15000
rect 8114 14498 8170 15000
rect 8390 14498 8446 15000
rect 5552 14470 5686 14498
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 4804 14000 4856 14006
rect 4804 13942 4856 13948
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 3976 13796 4028 13802
rect 3976 13738 4028 13744
rect 3988 10690 4016 13738
rect 4068 13184 4120 13190
rect 4068 13126 4120 13132
rect 4080 11558 4108 13126
rect 4160 12912 4212 12918
rect 4160 12854 4212 12860
rect 4172 12374 4200 12854
rect 4160 12368 4212 12374
rect 4160 12310 4212 12316
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4160 12164 4212 12170
rect 4160 12106 4212 12112
rect 4068 11552 4120 11558
rect 4068 11494 4120 11500
rect 4172 11257 4200 12106
rect 4158 11248 4214 11257
rect 4068 11212 4120 11218
rect 4158 11183 4214 11192
rect 4068 11154 4120 11160
rect 4080 10810 4108 11154
rect 4068 10804 4120 10810
rect 4068 10746 4120 10752
rect 3988 10662 4108 10690
rect 3744 10300 3776 10356
rect 3832 10300 3856 10356
rect 3912 10300 3944 10356
rect 3744 10276 3944 10300
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3744 10220 3776 10276
rect 3832 10220 3856 10276
rect 3912 10220 3944 10276
rect 3344 9900 3376 9956
rect 3432 9900 3456 9956
rect 3512 9900 3544 9956
rect 3344 9876 3544 9900
rect 3344 9820 3376 9876
rect 3432 9820 3456 9876
rect 3512 9820 3544 9876
rect 2944 9500 2976 9556
rect 3032 9500 3056 9556
rect 3112 9500 3144 9556
rect 3240 9580 3292 9586
rect 3240 9522 3292 9528
rect 2944 9476 3144 9500
rect 2780 9444 2832 9450
rect 2780 9386 2832 9392
rect 2944 9420 2976 9476
rect 3032 9420 3056 9476
rect 3112 9420 3144 9476
rect 2544 9222 2554 9274
rect 2606 9222 2618 9274
rect 2670 9222 2682 9274
rect 2734 9222 2744 9274
rect 2544 9156 2744 9222
rect 2544 9100 2576 9156
rect 2632 9100 2656 9156
rect 2712 9100 2744 9156
rect 2544 9076 2744 9100
rect 2544 9020 2576 9076
rect 2632 9020 2656 9076
rect 2712 9020 2744 9076
rect 2780 9104 2832 9110
rect 2780 9046 2832 9052
rect 2228 8288 2280 8294
rect 2228 8230 2280 8236
rect 2332 7750 2360 8894
rect 2412 8832 2464 8838
rect 2412 8774 2464 8780
rect 2424 8566 2452 8774
rect 2412 8560 2464 8566
rect 2412 8502 2464 8508
rect 2544 8186 2744 9020
rect 2544 8134 2554 8186
rect 2606 8134 2618 8186
rect 2670 8134 2682 8186
rect 2734 8134 2744 8186
rect 2228 7744 2280 7750
rect 2228 7686 2280 7692
rect 2320 7744 2372 7750
rect 2320 7686 2372 7692
rect 2240 7478 2268 7686
rect 2228 7472 2280 7478
rect 2228 7414 2280 7420
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 2320 7268 2372 7274
rect 2320 7210 2372 7216
rect 2332 5234 2360 7210
rect 2320 5228 2372 5234
rect 2320 5170 2372 5176
rect 2332 4758 2360 5170
rect 2424 5166 2452 7278
rect 2544 7098 2744 8134
rect 2792 7886 2820 9046
rect 2944 8730 3144 9420
rect 3240 8968 3292 8974
rect 3240 8910 3292 8916
rect 3252 8809 3280 8910
rect 3238 8800 3294 8809
rect 3238 8735 3294 8744
rect 2944 8678 2954 8730
rect 3006 8678 3018 8730
rect 3070 8678 3082 8730
rect 3134 8678 3144 8730
rect 2780 7880 2832 7886
rect 2780 7822 2832 7828
rect 2544 7046 2554 7098
rect 2606 7046 2618 7098
rect 2670 7046 2682 7098
rect 2734 7046 2744 7098
rect 2544 6010 2744 7046
rect 2544 5958 2554 6010
rect 2606 5958 2618 6010
rect 2670 5958 2682 6010
rect 2734 5958 2744 6010
rect 2412 5160 2464 5166
rect 2412 5102 2464 5108
rect 2544 5156 2744 5958
rect 2544 5100 2576 5156
rect 2632 5100 2656 5156
rect 2712 5100 2744 5156
rect 2544 5076 2744 5100
rect 2544 5020 2576 5076
rect 2632 5020 2656 5076
rect 2712 5020 2744 5076
rect 2544 4922 2744 5020
rect 2544 4870 2554 4922
rect 2606 4870 2618 4922
rect 2670 4870 2682 4922
rect 2734 4870 2744 4922
rect 2320 4752 2372 4758
rect 2320 4694 2372 4700
rect 2544 4094 2744 4870
rect 2944 7642 3144 8678
rect 3238 8664 3294 8673
rect 3238 8599 3294 8608
rect 3252 8566 3280 8599
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3240 7880 3292 7886
rect 3240 7822 3292 7828
rect 2944 7590 2954 7642
rect 3006 7590 3018 7642
rect 3070 7590 3082 7642
rect 3134 7590 3144 7642
rect 2944 6554 3144 7590
rect 3252 7546 3280 7822
rect 3240 7540 3292 7546
rect 3240 7482 3292 7488
rect 2944 6502 2954 6554
rect 3006 6502 3018 6554
rect 3070 6502 3082 6554
rect 3134 6502 3144 6554
rect 2944 5556 3144 6502
rect 2944 5500 2976 5556
rect 3032 5500 3056 5556
rect 3112 5500 3144 5556
rect 2944 5476 3144 5500
rect 2944 5466 2976 5476
rect 3032 5466 3056 5476
rect 3112 5466 3144 5476
rect 2944 5414 2954 5466
rect 3006 5414 3018 5420
rect 3070 5414 3082 5420
rect 3134 5414 3144 5466
rect 2780 4616 2832 4622
rect 2780 4558 2832 4564
rect 2792 2774 2820 4558
rect 2944 4378 3144 5414
rect 2944 4326 2954 4378
rect 3006 4326 3018 4378
rect 3070 4326 3082 4378
rect 3134 4326 3144 4378
rect 2944 4094 3144 4326
rect 3344 5956 3544 9820
rect 3608 9716 3660 9722
rect 3608 9658 3660 9664
rect 3620 8498 3648 9658
rect 3608 8492 3660 8498
rect 3608 8434 3660 8440
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3620 7954 3648 8230
rect 3608 7948 3660 7954
rect 3608 7890 3660 7896
rect 3744 6356 3944 10220
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 9042 4016 9454
rect 4080 9110 4108 10662
rect 4160 10668 4212 10674
rect 4160 10610 4212 10616
rect 4172 9994 4200 10610
rect 4160 9988 4212 9994
rect 4160 9930 4212 9936
rect 4172 9722 4200 9930
rect 4160 9716 4212 9722
rect 4160 9658 4212 9664
rect 4264 9466 4292 12174
rect 4344 10464 4396 10470
rect 4344 10406 4396 10412
rect 4356 9654 4384 10406
rect 4344 9648 4396 9654
rect 4344 9590 4396 9596
rect 4264 9438 4384 9466
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4068 9104 4120 9110
rect 4068 9046 4120 9052
rect 3976 9036 4028 9042
rect 3976 8978 4028 8984
rect 4264 8922 4292 9318
rect 4080 8894 4292 8922
rect 4080 7002 4108 8894
rect 4356 8362 4384 9438
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4448 8090 4476 13874
rect 4896 13728 4948 13734
rect 4896 13670 4948 13676
rect 4528 13320 4580 13326
rect 4528 13262 4580 13268
rect 4540 12850 4568 13262
rect 4528 12844 4580 12850
rect 4528 12786 4580 12792
rect 4620 12232 4672 12238
rect 4620 12174 4672 12180
rect 4528 12096 4580 12102
rect 4528 12038 4580 12044
rect 4540 11830 4568 12038
rect 4528 11824 4580 11830
rect 4528 11766 4580 11772
rect 4540 10674 4568 11766
rect 4632 11354 4660 12174
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 10668 4580 10674
rect 4528 10610 4580 10616
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4436 8084 4488 8090
rect 4436 8026 4488 8032
rect 4068 6996 4120 7002
rect 4068 6938 4120 6944
rect 3744 6300 3776 6356
rect 3832 6300 3856 6356
rect 3912 6300 3944 6356
rect 3744 6276 3944 6300
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3744 6220 3776 6276
rect 3832 6220 3856 6276
rect 3912 6220 3944 6276
rect 3344 5900 3376 5956
rect 3432 5900 3456 5956
rect 3512 5900 3544 5956
rect 3344 5876 3544 5900
rect 3344 5820 3376 5876
rect 3432 5820 3456 5876
rect 3512 5820 3544 5876
rect 3344 4094 3544 5820
rect 3620 5778 3648 6190
rect 3608 5772 3660 5778
rect 3608 5714 3660 5720
rect 3620 4146 3648 5714
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3620 3602 3648 4082
rect 3608 3596 3660 3602
rect 3608 3538 3660 3544
rect 2792 2746 3004 2774
rect 2136 2644 2188 2650
rect 2136 2586 2188 2592
rect 386 2544 442 2553
rect 386 2479 442 2488
rect 1950 2544 2006 2553
rect 1950 2479 2006 2488
rect 400 2009 428 2479
rect 2976 2446 3004 2746
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 900 2356 1100 2365
rect 900 2300 932 2356
rect 988 2300 1012 2356
rect 1068 2300 1100 2356
rect 900 2276 1100 2300
rect 900 2220 932 2276
rect 988 2220 1012 2276
rect 1068 2220 1100 2276
rect 900 2211 1100 2220
rect 386 2000 442 2009
rect 386 1935 442 1944
rect 1500 1956 1700 1965
rect 1500 1900 1532 1956
rect 1588 1900 1612 1956
rect 1668 1900 1700 1956
rect 1500 1876 1700 1900
rect 1500 1820 1532 1876
rect 1588 1820 1612 1876
rect 1668 1820 1700 1876
rect 1500 1811 1700 1820
rect 2976 1562 3004 2382
rect 3744 2356 3944 6220
rect 4160 5160 4212 5166
rect 4160 5102 4212 5108
rect 4172 3738 4200 5102
rect 4632 4826 4660 9454
rect 4724 7478 4752 11494
rect 4908 9382 4936 13670
rect 5368 13394 5396 14282
rect 5356 13388 5408 13394
rect 5356 13330 5408 13336
rect 5080 13252 5132 13258
rect 5080 13194 5132 13200
rect 5092 12850 5120 13194
rect 5080 12844 5132 12850
rect 5080 12786 5132 12792
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 5092 11558 5120 12174
rect 5552 12102 5580 14470
rect 5630 14400 5686 14470
rect 5736 14470 5962 14498
rect 5632 13796 5684 13802
rect 5632 13738 5684 13744
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5080 11552 5132 11558
rect 5080 11494 5132 11500
rect 5356 11144 5408 11150
rect 5356 11086 5408 11092
rect 5172 11076 5224 11082
rect 5172 11018 5224 11024
rect 4988 10464 5040 10470
rect 4988 10406 5040 10412
rect 4896 9376 4948 9382
rect 4896 9318 4948 9324
rect 4896 9036 4948 9042
rect 4896 8978 4948 8984
rect 4804 7744 4856 7750
rect 4804 7686 4856 7692
rect 4712 7472 4764 7478
rect 4712 7414 4764 7420
rect 4816 6798 4844 7686
rect 4908 7410 4936 8978
rect 5000 8974 5028 10406
rect 5184 10198 5212 11018
rect 5368 10810 5396 11086
rect 5356 10804 5408 10810
rect 5356 10746 5408 10752
rect 5644 10742 5672 13738
rect 5736 13530 5764 14470
rect 5906 14400 5962 14470
rect 6012 14470 6238 14498
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5724 13524 5776 13530
rect 5724 13466 5776 13472
rect 5920 13462 5948 13670
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 6012 13308 6040 14470
rect 6182 14400 6238 14470
rect 6288 14470 6514 14498
rect 6288 14090 6316 14470
rect 6458 14400 6514 14470
rect 6564 14470 6790 14498
rect 6564 14362 6592 14470
rect 6734 14400 6790 14470
rect 6840 14470 7066 14498
rect 5920 13280 6040 13308
rect 6104 14062 6316 14090
rect 6472 14334 6592 14362
rect 5816 12640 5868 12646
rect 5816 12582 5868 12588
rect 5632 10736 5684 10742
rect 5632 10678 5684 10684
rect 5356 10668 5408 10674
rect 5356 10610 5408 10616
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5172 10192 5224 10198
rect 5172 10134 5224 10140
rect 5080 10056 5132 10062
rect 5080 9998 5132 10004
rect 5092 9042 5120 9998
rect 5172 9988 5224 9994
rect 5172 9930 5224 9936
rect 5184 9110 5212 9930
rect 5368 9586 5396 10610
rect 5552 10554 5580 10610
rect 5460 10526 5580 10554
rect 5356 9580 5408 9586
rect 5356 9522 5408 9528
rect 5172 9104 5224 9110
rect 5172 9046 5224 9052
rect 5080 9036 5132 9042
rect 5080 8978 5132 8984
rect 5368 8974 5396 9522
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5356 8968 5408 8974
rect 5356 8910 5408 8916
rect 5172 8900 5224 8906
rect 5172 8842 5224 8848
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5092 7410 5120 8570
rect 4896 7404 4948 7410
rect 4896 7346 4948 7352
rect 5080 7404 5132 7410
rect 5080 7346 5132 7352
rect 4804 6792 4856 6798
rect 4804 6734 4856 6740
rect 4816 6254 4844 6734
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4908 5794 4936 7346
rect 5092 6866 5120 7346
rect 5080 6860 5132 6866
rect 5080 6802 5132 6808
rect 5092 6458 5120 6802
rect 5080 6452 5132 6458
rect 5080 6394 5132 6400
rect 4816 5778 4936 5794
rect 4804 5772 4936 5778
rect 4856 5766 4936 5772
rect 4804 5714 4856 5720
rect 5184 5574 5212 8842
rect 5460 7274 5488 10526
rect 5644 10198 5672 10678
rect 5724 10600 5776 10606
rect 5724 10542 5776 10548
rect 5736 10266 5764 10542
rect 5724 10260 5776 10266
rect 5724 10202 5776 10208
rect 5632 10192 5684 10198
rect 5632 10134 5684 10140
rect 5540 10056 5592 10062
rect 5540 9998 5592 10004
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5552 9654 5580 9998
rect 5540 9648 5592 9654
rect 5540 9590 5592 9596
rect 5644 8634 5672 9998
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5736 7818 5764 8570
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5724 7812 5776 7818
rect 5724 7754 5776 7760
rect 5644 7410 5672 7754
rect 5736 7410 5764 7754
rect 5632 7404 5684 7410
rect 5632 7346 5684 7352
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 5540 7200 5592 7206
rect 5540 7142 5592 7148
rect 5552 6730 5580 7142
rect 5540 6724 5592 6730
rect 5540 6666 5592 6672
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5264 6316 5316 6322
rect 5264 6258 5316 6264
rect 5172 5568 5224 5574
rect 5172 5510 5224 5516
rect 4620 4820 4672 4826
rect 4620 4762 4672 4768
rect 5276 4622 5304 6258
rect 5264 4616 5316 4622
rect 5264 4558 5316 4564
rect 5276 4214 5304 4558
rect 5356 4480 5408 4486
rect 5356 4422 5408 4428
rect 5368 4214 5396 4422
rect 5264 4208 5316 4214
rect 5264 4154 5316 4156
rect 5092 4150 5316 4154
rect 5356 4208 5408 4214
rect 5356 4150 5408 4156
rect 5092 4126 5304 4150
rect 4160 3732 4212 3738
rect 4160 3674 4212 3680
rect 4988 3732 5040 3738
rect 4988 3674 5040 3680
rect 4896 3596 4948 3602
rect 4896 3538 4948 3544
rect 3744 2300 3776 2356
rect 3832 2300 3856 2356
rect 3912 2300 3944 2356
rect 3744 2276 3944 2300
rect 3744 2220 3776 2276
rect 3832 2220 3856 2276
rect 3912 2220 3944 2276
rect 2964 1556 3016 1562
rect 2964 1498 3016 1504
rect 3744 1040 3944 2220
rect 4908 1970 4936 3538
rect 5000 2446 5028 3674
rect 5092 3398 5120 4126
rect 5368 4026 5396 4150
rect 5460 4146 5488 6394
rect 5736 6118 5764 7346
rect 5724 6112 5776 6118
rect 5724 6054 5776 6060
rect 5828 5302 5856 12582
rect 5920 10198 5948 13280
rect 6104 13138 6132 14062
rect 6276 13932 6328 13938
rect 6276 13874 6328 13880
rect 6184 13524 6236 13530
rect 6184 13466 6236 13472
rect 6012 13110 6132 13138
rect 6012 12442 6040 13110
rect 6092 12640 6144 12646
rect 6092 12582 6144 12588
rect 6000 12436 6052 12442
rect 6000 12378 6052 12384
rect 6104 12170 6132 12582
rect 6196 12322 6224 13466
rect 6288 12442 6316 13874
rect 6472 13870 6500 14334
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6544 13626 6744 14192
rect 6840 14074 6868 14470
rect 7010 14400 7066 14470
rect 7116 14470 7342 14498
rect 7116 14346 7144 14470
rect 7286 14400 7342 14470
rect 7392 14470 7618 14498
rect 7392 14362 7420 14470
rect 7562 14400 7618 14470
rect 7668 14470 7894 14498
rect 7668 14362 7696 14470
rect 7838 14400 7894 14470
rect 8036 14470 8170 14498
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7208 14334 7420 14362
rect 7576 14334 7696 14362
rect 6944 14170 7144 14192
rect 6944 14118 6954 14170
rect 7006 14118 7018 14170
rect 7070 14118 7082 14170
rect 7134 14118 7144 14170
rect 6828 14068 6880 14074
rect 6828 14010 6880 14016
rect 6544 13574 6554 13626
rect 6606 13574 6618 13626
rect 6670 13574 6682 13626
rect 6734 13574 6744 13626
rect 6460 13320 6512 13326
rect 6460 13262 6512 13268
rect 6368 13252 6420 13258
rect 6368 13194 6420 13200
rect 6380 12918 6408 13194
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6472 12442 6500 13262
rect 6544 13156 6744 13574
rect 6544 13100 6576 13156
rect 6632 13100 6656 13156
rect 6712 13100 6744 13156
rect 6544 13076 6744 13100
rect 6544 13020 6576 13076
rect 6632 13020 6656 13076
rect 6712 13020 6744 13076
rect 6544 12538 6744 13020
rect 6944 13556 7144 14118
rect 7208 13734 7236 14334
rect 7344 13956 7544 14192
rect 7344 13900 7376 13956
rect 7432 13900 7456 13956
rect 7512 13900 7544 13956
rect 7344 13876 7544 13900
rect 7344 13820 7376 13876
rect 7432 13820 7456 13876
rect 7512 13820 7544 13876
rect 7196 13728 7248 13734
rect 7196 13670 7248 13676
rect 6944 13500 6976 13556
rect 7032 13500 7056 13556
rect 7112 13500 7144 13556
rect 6944 13476 7144 13500
rect 6944 13420 6976 13476
rect 7032 13420 7056 13476
rect 7112 13420 7144 13476
rect 6944 13082 7144 13420
rect 6944 13030 6954 13082
rect 7006 13030 7018 13082
rect 7070 13030 7082 13082
rect 7134 13030 7144 13082
rect 6828 12776 6880 12782
rect 6828 12718 6880 12724
rect 6544 12486 6554 12538
rect 6606 12486 6618 12538
rect 6670 12486 6682 12538
rect 6734 12486 6744 12538
rect 6276 12436 6328 12442
rect 6276 12378 6328 12384
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6196 12294 6316 12322
rect 6288 12238 6316 12294
rect 6276 12232 6328 12238
rect 6276 12174 6328 12180
rect 6092 12164 6144 12170
rect 6092 12106 6144 12112
rect 6368 12164 6420 12170
rect 6368 12106 6420 12112
rect 6380 11762 6408 12106
rect 6000 11756 6052 11762
rect 6000 11698 6052 11704
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6012 11626 6040 11698
rect 6092 11688 6144 11694
rect 6092 11630 6144 11636
rect 6460 11688 6512 11694
rect 6460 11630 6512 11636
rect 6000 11620 6052 11626
rect 6000 11562 6052 11568
rect 6012 10742 6040 11562
rect 6104 11054 6132 11630
rect 6274 11384 6330 11393
rect 6274 11319 6330 11328
rect 6288 11150 6316 11319
rect 6276 11144 6328 11150
rect 6276 11086 6328 11092
rect 6104 11026 6224 11054
rect 6000 10736 6052 10742
rect 6000 10678 6052 10684
rect 6196 10674 6224 11026
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6184 10532 6236 10538
rect 6184 10474 6236 10480
rect 5908 10192 5960 10198
rect 5908 10134 5960 10140
rect 6000 10056 6052 10062
rect 6000 9998 6052 10004
rect 5908 8560 5960 8566
rect 5908 8502 5960 8508
rect 5920 8022 5948 8502
rect 5908 8016 5960 8022
rect 5908 7958 5960 7964
rect 5908 7268 5960 7274
rect 5908 7210 5960 7216
rect 5920 6322 5948 7210
rect 5908 6316 5960 6322
rect 5908 6258 5960 6264
rect 5816 5296 5868 5302
rect 5816 5238 5868 5244
rect 5920 5114 5948 6258
rect 6012 5370 6040 9998
rect 6196 8906 6224 10474
rect 6288 9722 6316 11086
rect 6472 10062 6500 11630
rect 6544 11450 6744 12486
rect 6544 11398 6554 11450
rect 6606 11398 6618 11450
rect 6670 11398 6682 11450
rect 6734 11398 6744 11450
rect 6544 10362 6744 11398
rect 6544 10310 6554 10362
rect 6606 10310 6618 10362
rect 6670 10310 6682 10362
rect 6734 10310 6744 10362
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6276 9716 6328 9722
rect 6276 9658 6328 9664
rect 6380 9586 6408 9930
rect 6460 9920 6512 9926
rect 6460 9862 6512 9868
rect 6368 9580 6420 9586
rect 6368 9522 6420 9528
rect 6472 9518 6500 9862
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6544 9274 6744 10310
rect 6544 9222 6554 9274
rect 6606 9222 6618 9274
rect 6670 9222 6682 9274
rect 6734 9222 6744 9274
rect 6368 9172 6420 9178
rect 6368 9114 6420 9120
rect 6460 9172 6512 9178
rect 6460 9114 6512 9120
rect 6544 9156 6744 9222
rect 6840 9178 6868 12718
rect 6944 11994 7144 13030
rect 7196 12776 7248 12782
rect 7196 12718 7248 12724
rect 6944 11942 6954 11994
rect 7006 11942 7018 11994
rect 7070 11942 7082 11994
rect 7134 11942 7144 11994
rect 6944 10906 7144 11942
rect 7208 11354 7236 12718
rect 7196 11348 7248 11354
rect 7196 11290 7248 11296
rect 6944 10854 6954 10906
rect 7006 10854 7018 10906
rect 7070 10854 7082 10906
rect 7134 10854 7144 10906
rect 6944 9818 7144 10854
rect 6944 9766 6954 9818
rect 7006 9766 7018 9818
rect 7070 9766 7082 9818
rect 7134 9766 7144 9818
rect 6944 9556 7144 9766
rect 6944 9500 6976 9556
rect 7032 9500 7056 9556
rect 7112 9500 7144 9556
rect 6944 9476 7144 9500
rect 6944 9420 6976 9476
rect 7032 9420 7056 9476
rect 7112 9420 7144 9476
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 6104 6254 6132 7822
rect 6196 7002 6224 8842
rect 6380 8498 6408 9114
rect 6472 8634 6500 9114
rect 6544 9100 6576 9156
rect 6632 9100 6656 9156
rect 6712 9100 6744 9156
rect 6828 9172 6880 9178
rect 6828 9114 6880 9120
rect 6544 9076 6744 9100
rect 6544 9020 6576 9076
rect 6632 9020 6656 9076
rect 6712 9020 6744 9076
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6368 8492 6420 8498
rect 6368 8434 6420 8440
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6288 7410 6316 7754
rect 6368 7744 6420 7750
rect 6368 7686 6420 7692
rect 6276 7404 6328 7410
rect 6276 7346 6328 7352
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6092 6248 6144 6254
rect 6092 6190 6144 6196
rect 6184 6112 6236 6118
rect 6184 6054 6236 6060
rect 6196 5710 6224 6054
rect 6288 5778 6316 7346
rect 6380 6798 6408 7686
rect 6368 6792 6420 6798
rect 6368 6734 6420 6740
rect 6472 5914 6500 8366
rect 6544 8186 6744 9020
rect 6828 8832 6880 8838
rect 6828 8774 6880 8780
rect 6544 8134 6554 8186
rect 6606 8134 6618 8186
rect 6670 8134 6682 8186
rect 6734 8134 6744 8186
rect 6544 7098 6744 8134
rect 6840 7478 6868 8774
rect 6944 8730 7144 9420
rect 7344 9956 7544 13820
rect 7576 13546 7604 14334
rect 8036 14278 8064 14470
rect 8114 14400 8170 14470
rect 8312 14470 8446 14498
rect 8024 14272 8076 14278
rect 8024 14214 8076 14220
rect 7576 13518 7696 13546
rect 7668 13462 7696 13518
rect 7656 13456 7708 13462
rect 7656 13398 7708 13404
rect 7656 13320 7708 13326
rect 7344 9900 7376 9956
rect 7432 9900 7456 9956
rect 7512 9900 7544 9956
rect 7344 9876 7544 9900
rect 7344 9820 7376 9876
rect 7432 9820 7456 9876
rect 7512 9820 7544 9876
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 8974 7236 9318
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 6944 8678 6954 8730
rect 7006 8678 7018 8730
rect 7070 8678 7082 8730
rect 7134 8678 7144 8730
rect 6944 7642 7144 8678
rect 7208 8498 7236 8910
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 7196 8288 7248 8294
rect 7194 8256 7196 8265
rect 7248 8256 7250 8265
rect 7194 8191 7250 8200
rect 6944 7590 6954 7642
rect 7006 7590 7018 7642
rect 7070 7590 7082 7642
rect 7134 7590 7144 7642
rect 6828 7472 6880 7478
rect 6828 7414 6880 7420
rect 6544 7046 6554 7098
rect 6606 7046 6618 7098
rect 6670 7046 6682 7098
rect 6734 7046 6744 7098
rect 6544 6010 6744 7046
rect 6544 5958 6554 6010
rect 6606 5958 6618 6010
rect 6670 5958 6682 6010
rect 6734 5958 6744 6010
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6368 5840 6420 5846
rect 6368 5782 6420 5788
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6184 5704 6236 5710
rect 6184 5646 6236 5652
rect 6000 5364 6052 5370
rect 6000 5306 6052 5312
rect 5828 5086 5948 5114
rect 5828 4298 5856 5086
rect 6012 4570 6040 5306
rect 6380 5234 6408 5782
rect 6368 5228 6420 5234
rect 6368 5170 6420 5176
rect 6544 5156 6744 5958
rect 6544 5100 6576 5156
rect 6632 5100 6656 5156
rect 6712 5100 6744 5156
rect 6544 5076 6744 5100
rect 6544 5020 6576 5076
rect 6632 5020 6656 5076
rect 6712 5020 6744 5076
rect 6544 4922 6744 5020
rect 6544 4870 6554 4922
rect 6606 4870 6618 4922
rect 6670 4870 6682 4922
rect 6734 4870 6744 4922
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6012 4554 6132 4570
rect 6012 4548 6144 4554
rect 6012 4542 6092 4548
rect 6092 4490 6144 4496
rect 5828 4270 6040 4298
rect 5906 4176 5962 4185
rect 5448 4140 5500 4146
rect 6012 4146 6040 4270
rect 6288 4185 6316 4626
rect 6274 4176 6330 4185
rect 5906 4111 5962 4120
rect 6000 4140 6052 4146
rect 5448 4082 5500 4088
rect 5184 3998 5396 4026
rect 5080 3392 5132 3398
rect 5080 3334 5132 3340
rect 4988 2440 5040 2446
rect 4988 2382 5040 2388
rect 5184 2038 5212 3998
rect 5264 3936 5316 3942
rect 5264 3878 5316 3884
rect 5276 2446 5304 3878
rect 5460 3738 5488 4082
rect 5448 3732 5500 3738
rect 5448 3674 5500 3680
rect 5920 3602 5948 4111
rect 6274 4111 6330 4120
rect 6000 4082 6052 4088
rect 6544 3834 6744 4870
rect 6544 3782 6554 3834
rect 6606 3782 6618 3834
rect 6670 3782 6682 3834
rect 6734 3782 6744 3834
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 5448 3460 5500 3466
rect 5448 3402 5500 3408
rect 6276 3460 6328 3466
rect 6276 3402 6328 3408
rect 5460 2650 5488 3402
rect 5724 3052 5776 3058
rect 5724 2994 5776 3000
rect 5632 2984 5684 2990
rect 5632 2926 5684 2932
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5644 2553 5672 2926
rect 5630 2544 5686 2553
rect 5630 2479 5686 2488
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 5172 2032 5224 2038
rect 5172 1974 5224 1980
rect 4896 1964 4948 1970
rect 4896 1906 4948 1912
rect 5736 1766 5764 2994
rect 6288 1970 6316 3402
rect 6458 3224 6514 3233
rect 6458 3159 6460 3168
rect 6512 3159 6514 3168
rect 6460 3130 6512 3136
rect 6472 2038 6500 3130
rect 6544 2746 6744 3782
rect 6944 6554 7144 7590
rect 7196 7200 7248 7206
rect 7196 7142 7248 7148
rect 6944 6502 6954 6554
rect 7006 6502 7018 6554
rect 7070 6502 7082 6554
rect 7134 6502 7144 6554
rect 6944 5556 7144 6502
rect 7208 6254 7236 7142
rect 7196 6248 7248 6254
rect 7196 6190 7248 6196
rect 6944 5500 6976 5556
rect 7032 5500 7056 5556
rect 7112 5500 7144 5556
rect 6944 5476 7144 5500
rect 6944 5466 6976 5476
rect 7032 5466 7056 5476
rect 7112 5466 7144 5476
rect 6944 5414 6954 5466
rect 7006 5414 7018 5420
rect 7070 5414 7082 5420
rect 7134 5414 7144 5466
rect 6944 4378 7144 5414
rect 6944 4326 6954 4378
rect 7006 4326 7018 4378
rect 7070 4326 7082 4378
rect 7134 4326 7144 4378
rect 6944 3290 7144 4326
rect 7208 4078 7236 6190
rect 7344 5956 7544 9820
rect 7576 13280 7656 13308
rect 7576 8650 7604 13280
rect 7656 13262 7708 13268
rect 7656 12912 7708 12918
rect 7656 12854 7708 12860
rect 7668 11898 7696 12854
rect 7656 11892 7708 11898
rect 7656 11834 7708 11840
rect 7744 10356 7944 14192
rect 8116 13932 8168 13938
rect 8116 13874 8168 13880
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7744 10300 7776 10356
rect 7832 10300 7856 10356
rect 7912 10300 7944 10356
rect 7744 10276 7944 10300
rect 7744 10220 7776 10276
rect 7832 10220 7856 10276
rect 7912 10220 7944 10276
rect 7656 10192 7708 10198
rect 7656 10134 7708 10140
rect 7668 8974 7696 10134
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7576 8622 7696 8650
rect 7668 8566 7696 8622
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7206 7696 8230
rect 7656 7200 7708 7206
rect 7656 7142 7708 7148
rect 7656 6928 7708 6934
rect 7344 5900 7376 5956
rect 7432 5900 7456 5956
rect 7512 5900 7544 5956
rect 7344 5876 7544 5900
rect 7344 5820 7376 5876
rect 7432 5820 7456 5876
rect 7512 5820 7544 5876
rect 7196 4072 7248 4078
rect 7196 4014 7248 4020
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 6944 3238 6954 3290
rect 7006 3238 7018 3290
rect 7070 3238 7082 3290
rect 7134 3238 7144 3290
rect 6828 3120 6880 3126
rect 6828 3062 6880 3068
rect 6544 2694 6554 2746
rect 6606 2694 6618 2746
rect 6670 2694 6682 2746
rect 6734 2694 6744 2746
rect 6460 2032 6512 2038
rect 6460 1974 6512 1980
rect 6276 1964 6328 1970
rect 6276 1906 6328 1912
rect 5724 1760 5776 1766
rect 5724 1702 5776 1708
rect 6544 1658 6744 2694
rect 6840 2650 6868 3062
rect 6828 2644 6880 2650
rect 6828 2586 6880 2592
rect 6828 2304 6880 2310
rect 6828 2246 6880 2252
rect 6840 2106 6868 2246
rect 6944 2202 7144 3238
rect 7208 3058 7236 3538
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6944 2150 6954 2202
rect 7006 2150 7018 2202
rect 7070 2150 7082 2202
rect 7134 2150 7144 2202
rect 6828 2100 6880 2106
rect 6828 2042 6880 2048
rect 6544 1606 6554 1658
rect 6606 1606 6618 1658
rect 6670 1606 6682 1658
rect 6734 1606 6744 1658
rect 6544 1156 6744 1606
rect 6544 1100 6576 1156
rect 6632 1100 6656 1156
rect 6712 1100 6744 1156
rect 6544 1076 6744 1100
rect 6544 1020 6576 1076
rect 6632 1020 6656 1076
rect 6712 1020 6744 1076
rect 6944 1556 7144 2150
rect 6944 1500 6976 1556
rect 7032 1500 7056 1556
rect 7112 1500 7144 1556
rect 6944 1476 7144 1500
rect 6944 1420 6976 1476
rect 7032 1420 7056 1476
rect 7112 1420 7144 1476
rect 6944 1114 7144 1420
rect 6944 1062 6954 1114
rect 7006 1062 7018 1114
rect 7070 1062 7082 1114
rect 7134 1062 7144 1114
rect 6944 1040 7144 1062
rect 7344 1956 7544 5820
rect 7344 1900 7376 1956
rect 7432 1900 7456 1956
rect 7512 1900 7544 1956
rect 7344 1876 7544 1900
rect 7344 1820 7376 1876
rect 7432 1820 7456 1876
rect 7512 1820 7544 1876
rect 7344 1040 7544 1820
rect 7576 6876 7656 6882
rect 7576 6870 7708 6876
rect 7576 6854 7696 6870
rect 7576 1442 7604 6854
rect 7656 6792 7708 6798
rect 7656 6734 7708 6740
rect 7668 3670 7696 6734
rect 7744 6356 7944 10220
rect 8036 10062 8064 12174
rect 8128 11898 8156 13874
rect 8208 13184 8260 13190
rect 8208 13126 8260 13132
rect 8116 11892 8168 11898
rect 8116 11834 8168 11840
rect 8220 11762 8248 13126
rect 8312 12986 8340 14470
rect 8390 14400 8446 14470
rect 8666 14498 8722 15000
rect 8666 14470 8800 14498
rect 8666 14400 8722 14470
rect 8576 13932 8628 13938
rect 8576 13874 8628 13880
rect 8588 13818 8616 13874
rect 8484 13796 8536 13802
rect 8588 13790 8708 13818
rect 8484 13738 8536 13744
rect 8300 12980 8352 12986
rect 8300 12922 8352 12928
rect 8392 12844 8444 12850
rect 8392 12786 8444 12792
rect 8404 12730 8432 12786
rect 8312 12702 8432 12730
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8128 10713 8156 11018
rect 8312 10810 8340 12702
rect 8496 12594 8524 13738
rect 8576 13728 8628 13734
rect 8576 13670 8628 13676
rect 8588 13394 8616 13670
rect 8576 13388 8628 13394
rect 8576 13330 8628 13336
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8404 12566 8524 12594
rect 8404 12345 8432 12566
rect 8482 12472 8538 12481
rect 8482 12407 8538 12416
rect 8390 12336 8446 12345
rect 8390 12271 8446 12280
rect 8496 12186 8524 12407
rect 8404 12158 8524 12186
rect 8404 11098 8432 12158
rect 8484 12096 8536 12102
rect 8484 12038 8536 12044
rect 8496 11830 8524 12038
rect 8484 11824 8536 11830
rect 8484 11766 8536 11772
rect 8588 11529 8616 13194
rect 8680 12646 8708 13790
rect 8668 12640 8720 12646
rect 8666 12608 8668 12617
rect 8720 12608 8722 12617
rect 8666 12543 8722 12552
rect 8772 12434 8800 14470
rect 8942 14400 8998 15000
rect 9218 14498 9274 15000
rect 9048 14470 9274 14498
rect 8852 13728 8904 13734
rect 8852 13670 8904 13676
rect 8864 13530 8892 13670
rect 8852 13524 8904 13530
rect 8852 13466 8904 13472
rect 8852 13320 8904 13326
rect 8852 13262 8904 13268
rect 8864 12889 8892 13262
rect 8850 12880 8906 12889
rect 8850 12815 8906 12824
rect 8680 12406 8800 12434
rect 8574 11520 8630 11529
rect 8574 11455 8630 11464
rect 8404 11070 8616 11098
rect 8484 11008 8536 11014
rect 8484 10950 8536 10956
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8208 10736 8260 10742
rect 8114 10704 8170 10713
rect 8208 10678 8260 10684
rect 8114 10639 8170 10648
rect 8220 10198 8248 10678
rect 8496 10674 8524 10950
rect 8484 10668 8536 10674
rect 8484 10610 8536 10616
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8312 10062 8340 10406
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8300 10056 8352 10062
rect 8300 9998 8352 10004
rect 8036 9042 8064 9998
rect 8484 9648 8536 9654
rect 8484 9590 8536 9596
rect 8208 9580 8260 9586
rect 8208 9522 8260 9528
rect 8116 9376 8168 9382
rect 8116 9318 8168 9324
rect 8024 9036 8076 9042
rect 8024 8978 8076 8984
rect 8128 8922 8156 9318
rect 7744 6300 7776 6356
rect 7832 6300 7856 6356
rect 7912 6300 7944 6356
rect 7744 6276 7944 6300
rect 7744 6220 7776 6276
rect 7832 6220 7856 6276
rect 7912 6220 7944 6276
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7656 3528 7708 3534
rect 7656 3470 7708 3476
rect 7668 3058 7696 3470
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7656 2372 7708 2378
rect 7656 2314 7708 2320
rect 7744 2356 7944 6220
rect 8036 8894 8156 8922
rect 8036 5710 8064 8894
rect 8116 8832 8168 8838
rect 8116 8774 8168 8780
rect 8128 6798 8156 8774
rect 8220 8090 8248 9522
rect 8496 9110 8524 9590
rect 8484 9104 8536 9110
rect 8484 9046 8536 9052
rect 8208 8084 8260 8090
rect 8208 8026 8260 8032
rect 8392 7948 8444 7954
rect 8392 7890 8444 7896
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8312 7546 8340 7822
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8404 7449 8432 7890
rect 8390 7440 8446 7449
rect 8390 7375 8446 7384
rect 8588 7002 8616 11070
rect 8680 10538 8708 12406
rect 8760 12232 8812 12238
rect 8864 12220 8892 12815
rect 8944 12640 8996 12646
rect 8944 12582 8996 12588
rect 8812 12192 8892 12220
rect 8760 12174 8812 12180
rect 8760 11212 8812 11218
rect 8760 11154 8812 11160
rect 8668 10532 8720 10538
rect 8668 10474 8720 10480
rect 8772 10062 8800 11154
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8680 7478 8708 8434
rect 8772 7886 8800 8910
rect 8956 8498 8984 12582
rect 9048 11558 9076 14470
rect 9218 14400 9274 14470
rect 9588 14000 9640 14006
rect 9586 13968 9588 13977
rect 9640 13968 9642 13977
rect 9586 13903 9642 13912
rect 9588 13456 9640 13462
rect 9588 13398 9640 13404
rect 9128 13252 9180 13258
rect 9128 13194 9180 13200
rect 9140 12238 9168 13194
rect 9600 13161 9628 13398
rect 9586 13152 9642 13161
rect 9586 13087 9642 13096
rect 9128 12232 9180 12238
rect 9128 12174 9180 12180
rect 9036 11552 9088 11558
rect 9036 11494 9088 11500
rect 9140 11082 9168 12174
rect 9128 11076 9180 11082
rect 9128 11018 9180 11024
rect 9140 10062 9168 11018
rect 9588 10124 9640 10130
rect 9588 10066 9640 10072
rect 9128 10056 9180 10062
rect 9128 9998 9180 10004
rect 9140 9722 9168 9998
rect 9600 9897 9628 10066
rect 9586 9888 9642 9897
rect 9586 9823 9642 9832
rect 9128 9716 9180 9722
rect 9128 9658 9180 9664
rect 9140 8974 9168 9658
rect 9586 9072 9642 9081
rect 9586 9007 9642 9016
rect 9128 8968 9180 8974
rect 9128 8910 9180 8916
rect 8944 8492 8996 8498
rect 8944 8434 8996 8440
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 9140 7818 9168 8910
rect 9600 8430 9628 9007
rect 9588 8424 9640 8430
rect 9588 8366 9640 8372
rect 9128 7812 9180 7818
rect 9128 7754 9180 7760
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8576 6996 8628 7002
rect 8576 6938 8628 6944
rect 8956 6798 8984 7346
rect 8116 6792 8168 6798
rect 8116 6734 8168 6740
rect 8576 6792 8628 6798
rect 8576 6734 8628 6740
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8484 6656 8536 6662
rect 8484 6598 8536 6604
rect 8496 6390 8524 6598
rect 8484 6384 8536 6390
rect 8484 6326 8536 6332
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8300 6112 8352 6118
rect 8300 6054 8352 6060
rect 8312 5710 8340 6054
rect 8404 5914 8432 6258
rect 8392 5908 8444 5914
rect 8392 5850 8444 5856
rect 8588 5710 8616 6734
rect 8850 6624 8906 6633
rect 8850 6559 8906 6568
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8576 5704 8628 5710
rect 8576 5646 8628 5652
rect 8864 5302 8892 6559
rect 8956 5642 8984 6734
rect 9586 5808 9642 5817
rect 9586 5743 9588 5752
rect 9640 5743 9642 5752
rect 9588 5714 9640 5720
rect 8944 5636 8996 5642
rect 8944 5578 8996 5584
rect 9036 5568 9088 5574
rect 9036 5510 9088 5516
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8208 4684 8260 4690
rect 8208 4626 8260 4632
rect 8944 4684 8996 4690
rect 8944 4626 8996 4632
rect 8220 4185 8248 4626
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4282 8340 4558
rect 8576 4548 8628 4554
rect 8576 4490 8628 4496
rect 8484 4480 8536 4486
rect 8484 4422 8536 4428
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8496 4214 8524 4422
rect 8484 4208 8536 4214
rect 8206 4176 8262 4185
rect 8484 4150 8536 4156
rect 8206 4111 8262 4120
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 8404 3738 8432 4082
rect 8392 3732 8444 3738
rect 8392 3674 8444 3680
rect 8588 3398 8616 4490
rect 8956 3534 8984 4626
rect 8944 3528 8996 3534
rect 8944 3470 8996 3476
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8588 3058 8616 3334
rect 8576 3052 8628 3058
rect 8576 2994 8628 3000
rect 8300 2984 8352 2990
rect 8300 2926 8352 2932
rect 8024 2848 8076 2854
rect 8024 2790 8076 2796
rect 8036 2446 8064 2790
rect 8024 2440 8076 2446
rect 8024 2382 8076 2388
rect 7668 2106 7696 2314
rect 7744 2300 7776 2356
rect 7832 2300 7856 2356
rect 7912 2300 7944 2356
rect 7744 2276 7944 2300
rect 7744 2220 7776 2276
rect 7832 2220 7856 2276
rect 7912 2220 7944 2276
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7576 1414 7696 1442
rect 7668 1358 7696 1414
rect 7656 1352 7708 1358
rect 7656 1294 7708 1300
rect 7744 1040 7944 2220
rect 8312 1834 8340 2926
rect 8588 2446 8616 2994
rect 9048 2446 9076 5510
rect 9588 5160 9640 5166
rect 9588 5102 9640 5108
rect 9600 5001 9628 5102
rect 9586 4992 9642 5001
rect 9586 4927 9642 4936
rect 9126 3360 9182 3369
rect 9126 3295 9182 3304
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 9036 2440 9088 2446
rect 9036 2382 9088 2388
rect 8588 1970 8616 2382
rect 9048 2038 9076 2382
rect 9036 2032 9088 2038
rect 9036 1974 9088 1980
rect 8576 1964 8628 1970
rect 8576 1906 8628 1912
rect 8300 1828 8352 1834
rect 8300 1770 8352 1776
rect 9140 1426 9168 3295
rect 9588 1896 9640 1902
rect 9588 1838 9640 1844
rect 9600 1737 9628 1838
rect 9586 1728 9642 1737
rect 9586 1663 9642 1672
rect 9128 1420 9180 1426
rect 9128 1362 9180 1368
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 6544 988 6744 1020
rect 9048 921 9076 1294
rect 9034 912 9090 921
rect 9034 847 9090 856
<< via2 >>
rect 478 11736 534 11792
rect 1030 10920 1086 10976
rect 478 10124 534 10160
rect 478 10104 480 10124
rect 480 10104 532 10124
rect 532 10104 534 10124
rect 386 9288 442 9344
rect 1398 12824 1454 12880
rect 1398 12552 1454 12608
rect 938 7656 994 7712
rect 478 6024 534 6080
rect 386 5208 442 5264
rect 386 4392 442 4448
rect 1214 6840 1270 6896
rect 1030 3576 1086 3632
rect 3376 13900 3432 13956
rect 3456 13900 3512 13956
rect 2976 13500 3032 13556
rect 3056 13500 3112 13556
rect 2976 13420 3032 13476
rect 3056 13420 3112 13476
rect 2576 13100 2632 13156
rect 2656 13100 2712 13156
rect 2576 13020 2632 13076
rect 2656 13020 2712 13076
rect 2134 11192 2190 11248
rect 2318 12164 2374 12200
rect 2318 12144 2320 12164
rect 2320 12144 2372 12164
rect 2372 12144 2374 12164
rect 2042 8608 2098 8664
rect 1582 3168 1638 3224
rect 938 2760 994 2816
rect 3376 13820 3432 13876
rect 3456 13820 3512 13876
rect 2410 11328 2466 11384
rect 3606 12144 3662 12200
rect 4158 11192 4214 11248
rect 3776 10300 3832 10356
rect 3856 10300 3912 10356
rect 3776 10220 3832 10276
rect 3856 10220 3912 10276
rect 3376 9900 3432 9956
rect 3456 9900 3512 9956
rect 3376 9820 3432 9876
rect 3456 9820 3512 9876
rect 2976 9500 3032 9556
rect 3056 9500 3112 9556
rect 2976 9420 3032 9476
rect 3056 9420 3112 9476
rect 2576 9100 2632 9156
rect 2656 9100 2712 9156
rect 2576 9020 2632 9076
rect 2656 9020 2712 9076
rect 3238 8744 3294 8800
rect 2576 5100 2632 5156
rect 2656 5100 2712 5156
rect 2576 5020 2632 5076
rect 2656 5020 2712 5076
rect 3238 8608 3294 8664
rect 2976 5500 3032 5556
rect 3056 5500 3112 5556
rect 2976 5466 3032 5476
rect 3056 5466 3112 5476
rect 2976 5420 3006 5466
rect 3006 5420 3018 5466
rect 3018 5420 3032 5466
rect 3056 5420 3070 5466
rect 3070 5420 3082 5466
rect 3082 5420 3112 5466
rect 3776 6300 3832 6356
rect 3856 6300 3912 6356
rect 3776 6220 3832 6276
rect 3856 6220 3912 6276
rect 3376 5900 3432 5956
rect 3456 5900 3512 5956
rect 3376 5820 3432 5876
rect 3456 5820 3512 5876
rect 386 2488 442 2544
rect 1950 2488 2006 2544
rect 932 2300 988 2356
rect 1012 2300 1068 2356
rect 932 2220 988 2276
rect 1012 2220 1068 2276
rect 386 1944 442 2000
rect 1532 1900 1588 1956
rect 1612 1900 1668 1956
rect 1532 1820 1588 1876
rect 1612 1820 1668 1876
rect 3776 2300 3832 2356
rect 3856 2300 3912 2356
rect 3776 2220 3832 2276
rect 3856 2220 3912 2276
rect 6576 13100 6632 13156
rect 6656 13100 6712 13156
rect 6576 13020 6632 13076
rect 6656 13020 6712 13076
rect 7376 13900 7432 13956
rect 7456 13900 7512 13956
rect 7376 13820 7432 13876
rect 7456 13820 7512 13876
rect 6976 13500 7032 13556
rect 7056 13500 7112 13556
rect 6976 13420 7032 13476
rect 7056 13420 7112 13476
rect 6274 11328 6330 11384
rect 6976 9500 7032 9556
rect 7056 9500 7112 9556
rect 6976 9420 7032 9476
rect 7056 9420 7112 9476
rect 6576 9100 6632 9156
rect 6656 9100 6712 9156
rect 6576 9020 6632 9076
rect 6656 9020 6712 9076
rect 7376 9900 7432 9956
rect 7456 9900 7512 9956
rect 7376 9820 7432 9876
rect 7456 9820 7512 9876
rect 7194 8236 7196 8256
rect 7196 8236 7248 8256
rect 7248 8236 7250 8256
rect 7194 8200 7250 8236
rect 6576 5100 6632 5156
rect 6656 5100 6712 5156
rect 6576 5020 6632 5076
rect 6656 5020 6712 5076
rect 5906 4120 5962 4176
rect 6274 4120 6330 4176
rect 5630 2488 5686 2544
rect 6458 3188 6514 3224
rect 6458 3168 6460 3188
rect 6460 3168 6512 3188
rect 6512 3168 6514 3188
rect 6976 5500 7032 5556
rect 7056 5500 7112 5556
rect 6976 5466 7032 5476
rect 7056 5466 7112 5476
rect 6976 5420 7006 5466
rect 7006 5420 7018 5466
rect 7018 5420 7032 5466
rect 7056 5420 7070 5466
rect 7070 5420 7082 5466
rect 7082 5420 7112 5466
rect 7776 10300 7832 10356
rect 7856 10300 7912 10356
rect 7776 10220 7832 10276
rect 7856 10220 7912 10276
rect 7376 5900 7432 5956
rect 7456 5900 7512 5956
rect 7376 5820 7432 5876
rect 7456 5820 7512 5876
rect 6576 1100 6632 1156
rect 6656 1100 6712 1156
rect 6576 1020 6632 1076
rect 6656 1020 6712 1076
rect 6976 1500 7032 1556
rect 7056 1500 7112 1556
rect 6976 1420 7032 1476
rect 7056 1420 7112 1476
rect 7376 1900 7432 1956
rect 7456 1900 7512 1956
rect 7376 1820 7432 1876
rect 7456 1820 7512 1876
rect 8482 12416 8538 12472
rect 8390 12280 8446 12336
rect 8666 12588 8668 12608
rect 8668 12588 8720 12608
rect 8720 12588 8722 12608
rect 8666 12552 8722 12588
rect 8850 12824 8906 12880
rect 8574 11464 8630 11520
rect 8114 10648 8170 10704
rect 7776 6300 7832 6356
rect 7856 6300 7912 6356
rect 7776 6220 7832 6276
rect 7856 6220 7912 6276
rect 8390 7384 8446 7440
rect 9586 13948 9588 13968
rect 9588 13948 9640 13968
rect 9640 13948 9642 13968
rect 9586 13912 9642 13948
rect 9586 13096 9642 13152
rect 9586 9832 9642 9888
rect 9586 9016 9642 9072
rect 8850 6568 8906 6624
rect 9586 5772 9642 5808
rect 9586 5752 9588 5772
rect 9588 5752 9640 5772
rect 9640 5752 9642 5772
rect 8206 4120 8262 4176
rect 7776 2300 7832 2356
rect 7856 2300 7912 2356
rect 7776 2220 7832 2276
rect 7856 2220 7912 2276
rect 9586 4936 9642 4992
rect 9126 3304 9182 3360
rect 9586 1672 9642 1728
rect 9034 856 9090 912
<< metal3 >>
rect 596 13956 9432 13988
rect 9600 13973 10200 14000
rect 596 13900 3376 13956
rect 3432 13900 3456 13956
rect 3512 13900 7376 13956
rect 7432 13900 7456 13956
rect 7512 13900 9432 13956
rect 9581 13968 10200 13973
rect 9581 13912 9586 13968
rect 9642 13912 10200 13968
rect 9581 13907 10200 13912
rect 596 13876 9432 13900
rect 9600 13880 10200 13907
rect 596 13820 3376 13876
rect 3432 13820 3456 13876
rect 3512 13820 7376 13876
rect 7432 13820 7456 13876
rect 7512 13820 9432 13876
rect 596 13788 9432 13820
rect 596 13556 9432 13588
rect 596 13500 2976 13556
rect 3032 13500 3056 13556
rect 3112 13500 6976 13556
rect 7032 13500 7056 13556
rect 7112 13500 9432 13556
rect 596 13476 9432 13500
rect 596 13420 2976 13476
rect 3032 13420 3056 13476
rect 3112 13420 6976 13476
rect 7032 13420 7056 13476
rect 7112 13420 9432 13476
rect 596 13388 9432 13420
rect 596 13156 9432 13188
rect 9600 13157 10200 13184
rect 596 13100 2576 13156
rect 2632 13100 2656 13156
rect 2712 13100 6576 13156
rect 6632 13100 6656 13156
rect 6712 13100 9432 13156
rect 596 13076 9432 13100
rect 9581 13152 10200 13157
rect 9581 13096 9586 13152
rect 9642 13096 10200 13152
rect 9581 13091 10200 13096
rect 596 13020 2576 13076
rect 2632 13020 2656 13076
rect 2712 13020 6576 13076
rect 6632 13020 6656 13076
rect 6712 13020 9432 13076
rect 9600 13064 10200 13091
rect 596 12988 9432 13020
rect 1393 12882 1459 12885
rect 8845 12882 8911 12885
rect 1393 12880 8911 12882
rect 1393 12824 1398 12880
rect 1454 12824 8850 12880
rect 8906 12824 8911 12880
rect 1393 12822 8911 12824
rect 1393 12819 1459 12822
rect 8845 12819 8911 12822
rect -200 12610 400 12640
rect 1393 12610 1459 12613
rect 8661 12610 8727 12613
rect -200 12608 1459 12610
rect -200 12552 1398 12608
rect 1454 12552 1459 12608
rect -200 12550 1459 12552
rect -200 12520 400 12550
rect 1393 12547 1459 12550
rect 8526 12608 8727 12610
rect 8526 12552 8666 12608
rect 8722 12552 8727 12608
rect 8526 12550 8727 12552
rect 8526 12477 8586 12550
rect 8661 12547 8727 12550
rect 8477 12472 8586 12477
rect 8477 12416 8482 12472
rect 8538 12416 8586 12472
rect 8477 12414 8586 12416
rect 8477 12411 8543 12414
rect 8385 12338 8451 12341
rect 9600 12338 10200 12368
rect 8385 12336 10200 12338
rect 8385 12280 8390 12336
rect 8446 12280 10200 12336
rect 8385 12278 10200 12280
rect 8385 12275 8451 12278
rect 9600 12248 10200 12278
rect 2313 12202 2379 12205
rect 3601 12202 3667 12205
rect 2313 12200 3667 12202
rect 2313 12144 2318 12200
rect 2374 12144 3606 12200
rect 3662 12144 3667 12200
rect 2313 12142 3667 12144
rect 2313 12139 2379 12142
rect 3601 12139 3667 12142
rect -200 11794 400 11824
rect 473 11794 539 11797
rect -200 11792 539 11794
rect -200 11736 478 11792
rect 534 11736 539 11792
rect -200 11734 539 11736
rect -200 11704 400 11734
rect 473 11731 539 11734
rect 8569 11522 8635 11525
rect 9600 11522 10200 11552
rect 8569 11520 10200 11522
rect 8569 11464 8574 11520
rect 8630 11464 10200 11520
rect 8569 11462 10200 11464
rect 8569 11459 8635 11462
rect 9600 11432 10200 11462
rect 2405 11386 2471 11389
rect 6269 11386 6335 11389
rect 2405 11384 6335 11386
rect 2405 11328 2410 11384
rect 2466 11328 6274 11384
rect 6330 11328 6335 11384
rect 2405 11326 6335 11328
rect 2405 11323 2471 11326
rect 6269 11323 6335 11326
rect 2129 11250 2195 11253
rect 4153 11250 4219 11253
rect 2129 11248 4219 11250
rect 2129 11192 2134 11248
rect 2190 11192 4158 11248
rect 4214 11192 4219 11248
rect 2129 11190 4219 11192
rect 2129 11187 2195 11190
rect 4153 11187 4219 11190
rect -200 10978 400 11008
rect 1025 10978 1091 10981
rect -200 10976 1091 10978
rect -200 10920 1030 10976
rect 1086 10920 1091 10976
rect -200 10918 1091 10920
rect -200 10888 400 10918
rect 1025 10915 1091 10918
rect 8109 10706 8175 10709
rect 9600 10706 10200 10736
rect 8109 10704 10200 10706
rect 8109 10648 8114 10704
rect 8170 10648 10200 10704
rect 8109 10646 10200 10648
rect 8109 10643 8175 10646
rect 9600 10616 10200 10646
rect 596 10356 9432 10388
rect 596 10300 3776 10356
rect 3832 10300 3856 10356
rect 3912 10300 7776 10356
rect 7832 10300 7856 10356
rect 7912 10300 9432 10356
rect 596 10276 9432 10300
rect 596 10220 3776 10276
rect 3832 10220 3856 10276
rect 3912 10220 7776 10276
rect 7832 10220 7856 10276
rect 7912 10220 9432 10276
rect -200 10162 400 10192
rect 596 10188 9432 10220
rect 473 10162 539 10165
rect -200 10160 539 10162
rect -200 10104 478 10160
rect 534 10104 539 10160
rect -200 10102 539 10104
rect -200 10072 400 10102
rect 473 10099 539 10102
rect 596 9956 9432 9988
rect 596 9900 3376 9956
rect 3432 9900 3456 9956
rect 3512 9900 7376 9956
rect 7432 9900 7456 9956
rect 7512 9900 9432 9956
rect 596 9876 9432 9900
rect 9600 9893 10200 9920
rect 596 9820 3376 9876
rect 3432 9820 3456 9876
rect 3512 9820 7376 9876
rect 7432 9820 7456 9876
rect 7512 9820 9432 9876
rect 9581 9888 10200 9893
rect 9581 9832 9586 9888
rect 9642 9832 10200 9888
rect 9581 9827 10200 9832
rect 596 9788 9432 9820
rect 9600 9800 10200 9827
rect 596 9556 9432 9588
rect 596 9500 2976 9556
rect 3032 9500 3056 9556
rect 3112 9500 6976 9556
rect 7032 9500 7056 9556
rect 7112 9500 9432 9556
rect 596 9476 9432 9500
rect 596 9420 2976 9476
rect 3032 9420 3056 9476
rect 3112 9420 6976 9476
rect 7032 9420 7056 9476
rect 7112 9420 9432 9476
rect 596 9388 9432 9420
rect -200 9349 400 9376
rect -200 9344 447 9349
rect -200 9288 386 9344
rect 442 9288 447 9344
rect -200 9283 447 9288
rect -200 9256 400 9283
rect 596 9156 9432 9188
rect 596 9100 2576 9156
rect 2632 9100 2656 9156
rect 2712 9100 6576 9156
rect 6632 9100 6656 9156
rect 6712 9100 9432 9156
rect 596 9076 9432 9100
rect 9600 9077 10200 9104
rect 596 9020 2576 9076
rect 2632 9020 2656 9076
rect 2712 9020 6576 9076
rect 6632 9020 6656 9076
rect 6712 9020 9432 9076
rect 596 8988 9432 9020
rect 9581 9072 10200 9077
rect 9581 9016 9586 9072
rect 9642 9016 10200 9072
rect 9581 9011 10200 9016
rect 9600 8984 10200 9011
rect 3233 8802 3299 8805
rect 1580 8800 3299 8802
rect 1580 8744 3238 8800
rect 3294 8744 3299 8800
rect 1580 8742 3299 8744
rect -200 8530 400 8560
rect 1580 8530 1640 8742
rect 3233 8739 3299 8742
rect 2037 8666 2103 8669
rect 3233 8666 3299 8669
rect 2037 8664 3299 8666
rect 2037 8608 2042 8664
rect 2098 8608 3238 8664
rect 3294 8608 3299 8664
rect 2037 8606 3299 8608
rect 2037 8603 2103 8606
rect 3233 8603 3299 8606
rect -200 8470 1640 8530
rect -200 8440 400 8470
rect 7189 8258 7255 8261
rect 9600 8258 10200 8288
rect 7189 8256 10200 8258
rect 7189 8200 7194 8256
rect 7250 8200 10200 8256
rect 7189 8198 10200 8200
rect 7189 8195 7255 8198
rect 9600 8168 10200 8198
rect -200 7714 400 7744
rect 933 7714 999 7717
rect -200 7712 999 7714
rect -200 7656 938 7712
rect 994 7656 999 7712
rect -200 7654 999 7656
rect -200 7624 400 7654
rect 933 7651 999 7654
rect 8385 7442 8451 7445
rect 9600 7442 10200 7472
rect 8385 7440 10200 7442
rect 8385 7384 8390 7440
rect 8446 7384 10200 7440
rect 8385 7382 10200 7384
rect 8385 7379 8451 7382
rect 9600 7352 10200 7382
rect -200 6898 400 6928
rect 1209 6898 1275 6901
rect -200 6896 1275 6898
rect -200 6840 1214 6896
rect 1270 6840 1275 6896
rect -200 6838 1275 6840
rect -200 6808 400 6838
rect 1209 6835 1275 6838
rect 8845 6626 8911 6629
rect 9600 6626 10200 6656
rect 8845 6624 10200 6626
rect 8845 6568 8850 6624
rect 8906 6568 10200 6624
rect 8845 6566 10200 6568
rect 8845 6563 8911 6566
rect 9600 6536 10200 6566
rect 596 6356 9432 6388
rect 596 6300 3776 6356
rect 3832 6300 3856 6356
rect 3912 6300 7776 6356
rect 7832 6300 7856 6356
rect 7912 6300 9432 6356
rect 596 6276 9432 6300
rect 596 6220 3776 6276
rect 3832 6220 3856 6276
rect 3912 6220 7776 6276
rect 7832 6220 7856 6276
rect 7912 6220 9432 6276
rect 596 6188 9432 6220
rect -200 6082 400 6112
rect 473 6082 539 6085
rect -200 6080 539 6082
rect -200 6024 478 6080
rect 534 6024 539 6080
rect -200 6022 539 6024
rect -200 5992 400 6022
rect 473 6019 539 6022
rect 596 5956 9432 5988
rect 596 5900 3376 5956
rect 3432 5900 3456 5956
rect 3512 5900 7376 5956
rect 7432 5900 7456 5956
rect 7512 5900 9432 5956
rect 596 5876 9432 5900
rect 596 5820 3376 5876
rect 3432 5820 3456 5876
rect 3512 5820 7376 5876
rect 7432 5820 7456 5876
rect 7512 5820 9432 5876
rect 596 5788 9432 5820
rect 9600 5813 10200 5840
rect 9581 5808 10200 5813
rect 9581 5752 9586 5808
rect 9642 5752 10200 5808
rect 9581 5747 10200 5752
rect 9600 5720 10200 5747
rect 596 5556 9432 5588
rect 596 5500 2976 5556
rect 3032 5500 3056 5556
rect 3112 5500 6976 5556
rect 7032 5500 7056 5556
rect 7112 5500 9432 5556
rect 596 5476 9432 5500
rect 596 5420 2976 5476
rect 3032 5420 3056 5476
rect 3112 5420 6976 5476
rect 7032 5420 7056 5476
rect 7112 5420 9432 5476
rect 596 5388 9432 5420
rect -200 5269 400 5296
rect -200 5264 447 5269
rect -200 5208 386 5264
rect 442 5208 447 5264
rect -200 5203 447 5208
rect -200 5176 400 5203
rect 596 5156 9432 5188
rect 596 5100 2576 5156
rect 2632 5100 2656 5156
rect 2712 5100 6576 5156
rect 6632 5100 6656 5156
rect 6712 5100 9432 5156
rect 596 5076 9432 5100
rect 596 5020 2576 5076
rect 2632 5020 2656 5076
rect 2712 5020 6576 5076
rect 6632 5020 6656 5076
rect 6712 5020 9432 5076
rect 596 4988 9432 5020
rect 9600 4997 10200 5024
rect 9581 4992 10200 4997
rect 9581 4936 9586 4992
rect 9642 4936 10200 4992
rect 9581 4931 10200 4936
rect 9600 4904 10200 4931
rect -200 4453 400 4480
rect -200 4448 447 4453
rect -200 4392 386 4448
rect 442 4392 447 4448
rect -200 4387 447 4392
rect -200 4360 400 4387
rect 5901 4178 5967 4181
rect 6269 4178 6335 4181
rect 5901 4176 6335 4178
rect 5901 4120 5906 4176
rect 5962 4120 6274 4176
rect 6330 4120 6335 4176
rect 5901 4118 6335 4120
rect 5901 4115 5967 4118
rect 6269 4115 6335 4118
rect 8201 4178 8267 4181
rect 9600 4178 10200 4208
rect 8201 4176 10200 4178
rect 8201 4120 8206 4176
rect 8262 4120 10200 4176
rect 8201 4118 10200 4120
rect 8201 4115 8267 4118
rect 9600 4088 10200 4118
rect -200 3634 400 3664
rect 1025 3634 1091 3637
rect -200 3632 1091 3634
rect -200 3576 1030 3632
rect 1086 3576 1091 3632
rect -200 3574 1091 3576
rect -200 3544 400 3574
rect 1025 3571 1091 3574
rect 9121 3362 9187 3365
rect 9600 3362 10200 3392
rect 9121 3360 10200 3362
rect 9121 3304 9126 3360
rect 9182 3304 10200 3360
rect 9121 3302 10200 3304
rect 9121 3299 9187 3302
rect 9600 3272 10200 3302
rect 1577 3226 1643 3229
rect 6453 3226 6519 3229
rect 1577 3224 6519 3226
rect 1577 3168 1582 3224
rect 1638 3168 6458 3224
rect 6514 3168 6519 3224
rect 1577 3166 6519 3168
rect 1577 3163 1643 3166
rect 6453 3163 6519 3166
rect -200 2818 400 2848
rect 933 2818 999 2821
rect -200 2816 999 2818
rect -200 2760 938 2816
rect 994 2760 999 2816
rect -200 2758 999 2760
rect -200 2728 400 2758
rect 933 2755 999 2758
rect 381 2546 447 2549
rect 1945 2546 2011 2549
rect 381 2544 2011 2546
rect 381 2488 386 2544
rect 442 2488 1950 2544
rect 2006 2488 2011 2544
rect 381 2486 2011 2488
rect 381 2483 447 2486
rect 1945 2483 2011 2486
rect 5625 2546 5691 2549
rect 9600 2546 10200 2576
rect 5625 2544 10200 2546
rect 5625 2488 5630 2544
rect 5686 2488 10200 2544
rect 5625 2486 10200 2488
rect 5625 2483 5691 2486
rect 9600 2456 10200 2486
rect 596 2356 9432 2388
rect 596 2300 932 2356
rect 988 2300 1012 2356
rect 1068 2300 3776 2356
rect 3832 2300 3856 2356
rect 3912 2300 7776 2356
rect 7832 2300 7856 2356
rect 7912 2300 9432 2356
rect 596 2276 9432 2300
rect 596 2220 932 2276
rect 988 2220 1012 2276
rect 1068 2220 3776 2276
rect 3832 2220 3856 2276
rect 3912 2220 7776 2276
rect 7832 2220 7856 2276
rect 7912 2220 9432 2276
rect 596 2188 9432 2220
rect -200 2005 400 2032
rect -200 2000 447 2005
rect -200 1944 386 2000
rect 442 1944 447 2000
rect -200 1939 447 1944
rect 596 1956 9432 1988
rect -200 1912 400 1939
rect 596 1900 1532 1956
rect 1588 1900 1612 1956
rect 1668 1900 7376 1956
rect 7432 1900 7456 1956
rect 7512 1900 9432 1956
rect 596 1876 9432 1900
rect 596 1820 1532 1876
rect 1588 1820 1612 1876
rect 1668 1820 7376 1876
rect 7432 1820 7456 1876
rect 7512 1820 9432 1876
rect 596 1788 9432 1820
rect 9600 1733 10200 1760
rect 9581 1728 10200 1733
rect 9581 1672 9586 1728
rect 9642 1672 10200 1728
rect 9581 1667 10200 1672
rect 9600 1640 10200 1667
rect 596 1556 9432 1588
rect 596 1500 6976 1556
rect 7032 1500 7056 1556
rect 7112 1500 9432 1556
rect 596 1476 9432 1500
rect 596 1420 6976 1476
rect 7032 1420 7056 1476
rect 7112 1420 9432 1476
rect 596 1388 9432 1420
rect 596 1156 9432 1188
rect 596 1100 6576 1156
rect 6632 1100 6656 1156
rect 6712 1100 9432 1156
rect 596 1076 9432 1100
rect 596 1020 6576 1076
rect 6632 1020 6656 1076
rect 6712 1020 9432 1076
rect 596 988 9432 1020
rect 9029 914 9095 917
rect 9600 914 10200 944
rect 9029 912 10200 914
rect 9029 856 9034 912
rect 9090 856 10200 912
rect 9029 854 10200 856
rect 9029 851 9095 854
rect 9600 824 10200 854
use sky130_fd_sc_hd__inv_2  _057_
timestamp 1562557784
transform 1 0 5612 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _058_
timestamp 1562557784
transform -1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2b_1  _059_
timestamp 21601
transform -1 0 8924 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _060_
timestamp 21601
transform 1 0 8556 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _061_
timestamp 21601
transform -1 0 8924 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _062_
timestamp 21601
transform 1 0 5888 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _063_
timestamp 21601
transform -1 0 8924 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _064_
timestamp 21601
transform 1 0 6808 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _065_
timestamp 21601
transform -1 0 5796 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _066_
timestamp 21601
transform -1 0 8924 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _067_
timestamp 21601
transform -1 0 6348 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _068_
timestamp 21601
transform 1 0 3496 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _069_
timestamp 21601
transform -1 0 8924 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _070_
timestamp 21601
transform 1 0 6808 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _071_
timestamp 21601
transform -1 0 5612 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nand2b_1  _072_
timestamp 21601
transform -1 0 2944 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _073_
timestamp 21601
transform -1 0 1840 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 21601
transform -1 0 2668 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _075_
timestamp 21601
transform -1 0 3220 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _076_
timestamp 21601
transform 1 0 3864 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _077_
timestamp 21601
transform -1 0 5704 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _078_
timestamp 21601
transform 1 0 8464 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _079_
timestamp 21601
transform -1 0 8924 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _080_
timestamp 21601
transform 1 0 3496 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _081_
timestamp 21601
transform 1 0 8464 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _082_
timestamp 21601
transform -1 0 8924 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _083_
timestamp 21601
transform 1 0 8648 0 -1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _084_
timestamp 21601
transform -1 0 8924 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _085_
timestamp 21601
transform 1 0 5612 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _086_
timestamp 21601
transform 1 0 8648 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _087_
timestamp 21601
transform -1 0 8924 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _088_
timestamp 21601
transform 1 0 6072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _089_
timestamp 21601
transform -1 0 8924 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _090_
timestamp 1562557784
transform -1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _091_
timestamp 1562557784
transform -1 0 6900 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _092_
timestamp 1562557784
transform -1 0 7544 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _093_
timestamp 1562557784
transform 1 0 6256 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _094_
timestamp 1562557784
transform 1 0 5060 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _095_
timestamp 1562557784
transform 1 0 4232 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _096_
timestamp 1562557784
transform 1 0 5520 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _097_
timestamp 1562557784
transform 1 0 2944 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _098_
timestamp 1562557784
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _099_
timestamp 1562557784
transform 1 0 8004 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _100_
timestamp 1562557784
transform 1 0 4784 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _101_
timestamp 1562557784
transform 1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1562557784
transform 1 0 1012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _103_
timestamp 21601
transform 1 0 1288 0 -1 8704
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _104_
timestamp 21601
transform 1 0 3496 0 1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _105_
timestamp 21601
transform 1 0 5980 0 1 2176
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _106_
timestamp 21601
transform 1 0 6348 0 -1 11968
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _107_
timestamp 21601
transform 1 0 3220 0 -1 13056
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _108_
timestamp 21601
transform 1 0 4692 0 1 11968
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _109_
timestamp 21601
transform 1 0 6532 0 -1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _110_
timestamp 21601
transform -1 0 7636 0 -1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _111_
timestamp 21601
transform 1 0 6532 0 -1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _112_
timestamp 21601
transform 1 0 4508 0 1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _113_
timestamp 21601
transform 1 0 6072 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _114_
timestamp 21601
transform 1 0 6532 0 -1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _115_
timestamp 21601
transform 1 0 6532 0 -1 13056
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_1  _116_
timestamp 21601
transform 1 0 920 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _117_
timestamp 21601
transform 1 0 1012 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _118_
timestamp 21601
transform 1 0 1932 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _119_
timestamp 21601
transform -1 0 3220 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _120_
timestamp 21601
transform 1 0 2760 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _121_
timestamp 21601
transform -1 0 4968 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _122_
timestamp 21601
transform 1 0 3864 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _123_
timestamp 21601
transform 1 0 4784 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _124_
timestamp 21601
transform 1 0 3680 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _125_
timestamp 21601
transform -1 0 5796 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _126_
timestamp 21601
transform -1 0 6716 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _127_
timestamp 21601
transform 1 0 4876 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _128_
timestamp 21601
transform 1 0 5888 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _129_
timestamp 21601
transform -1 0 6808 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _130_
timestamp 21601
transform -1 0 5152 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _131_
timestamp 21601
transform 1 0 3956 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfbbn_2  _132_
timestamp 21601
transform 1 0 6348 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_1  _133_
timestamp 21601
transform -1 0 2760 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 21601
transform -1 0 1472 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _136_
timestamp 21601
transform -1 0 6900 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[0\]
timestamp 21601
transform -1 0 1932 0 -1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[1\]
timestamp 21601
transform -1 0 1932 0 1 9792
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  BUF\[2\]
timestamp 21601
transform -1 0 1932 0 1 10880
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_2  fanout39
timestamp 21601
transform 1 0 6072 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  fanout40
timestamp 21601
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  fanout41
timestamp 21601
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  fanout42
timestamp 21601
transform -1 0 2300 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  fanout43
timestamp 21601
transform 1 0 1840 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23
timestamp 21601
transform 1 0 2760 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26
timestamp 21601
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29
timestamp 21601
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32
timestamp 21601
transform 1 0 3588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35
timestamp 21601
transform 1 0 3864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38
timestamp 21601
transform 1 0 4140 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41
timestamp 21601
transform 1 0 4416 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44
timestamp 21601
transform 1 0 4692 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 21601
transform 1 0 4968 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49
timestamp 21601
transform 1 0 5152 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52
timestamp 21601
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55
timestamp 21601
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58
timestamp 21601
transform 1 0 5980 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77
timestamp 21601
transform 1 0 7728 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_80
timestamp 21601
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_83
timestamp 21601
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_86
timestamp 21601
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_23
timestamp 21601
transform 1 0 2760 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_26
timestamp 21601
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_29
timestamp 21601
transform 1 0 3312 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 21601
transform 1 0 6716 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_72
timestamp 21601
transform 1 0 7268 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_75
timestamp 21601
transform 1 0 7544 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_77
timestamp 21601
transform 1 0 7728 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_80
timestamp 21601
transform 1 0 8004 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_1_83
timestamp 21601
transform 1 0 8280 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_86
timestamp 21601
transform 1 0 8556 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_2_28
timestamp 21601
transform 1 0 3220 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_31
timestamp 21601
transform 1 0 3496 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_34
timestamp 21601
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_37
timestamp 21601
transform 1 0 4048 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_2_40
timestamp 21601
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_2_43
timestamp 21601
transform 1 0 4600 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_57
timestamp 21601
transform 1 0 5888 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_91
timestamp 21601
transform 1 0 9016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_23
timestamp 21601
transform 1 0 2760 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_26
timestamp 21601
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_3_29
timestamp 21601
transform 1 0 3312 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_3_90
timestamp 21601
transform 1 0 8924 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_4_3
timestamp 21601
transform 1 0 920 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_6
timestamp 21601
transform 1 0 1196 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_9
timestamp 21601
transform 1 0 1472 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_12
timestamp 21601
transform 1 0 1748 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_15
timestamp 21601
transform 1 0 2024 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_18
timestamp 21601
transform 1 0 2300 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_21
timestamp 21601
transform 1 0 2576 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_24
timestamp 21601
transform 1 0 2852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 21601
transform 1 0 3128 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_29
timestamp 21601
transform 1 0 3312 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_4_32
timestamp 21601
transform 1 0 3588 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_35
timestamp 21601
transform 1 0 3864 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_4_80
timestamp 21601
transform 1 0 8004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 21601
transform 1 0 8280 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_90
timestamp 21601
transform 1 0 8924 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_5_3
timestamp 21601
transform 1 0 920 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_6
timestamp 21601
transform 1 0 1196 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_9
timestamp 21601
transform 1 0 1472 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_12
timestamp 21601
transform 1 0 1748 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_15
timestamp 21601
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_18
timestamp 21601
transform 1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_21
timestamp 21601
transform 1 0 2576 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_24
timestamp 21601
transform 1 0 2852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_27
timestamp 21601
transform 1 0 3128 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_5_30
timestamp 21601
transform 1 0 3404 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_5_57
timestamp 21601
transform 1 0 5888 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 21601
transform 1 0 6440 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_9
timestamp 21601
transform 1 0 1472 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_6_12
timestamp 21601
transform 1 0 1748 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_17
timestamp 21601
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_20
timestamp 21601
transform 1 0 2484 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_23
timestamp 21601
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_26
timestamp 21601
transform 1 0 3036 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_6_29
timestamp 21601
transform 1 0 3312 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_32
timestamp 21601
transform 1 0 3588 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_6_35
timestamp 21601
transform 1 0 3864 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_66
timestamp 21601
transform 1 0 6716 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_90
timestamp 21601
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_7_23
timestamp 21601
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_26
timestamp 21601
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_29
timestamp 21601
transform 1 0 3312 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_32
timestamp 21601
transform 1 0 3588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_35
timestamp 21601
transform 1 0 3864 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_38
timestamp 21601
transform 1 0 4140 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_41
timestamp 21601
transform 1 0 4416 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_7_44
timestamp 21601
transform 1 0 4692 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_7_47
timestamp 21601
transform 1 0 4968 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_57
timestamp 21601
transform 1 0 5888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_19
timestamp 21601
transform 1 0 2392 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_22
timestamp 21601
transform 1 0 2668 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 21601
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_29
timestamp 21601
transform 1 0 3312 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_32
timestamp 21601
transform 1 0 3588 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_35
timestamp 21601
transform 1 0 3864 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_38
timestamp 21601
transform 1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_41
timestamp 21601
transform 1 0 4416 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_8_44
timestamp 21601
transform 1 0 4692 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_8_90
timestamp 21601
transform 1 0 8924 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_9_6
timestamp 21601
transform 1 0 1196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_9
timestamp 21601
transform 1 0 1472 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_12
timestamp 21601
transform 1 0 1748 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_15
timestamp 21601
transform 1 0 2024 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_18
timestamp 21601
transform 1 0 2300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_21
timestamp 21601
transform 1 0 2576 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_24
timestamp 21601
transform 1 0 2852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_27
timestamp 21601
transform 1 0 3128 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_9_30
timestamp 21601
transform 1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_9_33
timestamp 21601
transform 1 0 3680 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 21601
transform 1 0 5704 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_57
timestamp 21601
transform 1 0 5888 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_3
timestamp 21601
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_6
timestamp 21601
transform 1 0 1196 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_9
timestamp 21601
transform 1 0 1472 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_12
timestamp 21601
transform 1 0 1748 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_15
timestamp 21601
transform 1 0 2024 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_18
timestamp 21601
transform 1 0 2300 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_21
timestamp 21601
transform 1 0 2576 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_24
timestamp 21601
transform 1 0 2852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 21601
transform 1 0 3128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_10_29
timestamp 21601
transform 1 0 3312 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_32
timestamp 21601
transform 1 0 3588 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_10_35
timestamp 21601
transform 1 0 3864 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_10_38
timestamp 21601
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_70
timestamp 21601
transform 1 0 7084 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_80
timestamp 21601
transform 1 0 8004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_90
timestamp 21601
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_11_9
timestamp 21601
transform 1 0 1472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_12
timestamp 21601
transform 1 0 1748 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_11_15
timestamp 21601
transform 1 0 2024 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_11_25
timestamp 21601
transform 1 0 2944 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_11_47
timestamp 21601
transform 1 0 4968 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_57
timestamp 21601
transform 1 0 5888 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 21601
transform 1 0 920 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_12_22
timestamp 21601
transform 1 0 2668 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 21601
transform 1 0 2944 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_29
timestamp 21601
transform 1 0 3312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_32
timestamp 21601
transform 1 0 3588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_12_35
timestamp 21601
transform 1 0 3864 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_12_45
timestamp 21601
transform 1 0 4784 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_48
timestamp 21601
transform 1 0 5060 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_12_51
timestamp 21601
transform 1 0 5336 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_12_67
timestamp 21601
transform 1 0 6808 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_90
timestamp 21601
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 21601
transform 1 0 920 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_40
timestamp 21601
transform 1 0 4324 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_43
timestamp 21601
transform 1 0 4600 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_46
timestamp 21601
transform 1 0 4876 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_49
timestamp 21601
transform 1 0 5152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_13_52
timestamp 21601
transform 1 0 5428 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 21601
transform 1 0 5704 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_57
timestamp 21601
transform 1 0 5888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 21601
transform 1 0 7452 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_19
timestamp 21601
transform 1 0 2392 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_35
timestamp 21601
transform 1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_38
timestamp 21601
transform 1 0 4140 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_41
timestamp 21601
transform 1 0 4416 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_44
timestamp 21601
transform 1 0 4692 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 21601
transform 1 0 8280 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_14_90
timestamp 21601
transform 1 0 8924 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_3
timestamp 21601
transform 1 0 920 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_24
timestamp 21601
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_34
timestamp 21601
transform 1 0 3772 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_15_61
timestamp 21601
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_90
timestamp 21601
transform 1 0 8924 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_18
timestamp 21601
transform 1 0 2300 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_90
timestamp 21601
transform 1 0 8924 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 21601
transform 1 0 5704 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_57
timestamp 21601
transform 1 0 5888 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_14
timestamp 21601
transform 1 0 1932 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_18_29
timestamp 21601
transform 1 0 3312 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_18_59
timestamp 21601
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_90
timestamp 21601
transform 1 0 8924 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_43
timestamp 21601
transform 1 0 4600 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_90
timestamp 21601
transform 1 0 8924 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_3
timestamp 21601
transform 1 0 920 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_20_29
timestamp 21601
transform 1 0 3312 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 21601
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_90
timestamp 21601
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_21_19
timestamp 21601
transform 1 0 2392 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_62
timestamp 21601
transform 1 0 6348 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_29
timestamp 21601
transform 1 0 3312 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_22_90
timestamp 21601
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_23_3
timestamp 21601
transform 1 0 920 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_90
timestamp 21601
transform 1 0 8924 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  gpio_control_block_mgmt_monitor_44
timestamp 1562557784
transform 1 0 6440 0 -1 8704
box -38 -48 314 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 600 0 1 1252
box 0 0 1 1
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 21601
transform 1 0 1748 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 21601
transform -1 0 8004 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 21601
transform 1 0 7544 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 21601
transform -1 0 6624 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 21601
transform -1 0 1748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 21601
transform -1 0 3220 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 21601
transform -1 0 4692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 21601
transform -1 0 4324 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 21601
transform 1 0 1748 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 21601
transform -1 0 4692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 21601
transform -1 0 5428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 21601
transform 1 0 2484 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 21601
transform 1 0 2484 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 21601
transform 1 0 3772 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 21601
transform -1 0 3220 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 21601
transform 1 0 6072 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 21601
transform 1 0 4140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 21601
transform -1 0 8464 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 21601
transform 1 0 4048 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 21601
transform 1 0 5888 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 21601
transform -1 0 5244 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 21601
transform 1 0 6716 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 21601
transform 1 0 6164 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 21601
transform 1 0 5152 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 21601
transform 1 0 4784 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 21601
transform -1 0 2944 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 21601
transform -1 0 8004 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 21601
transform 1 0 5060 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 21601
transform 1 0 920 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 21601
transform 1 0 2944 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 21601
transform 1 0 3312 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 21601
transform -1 0 2668 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 21601
transform -1 0 3864 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 21601
transform -1 0 5796 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 21601
transform 1 0 6624 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 21601
transform 1 0 6164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 21601
transform -1 0 8372 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 21601
transform 1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 21601
transform -1 0 3588 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 21601
transform 1 0 3496 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 21601
transform 1 0 1472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 21601
transform -1 0 1472 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 21601
transform -1 0 1472 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 21601
transform -1 0 1196 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input17
timestamp 21601
transform -1 0 9108 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 21601
transform -1 0 1196 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 21601
transform 1 0 2944 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 21601
transform -1 0 1196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  output21
timestamp 21601
transform 1 0 920 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output22
timestamp 21601
transform 1 0 6164 0 1 1088
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output23
timestamp 21601
transform -1 0 8372 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output24
timestamp 21601
transform -1 0 8372 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output25
timestamp 21601
transform -1 0 8372 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output26
timestamp 21601
transform -1 0 5060 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output27
timestamp 21601
transform -1 0 8372 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output28
timestamp 21601
transform 1 0 6900 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output29
timestamp 21601
transform -1 0 9108 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output30
timestamp 21601
transform -1 0 6900 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output31
timestamp 21601
transform 1 0 7636 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output32
timestamp 21601
transform 1 0 6900 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output33
timestamp 21601
transform 1 0 4324 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output34
timestamp 21601
transform 1 0 6164 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output35
timestamp 21601
transform -1 0 4876 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output36
timestamp 21601
transform -1 0 8372 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output37
timestamp 21601
transform 1 0 920 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_12  output38
timestamp 21601
transform -1 0 2392 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Left_3
timestamp 21601
transform 1 0 2484 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_2_Right_27
timestamp 21601
transform -1 0 9384 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Left_0
timestamp 21601
transform 1 0 2484 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_2_Right_4
timestamp 21601
transform -1 0 9384 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Left_1
timestamp 21601
transform 1 0 2484 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_2_Right_5
timestamp 21601
transform -1 0 9384 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Left_2
timestamp 21601
transform 1 0 2484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_2_Right_6
timestamp 21601
transform -1 0 9384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_28
timestamp 21601
transform 1 0 644 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_7
timestamp 21601
transform -1 0 9384 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_29
timestamp 21601
transform 1 0 644 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_8
timestamp 21601
transform -1 0 9384 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_30
timestamp 21601
transform 1 0 644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_9
timestamp 21601
transform -1 0 9384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_31
timestamp 21601
transform 1 0 644 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_10
timestamp 21601
transform -1 0 9384 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_32
timestamp 21601
transform 1 0 644 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_11
timestamp 21601
transform -1 0 9384 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_33
timestamp 21601
transform 1 0 644 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_12
timestamp 21601
transform -1 0 9384 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_34
timestamp 21601
transform 1 0 644 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_13
timestamp 21601
transform -1 0 9384 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_35
timestamp 21601
transform 1 0 644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_14
timestamp 21601
transform -1 0 9384 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_36
timestamp 21601
transform 1 0 644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_15
timestamp 21601
transform -1 0 9384 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_37
timestamp 21601
transform 1 0 644 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_16
timestamp 21601
transform -1 0 9384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_38
timestamp 21601
transform 1 0 644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_17
timestamp 21601
transform -1 0 9384 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_39
timestamp 21601
transform 1 0 644 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_18
timestamp 21601
transform -1 0 9384 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_40
timestamp 21601
transform 1 0 644 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_19
timestamp 21601
transform -1 0 9384 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_41
timestamp 21601
transform 1 0 644 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_20
timestamp 21601
transform -1 0 9384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_42
timestamp 21601
transform 1 0 644 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_21
timestamp 21601
transform -1 0 9384 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_43
timestamp 21601
transform 1 0 644 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_22
timestamp 21601
transform -1 0 9384 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_44
timestamp 21601
transform 1 0 644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_23
timestamp 21601
transform -1 0 9384 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_45
timestamp 21601
transform 1 0 644 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_24
timestamp 21601
transform -1 0 9384 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_46
timestamp 21601
transform 1 0 644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_25
timestamp 21601
transform -1 0 9384 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_47
timestamp 21601
transform 1 0 644 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_26
timestamp 21601
transform -1 0 9384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_2_84
timestamp 21601
transform 1 0 5060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_2_85
timestamp 21601
transform 1 0 7636 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_2_48
timestamp 21601
transform 1 0 7636 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_2_49
timestamp 21601
transform 1 0 5060 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_2_50
timestamp 21601
transform 1 0 7636 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_51
timestamp 21601
transform 1 0 3220 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_52
timestamp 21601
transform 1 0 5796 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_53
timestamp 21601
transform 1 0 8372 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_54
timestamp 21601
transform 1 0 5796 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_55
timestamp 21601
transform 1 0 3220 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_56
timestamp 21601
transform 1 0 8372 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_57
timestamp 21601
transform 1 0 5796 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_58
timestamp 21601
transform 1 0 3220 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_59
timestamp 21601
transform 1 0 8372 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_60
timestamp 21601
transform 1 0 5796 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_61
timestamp 21601
transform 1 0 3220 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_62
timestamp 21601
transform 1 0 8372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_63
timestamp 21601
transform 1 0 5796 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_64
timestamp 21601
transform 1 0 3220 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_65
timestamp 21601
transform 1 0 8372 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_66
timestamp 21601
transform 1 0 5796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_67
timestamp 21601
transform 1 0 3220 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_68
timestamp 21601
transform 1 0 8372 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_69
timestamp 21601
transform 1 0 5796 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_70
timestamp 21601
transform 1 0 3220 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_71
timestamp 21601
transform 1 0 8372 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_72
timestamp 21601
transform 1 0 5796 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_73
timestamp 21601
transform 1 0 3220 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_74
timestamp 21601
transform 1 0 8372 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_75
timestamp 21601
transform 1 0 5796 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_76
timestamp 21601
transform 1 0 3220 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_77
timestamp 21601
transform 1 0 8372 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_78
timestamp 21601
transform 1 0 5796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_79
timestamp 21601
transform 1 0 3220 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_80
timestamp 21601
transform 1 0 8372 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_81
timestamp 21601
transform 1 0 3220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_82
timestamp 21601
transform 1 0 5796 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_83
timestamp 21601
transform 1 0 8372 0 -1 14144
box -38 -48 130 592
<< labels >>
flabel metal2 s 5078 14400 5134 15000 0 FreeSans 224 90 0 0 gpio_defaults[0]
port 0 nsew signal input
flabel metal2 s 7838 14400 7894 15000 0 FreeSans 224 90 0 0 gpio_defaults[10]
port 1 nsew signal input
flabel metal2 s 8114 14400 8170 15000 0 FreeSans 224 90 0 0 gpio_defaults[11]
port 2 nsew signal input
flabel metal2 s 8390 14400 8446 15000 0 FreeSans 224 90 0 0 gpio_defaults[12]
port 3 nsew signal input
flabel metal2 s 8666 14400 8722 15000 0 FreeSans 224 90 0 0 gpio_defaults[13]
port 4 nsew signal input
flabel metal2 s 8942 14400 8998 15000 0 FreeSans 224 90 0 0 gpio_defaults[14]
port 5 nsew signal input
flabel metal2 s 9218 14400 9274 15000 0 FreeSans 224 90 0 0 gpio_defaults[15]
port 6 nsew signal input
flabel metal2 s 5354 14400 5410 15000 0 FreeSans 224 90 0 0 gpio_defaults[1]
port 7 nsew signal input
flabel metal2 s 5630 14400 5686 15000 0 FreeSans 224 90 0 0 gpio_defaults[2]
port 8 nsew signal input
flabel metal2 s 5906 14400 5962 15000 0 FreeSans 224 90 0 0 gpio_defaults[3]
port 9 nsew signal input
flabel metal2 s 6182 14400 6238 15000 0 FreeSans 224 90 0 0 gpio_defaults[4]
port 10 nsew signal input
flabel metal2 s 6458 14400 6514 15000 0 FreeSans 224 90 0 0 gpio_defaults[5]
port 11 nsew signal input
flabel metal2 s 6734 14400 6790 15000 0 FreeSans 224 90 0 0 gpio_defaults[6]
port 12 nsew signal input
flabel metal2 s 7010 14400 7066 15000 0 FreeSans 224 90 0 0 gpio_defaults[7]
port 13 nsew signal input
flabel metal2 s 7286 14400 7342 15000 0 FreeSans 224 90 0 0 gpio_defaults[8]
port 14 nsew signal input
flabel metal2 s 7562 14400 7618 15000 0 FreeSans 224 90 0 0 gpio_defaults[9]
port 15 nsew signal input
flabel metal3 s -200 5176 400 5296 0 FreeSans 480 0 0 0 mgmt_gpio_in
port 16 nsew signal output
flabel metal3 s -200 6808 400 6928 0 FreeSans 480 0 0 0 mgmt_gpio_oeb
port 17 nsew signal input
flabel metal3 s -200 5992 400 6112 0 FreeSans 480 0 0 0 mgmt_gpio_out
port 18 nsew signal input
flabel metal3 s 9600 3272 10200 3392 0 FreeSans 480 0 0 0 pad_gpio_ana_en
port 19 nsew signal output
flabel metal3 s 9600 5720 10200 5840 0 FreeSans 480 0 0 0 pad_gpio_ana_pol
port 20 nsew signal output
flabel metal3 s 9600 7352 10200 7472 0 FreeSans 480 0 0 0 pad_gpio_ana_sel
port 21 nsew signal output
flabel metal3 s 9600 4088 10200 4208 0 FreeSans 480 0 0 0 pad_gpio_dm[0]
port 22 nsew signal output
flabel metal3 s 9600 2456 10200 2576 0 FreeSans 480 0 0 0 pad_gpio_dm[1]
port 23 nsew signal output
flabel metal3 s 9600 9800 10200 9920 0 FreeSans 480 0 0 0 pad_gpio_dm[2]
port 24 nsew signal output
flabel metal3 s 9600 10616 10200 10736 0 FreeSans 480 0 0 0 pad_gpio_holdover
port 25 nsew signal output
flabel metal3 s 9600 8984 10200 9104 0 FreeSans 480 0 0 0 pad_gpio_hys_trim
port 26 nsew signal output
flabel metal3 s 9600 13064 10200 13184 0 FreeSans 480 0 0 0 pad_gpio_ib_mode_sel
port 27 nsew signal output
flabel metal3 s 9600 824 10200 944 0 FreeSans 480 0 0 0 pad_gpio_in
port 28 nsew signal input
flabel metal3 s 9600 6536 10200 6656 0 FreeSans 480 0 0 0 pad_gpio_inenb
port 29 nsew signal output
flabel metal3 s 9600 11432 10200 11552 0 FreeSans 480 0 0 0 pad_gpio_out
port 30 nsew signal output
flabel metal3 s 9600 13880 10200 14000 0 FreeSans 480 0 0 0 pad_gpio_outenb
port 31 nsew signal output
flabel metal3 s 9600 4904 10200 5024 0 FreeSans 480 0 0 0 pad_gpio_slew_ctl[0]
port 32 nsew signal output
flabel metal3 s 9600 8168 10200 8288 0 FreeSans 480 0 0 0 pad_gpio_slew_ctl[1]
port 33 nsew signal output
flabel metal3 s 9600 1640 10200 1760 0 FreeSans 480 0 0 0 pad_gpio_slow_sel
port 34 nsew signal output
flabel metal3 s 9600 12248 10200 12368 0 FreeSans 480 0 0 0 pad_gpio_vtrip_sel
port 35 nsew signal output
flabel metal3 s -200 1912 400 2032 0 FreeSans 480 0 0 0 resetn
port 36 nsew signal input
flabel metal3 s -200 10072 400 10192 0 FreeSans 480 0 0 0 resetn_out
port 37 nsew signal output
flabel metal3 s -200 2728 400 2848 0 FreeSans 480 0 0 0 serial_clock
port 38 nsew signal input
flabel metal3 s -200 10888 400 11008 0 FreeSans 480 0 0 0 serial_clock_out
port 39 nsew signal output
flabel metal3 s -200 4360 400 4480 0 FreeSans 480 0 0 0 serial_data_in
port 40 nsew signal input
flabel metal3 s -200 12520 400 12640 0 FreeSans 480 0 0 0 serial_data_out
port 41 nsew signal output
flabel metal3 s -200 3544 400 3664 0 FreeSans 480 0 0 0 serial_load
port 42 nsew signal input
flabel metal3 s -200 11704 400 11824 0 FreeSans 480 0 0 0 serial_load_out
port 43 nsew signal output
flabel metal3 s -200 9256 400 9376 0 FreeSans 480 0 0 0 user_gpio_in
port 44 nsew signal output
flabel metal3 s -200 8440 400 8560 0 FreeSans 480 0 0 0 user_gpio_oeb
port 45 nsew signal input
flabel metal3 s -200 7624 400 7744 0 FreeSans 480 0 0 0 user_gpio_out
port 46 nsew signal input
flabel metal2 s 2544 4094 2744 14192 0 FreeSans 896 90 0 0 vccd
port 47 nsew power bidirectional
flabel metal2 s 6544 988 6744 14192 0 FreeSans 896 90 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 988 9432 1188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 4988 9432 5188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 8988 9432 9188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal3 s 596 12988 9432 13188 0 FreeSans 960 0 0 0 vccd
port 47 nsew power bidirectional
flabel metal2 s 3344 4094 3544 14192 0 FreeSans 896 90 0 0 vccd1
port 48 nsew power bidirectional
flabel metal2 s 7344 1040 7544 14192 0 FreeSans 896 90 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 1788 9432 1988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 5788 9432 5988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 9788 9432 9988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal3 s 596 13788 9432 13988 0 FreeSans 960 0 0 0 vccd1
port 48 nsew power bidirectional
flabel metal2 s 2944 4094 3144 14192 0 FreeSans 896 90 0 0 vssd
port 49 nsew ground bidirectional
flabel metal2 s 6944 1040 7144 14192 0 FreeSans 896 90 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 1388 9432 1588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 5388 9432 5588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 9388 9432 9588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal3 s 596 13388 9432 13588 0 FreeSans 960 0 0 0 vssd
port 49 nsew ground bidirectional
flabel metal2 s 3744 1040 3944 14192 0 FreeSans 896 90 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal2 s 7744 1040 7944 14192 0 FreeSans 896 90 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal3 s 596 2188 9432 2388 0 FreeSans 960 0 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal3 s 596 6188 9432 6388 0 FreeSans 960 0 0 0 vssd1
port 50 nsew ground bidirectional
flabel metal3 s 596 10188 9432 10388 0 FreeSans 960 0 0 0 vssd1
port 50 nsew ground bidirectional
rlabel metal1 5934 2720 5934 2720 0 vccd
rlabel via2 1640 1928 1640 1928 0 vccd1
rlabel metal1 5934 2176 5934 2176 0 vssd
rlabel via2 1040 2328 1040 2328 0 vssd1
rlabel metal1 3174 8432 3174 8432 0 _000_
rlabel metal2 2438 8670 2438 8670 0 _001_
rlabel metal1 5336 10778 5336 10778 0 _002_
rlabel metal1 5113 11050 5113 11050 0 _003_
rlabel metal1 7958 2414 7958 2414 0 _004_
rlabel metal1 7452 2074 7452 2074 0 _005_
rlabel metal1 8372 13158 8372 13158 0 _006_
rlabel metal1 8195 11798 8195 11798 0 _007_
rlabel metal2 5106 13022 5106 13022 0 _008_
rlabel metal1 4048 12342 4048 12342 0 _009_
rlabel metal1 7544 13498 7544 13498 0 _010_
rlabel metal2 6118 12376 6118 12376 0 _011_
rlabel metal1 8464 3706 8464 3706 0 _012_
rlabel metal1 8287 4182 8287 4182 0 _013_
rlabel metal1 7406 1734 7406 1734 0 _014_
rlabel metal1 7820 2618 7820 2618 0 _015_
rlabel metal2 8510 10812 8510 10812 0 _016_
rlabel metal1 8372 10166 8372 10166 0 _017_
rlabel metal2 6394 7242 6394 7242 0 _018_
rlabel metal2 5566 6936 5566 6936 0 _019_
rlabel metal1 7958 7344 7958 7344 0 _020_
rlabel metal1 7038 8806 7038 8806 0 _021_
rlabel metal1 8464 5882 8464 5882 0 _022_
rlabel metal1 8287 6358 8287 6358 0 _023_
rlabel metal2 8372 12716 8372 12716 0 _024_
rlabel metal1 6992 11866 6992 11866 0 _025_
rlabel metal1 8372 8058 8372 8058 0 _026_
rlabel metal2 8510 9350 8510 9350 0 _027_
rlabel metal2 5750 10404 5750 10404 0 _028_
rlabel metal1 7636 3026 7636 3026 0 _029_
rlabel metal2 6394 9758 6394 9758 0 _030_
rlabel metal1 6716 12750 6716 12750 0 _031_
rlabel metal1 6486 6222 6486 6222 0 _032_
rlabel metal1 5658 7310 5658 7310 0 _033_
rlabel metal1 4462 6766 4462 6766 0 _034_
rlabel metal1 6118 4046 6118 4046 0 _035_
rlabel metal1 3864 11322 3864 11322 0 _036_
rlabel metal2 1242 12614 1242 12614 0 _037_
rlabel metal2 6394 11934 6394 11934 0 _038_
rlabel metal1 5474 2482 5474 2482 0 _039_
rlabel metal1 3174 11186 3174 11186 0 _040_
rlabel metal1 1242 8398 1242 8398 0 _041_
rlabel metal2 2346 10506 2346 10506 0 _042_
rlabel metal1 1702 13940 1702 13940 0 gpio_defaults[0]
rlabel metal1 5428 13294 5428 13294 0 gpio_defaults[10]
rlabel metal2 3266 14076 3266 14076 0 gpio_defaults[11]
rlabel metal1 3220 13294 3220 13294 0 gpio_defaults[12]
rlabel metal2 8747 14484 8747 14484 0 gpio_defaults[13]
rlabel metal2 9147 14484 9147 14484 0 gpio_defaults[15]
rlabel metal2 5605 14484 5605 14484 0 gpio_defaults[2]
rlabel metal2 1886 13396 1886 13396 0 gpio_defaults[3]
rlabel metal2 5980 13294 5980 13294 0 gpio_defaults[4]
rlabel metal2 6072 13124 6072 13124 0 gpio_defaults[5]
rlabel metal1 5382 13838 5382 13838 0 gpio_defaults[6]
rlabel metal1 1702 13838 1702 13838 0 gpio_defaults[7]
rlabel metal2 5382 13838 5382 13838 0 gpio_defaults[8]
rlabel metal1 6578 13804 6578 13804 0 gpio_defaults[9]
rlabel metal1 2031 1530 2031 1530 0 gpio_logic1
rlabel metal1 7452 5678 7452 5678 0 gpio_slew_ctl
rlabel metal1 1656 7922 1656 7922 0 mgmt_ena
rlabel metal3 360 5236 360 5236 0 mgmt_gpio_in
rlabel metal3 774 6868 774 6868 0 mgmt_gpio_oeb
rlabel metal3 406 6052 406 6052 0 mgmt_gpio_out
rlabel metal1 2744 8908 2744 8908 0 net1
rlabel metal2 2346 8313 2346 8313 0 net10
rlabel metal1 4232 13702 4232 13702 0 net11
rlabel metal2 4094 7939 4094 7939 0 net12
rlabel metal1 1656 13158 1656 13158 0 net13
rlabel metal2 8878 13073 8878 13073 0 net14
rlabel via1 1426 7531 1426 7531 0 net15
rlabel metal2 1150 7106 1150 7106 0 net16
rlabel metal2 2990 1972 2990 1972 0 net17
rlabel metal1 1196 4794 1196 4794 0 net18
rlabel metal1 2116 7854 2116 7854 0 net19
rlabel metal1 4094 9452 4094 9452 0 net2
rlabel metal1 1150 7480 1150 7480 0 net20
rlabel metal1 1196 4454 1196 4454 0 net21
rlabel metal1 7038 1326 7038 1326 0 net22
rlabel metal2 8326 5882 8326 5882 0 net23
rlabel metal1 8422 7514 8422 7514 0 net24
rlabel metal1 8652 4250 8652 4250 0 net25
rlabel metal1 5099 3026 5099 3026 0 net26
rlabel metal2 8326 10234 8326 10234 0 net27
rlabel metal1 6946 11084 6946 11084 0 net28
rlabel via1 8974 12614 8974 12614 0 net29
rlabel metal1 3542 8840 3542 8840 0 net3
rlabel metal1 6578 13294 6578 13294 0 net30
rlabel metal1 5756 12614 5756 12614 0 net31
rlabel metal1 7406 13294 7406 13294 0 net32
rlabel metal1 3128 8058 3128 8058 0 net33
rlabel metal2 6394 5508 6394 5508 0 net34
rlabel metal1 4738 1972 4738 1972 0 net35
rlabel metal1 8468 11866 8468 11866 0 net36
rlabel metal2 966 12342 966 12342 0 net37
rlabel metal1 2484 2618 2484 2618 0 net38
rlabel metal1 5067 3434 5067 3434 0 net39
rlabel metal1 2691 10982 2691 10982 0 net4
rlabel metal2 6210 5882 6210 5882 0 net40
rlabel metal1 8694 13872 8694 13872 0 net41
rlabel metal1 3864 8466 3864 8466 0 net42
rlabel metal2 2070 7752 2070 7752 0 net43
rlabel metal3 8426 8228 8426 8228 0 net44
rlabel metal1 2254 13158 2254 13158 0 net45
rlabel metal1 6578 13906 6578 13906 0 net46
rlabel metal2 8142 7786 8142 7786 0 net47
rlabel metal1 1242 13328 1242 13328 0 net48
rlabel metal2 966 13498 966 13498 0 net49
rlabel via1 8770 8942 8770 8942 0 net5
rlabel metal1 2484 13294 2484 13294 0 net50
rlabel metal2 2162 11169 2162 11169 0 net51
rlabel metal1 3496 13906 3496 13906 0 net52
rlabel metal1 2070 13702 2070 13702 0 net53
rlabel metal1 4048 13158 4048 13158 0 net54
rlabel metal1 1518 13260 1518 13260 0 net55
rlabel metal1 3588 13770 3588 13770 0 net56
rlabel metal1 3404 12750 3404 12750 0 net57
rlabel metal1 4324 9622 4324 9622 0 net58
rlabel metal1 2392 10234 2392 10234 0 net59
rlabel via1 6026 11730 6026 11730 0 net6
rlabel metal1 6394 7378 6394 7378 0 net60
rlabel metal2 5290 4012 5290 4012 0 net61
rlabel metal2 7222 3298 7222 3298 0 net62
rlabel metal1 4876 6766 4876 6766 0 net63
rlabel metal1 5704 9894 5704 9894 0 net64
rlabel metal1 3772 11186 3772 11186 0 net65
rlabel metal1 4761 4046 4761 4046 0 net66
rlabel metal1 7084 12750 7084 12750 0 net67
rlabel metal2 5474 3026 5474 3026 0 net68
rlabel via1 5106 11526 5106 11526 0 net69
rlabel metal1 5842 13770 5842 13770 0 net7
rlabel metal2 1702 8976 1702 8976 0 net70
rlabel metal1 6348 8874 6348 8874 0 net71
rlabel metal1 6624 11662 6624 11662 0 net72
rlabel metal1 3174 13158 3174 13158 0 net8
rlabel via2 8533 12444 8533 12444 0 net9
rlabel metal3 9392 3332 9392 3332 0 pad_gpio_ana_en
rlabel metal1 8740 5746 8740 5746 0 pad_gpio_ana_pol
rlabel metal3 9024 7412 9024 7412 0 pad_gpio_ana_sel
rlabel metal3 8932 4148 8932 4148 0 pad_gpio_dm[0]
rlabel metal2 5658 2737 5658 2737 0 pad_gpio_dm[1]
rlabel via2 9622 9860 9622 9860 0 pad_gpio_dm[2]
rlabel metal3 8886 10676 8886 10676 0 pad_gpio_holdover
rlabel metal1 9108 8398 9108 8398 0 pad_gpio_hys_trim
rlabel via2 9622 13124 9622 13124 0 pad_gpio_ib_mode_sel
rlabel metal2 9062 1105 9062 1105 0 pad_gpio_in
rlabel metal3 9254 6596 9254 6596 0 pad_gpio_inenb
rlabel metal1 8372 13226 8372 13226 0 pad_gpio_out
rlabel via2 9622 13940 9622 13940 0 pad_gpio_outenb
rlabel via2 9622 4964 9622 4964 0 pad_gpio_slew_ctl[0]
rlabel via2 9622 1700 9622 1700 0 pad_gpio_slow_sel
rlabel metal2 8464 12580 8464 12580 0 pad_gpio_vtrip_sel
rlabel metal3 1196 2516 1196 2516 0 resetn
rlabel metal3 406 10132 406 10132 0 resetn_out
rlabel metal2 966 3961 966 3961 0 serial_clock
rlabel metal3 682 10948 682 10948 0 serial_clock_out
rlabel metal3 360 4420 360 4420 0 serial_data_in
rlabel metal3 866 12580 866 12580 0 serial_data_out
rlabel metal2 1058 6035 1058 6035 0 serial_load
rlabel metal3 406 11764 406 11764 0 serial_load_out
rlabel metal1 2576 5134 2576 5134 0 shift_register\[0\]
rlabel metal1 4600 4658 4600 4658 0 shift_register\[10\]
rlabel metal1 7498 1802 7498 1802 0 shift_register\[11\]
rlabel metal1 7774 6766 7774 6766 0 shift_register\[12\]
rlabel metal1 5106 9078 5106 9078 0 shift_register\[13\]
rlabel metal1 3496 10234 3496 10234 0 shift_register\[14\]
rlabel metal2 6302 11237 6302 11237 0 shift_register\[15\]
rlabel metal2 2806 9724 2806 9724 0 shift_register\[1\]
rlabel metal1 3933 10506 3933 10506 0 shift_register\[2\]
rlabel metal1 2024 12750 2024 12750 0 shift_register\[3\]
rlabel metal1 4692 11662 4692 11662 0 shift_register\[4\]
rlabel metal1 3220 7514 3220 7514 0 shift_register\[5\]
rlabel metal1 5888 6222 5888 6222 0 shift_register\[6\]
rlabel metal1 6532 5882 6532 5882 0 shift_register\[7\]
rlabel metal1 5382 3910 5382 3910 0 shift_register\[8\]
rlabel metal1 4094 3706 4094 3706 0 shift_register\[9\]
rlabel metal3 360 9316 360 9316 0 user_gpio_in
rlabel metal3 958 8500 958 8500 0 user_gpio_oeb
rlabel metal3 636 7684 636 7684 0 user_gpio_out
<< properties >>
string FIXED_BBOX 0 0 10000 14800
<< end >>
