module project_id_rom_32bit (VPWR,
    VGND,
    gpio_defaults);
 input VPWR;
 input VGND;
 output [31:0] gpio_defaults;

 wire \gpio_defaults_high[0] ;
 wire \gpio_defaults_high[10] ;
 wire \gpio_defaults_high[11] ;
 wire \gpio_defaults_high[12] ;
 wire \gpio_defaults_high[13] ;
 wire \gpio_defaults_high[14] ;
 wire \gpio_defaults_high[15] ;
 wire \gpio_defaults_high[16] ;
 wire \gpio_defaults_high[17] ;
 wire \gpio_defaults_high[18] ;
 wire \gpio_defaults_high[19] ;
 wire \gpio_defaults_high[1] ;
 wire \gpio_defaults_high[20] ;
 wire \gpio_defaults_high[21] ;
 wire \gpio_defaults_high[22] ;
 wire \gpio_defaults_high[23] ;
 wire \gpio_defaults_high[24] ;
 wire \gpio_defaults_high[25] ;
 wire \gpio_defaults_high[26] ;
 wire \gpio_defaults_high[27] ;
 wire \gpio_defaults_high[28] ;
 wire \gpio_defaults_high[29] ;
 wire \gpio_defaults_high[2] ;
 wire \gpio_defaults_high[30] ;
 wire \gpio_defaults_high[31] ;
 wire \gpio_defaults_high[3] ;
 wire \gpio_defaults_high[4] ;
 wire \gpio_defaults_high[5] ;
 wire \gpio_defaults_high[6] ;
 wire \gpio_defaults_high[7] ;
 wire \gpio_defaults_high[8] ;
 wire \gpio_defaults_high[9] ;
 wire \gpio_defaults_low[0] ;
 wire \gpio_defaults_low[10] ;
 wire \gpio_defaults_low[11] ;
 wire \gpio_defaults_low[12] ;
 wire \gpio_defaults_low[13] ;
 wire \gpio_defaults_low[14] ;
 wire \gpio_defaults_low[15] ;
 wire \gpio_defaults_low[16] ;
 wire \gpio_defaults_low[17] ;
 wire \gpio_defaults_low[18] ;
 wire \gpio_defaults_low[19] ;
 wire \gpio_defaults_low[1] ;
 wire \gpio_defaults_low[20] ;
 wire \gpio_defaults_low[21] ;
 wire \gpio_defaults_low[22] ;
 wire \gpio_defaults_low[23] ;
 wire \gpio_defaults_low[24] ;
 wire \gpio_defaults_low[25] ;
 wire \gpio_defaults_low[26] ;
 wire \gpio_defaults_low[27] ;
 wire \gpio_defaults_low[28] ;
 wire \gpio_defaults_low[29] ;
 wire \gpio_defaults_low[2] ;
 wire \gpio_defaults_low[30] ;
 wire \gpio_defaults_low[31] ;
 wire \gpio_defaults_low[3] ;
 wire \gpio_defaults_low[4] ;
 wire \gpio_defaults_low[5] ;
 wire \gpio_defaults_low[6] ;
 wire \gpio_defaults_low[7] ;
 wire \gpio_defaults_low[8] ;
 wire \gpio_defaults_low[9] ;

 sky130_fd_sc_hd__conb_1 \gpio_default_value[0]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[0] ),
    .LO(\gpio_defaults_low[0] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[10]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[10] ),
    .LO(\gpio_defaults_low[10] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[11]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[11] ),
    .LO(\gpio_defaults_low[11] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[12]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[12] ),
    .LO(\gpio_defaults_low[12] ));
 sky130_fd_sc_hd__conb_1 sky130_fd_sc_hd__conb_1_12  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[13] ),
    .LO(\gpio_defaults_low[13] ));
sky130_fd_sc_hd__conb_1 \gpio_default_value[14]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[14] ),
    .LO(\gpio_defaults_low[14] ));
sky130_fd_sc_hd__conb_1 \gpio_default_value[15]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[15] ),
    .LO(\gpio_defaults_low[15] ));
sky130_fd_sc_hd__conb_1 \gpio_default_value[16]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[16] ),
    .LO(\gpio_defaults_low[16] ));
sky130_fd_sc_hd__conb_1 \gpio_default_value[17]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[17] ),
    .LO(\gpio_defaults_low[17] ));
sky130_fd_sc_hd__conb_1 \gpio_default_value[18]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[18] ),
    .LO(\gpio_defaults_low[18] ));
sky130_fd_sc_hd__conb_1 \gpio_default_value[19]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[19] ),
    .LO(\gpio_defaults_low[19] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[1]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[1] ),
    .LO(\gpio_defaults_low[1] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[20]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[20] ),
    .LO(\gpio_defaults_low[20] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[21]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[21] ),
    .LO(\gpio_defaults_low[21] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[22]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[22] ),
    .LO(\gpio_defaults_low[22] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[23]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[23] ),
    .LO(\gpio_defaults_low[23] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[24]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[24] ),
    .LO(\gpio_defaults_low[24] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[25]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[25] ),
    .LO(\gpio_defaults_low[25] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[26]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[26] ),
    .LO(\gpio_defaults_low[26] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[27]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[27] ),
    .LO(\gpio_defaults_low[27] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[28]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[28] ),
    .LO(\gpio_defaults_low[28] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[29]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[29] ),
    .LO(\gpio_defaults_low[29] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[2]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[2] ),
    .LO(\gpio_defaults_low[2] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[30]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[30] ),
    .LO(\gpio_defaults_low[30] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[31]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[31] ),
    .LO(\gpio_defaults_low[31] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[3]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[3] ),
    .LO(\gpio_defaults_low[3] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[4]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[4] ),
    .LO(\gpio_defaults_low[4] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[5]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[5] ),
    .LO(\gpio_defaults_low[5] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[6]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[6] ),
    .LO(\gpio_defaults_low[6] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[7]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[7] ),
    .LO(\gpio_defaults_low[7] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[8]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[8] ),
    .LO(\gpio_defaults_low[8] ));
 sky130_fd_sc_hd__conb_1 \gpio_default_value[9]  (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR),
    .HI(\gpio_defaults_high[9] ),
    .LO(\gpio_defaults_low[9] ));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_4 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_3 PHY_5 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_51 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_4 FILLER_1_57 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_6 FILLER_0_3 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_15 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_27 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__decap_12 FILLER_1_39 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_9 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_29 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_0_48 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_55 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 FILLER_1_61 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 sky130_fd_sc_hd__fill_1_0 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 sky130_fd_sc_hd__fill_1_1 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__fill_1 sky130_fd_sc_hd__fill_1_2 (.VGND(VGND),
    .VNB(VGND),
    .VPB(VPWR),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_7 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_8 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_9 (.VGND(VGND),
    .VPWR(VPWR));
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_10 (.VGND(VGND),
    .VPWR(VPWR));
 
 assign gpio_defaults[0]  = \gpio_defaults_low[0] ;
 assign gpio_defaults[1]  = \gpio_defaults_low[1] ;
 assign gpio_defaults[10] = \gpio_defaults_low[10] ;
 assign gpio_defaults[11] = \gpio_defaults_low[11] ;
 assign gpio_defaults[12] = \gpio_defaults_low[12] ;
 assign gpio_defaults[13] = \gpio_defaults_low[13] ;
 assign gpio_defaults[14] = \gpio_defaults_low[14] ;
 assign gpio_defaults[15] = \gpio_defaults_low[15] ;
 assign gpio_defaults[16] = \gpio_defaults_low[16] ;
 assign gpio_defaults[17] = \gpio_defaults_low[17] ;
 assign gpio_defaults[18] = \gpio_defaults_low[18] ;
 assign gpio_defaults[19] = \gpio_defaults_low[19] ;
 assign gpio_defaults[2]  = \gpio_defaults_low[2] ;
 assign gpio_defaults[20] = \gpio_defaults_low[20] ;
 assign gpio_defaults[21] = \gpio_defaults_low[21] ;
 assign gpio_defaults[22] = \gpio_defaults_low[22] ;
 assign gpio_defaults[23] = \gpio_defaults_low[23] ;
 assign gpio_defaults[24] = \gpio_defaults_low[24] ;
 assign gpio_defaults[25] = \gpio_defaults_low[25] ;
 assign gpio_defaults[26] = \gpio_defaults_low[26] ;
 assign gpio_defaults[27] = \gpio_defaults_low[27] ;
 assign gpio_defaults[28] = \gpio_defaults_low[28] ;
 assign gpio_defaults[29] = \gpio_defaults_low[29] ;
 assign gpio_defaults[3]  = \gpio_defaults_low[3] ;
 assign gpio_defaults[30] = \gpio_defaults_low[30] ;
 assign gpio_defaults[31] = \gpio_defaults_low[31] ;
 assign gpio_defaults[4]  = \gpio_defaults_low[4] ;
 assign gpio_defaults[5]  = \gpio_defaults_low[5] ;
 assign gpio_defaults[6]  = \gpio_defaults_low[6] ;
 assign gpio_defaults[7]  = \gpio_defaults_low[7] ;
 assign gpio_defaults[8]  = \gpio_defaults_low[8] ;
 assign gpio_defaults[9]  = \gpio_defaults_low[9] ;
endmodule
