VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vccd1_tie_high
  CLASS BLOCK ;
  FOREIGN vccd1_tie_high ;
  ORIGIN 0.000 0.000 ;
  SIZE 100.000 BY 17.000 ;
  PIN HI[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 8.370 15.000 8.650 17.000 ;
    END
  END HI[0]
  PIN HI[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 17.570 15.000 17.850 17.000 ;
    END
  END HI[10]
  PIN HI[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 18.490 15.000 18.770 17.000 ;
    END
  END HI[11]
  PIN HI[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 19.410 15.000 19.690 17.000 ;
    END
  END HI[12]
  PIN HI[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 20.330 15.000 20.610 17.000 ;
    END
  END HI[13]
  PIN HI[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 21.250 15.000 21.530 17.000 ;
    END
  END HI[14]
  PIN HI[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 22.170 15.000 22.450 17.000 ;
    END
  END HI[15]
  PIN HI[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 23.090 15.000 23.370 17.000 ;
    END
  END HI[16]
  PIN HI[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 24.010 15.000 24.290 17.000 ;
    END
  END HI[17]
  PIN HI[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 24.930 15.000 25.210 17.000 ;
    END
  END HI[18]
  PIN HI[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 25.850 15.000 26.130 17.000 ;
    END
  END HI[19]
  PIN HI[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 9.290 15.000 9.570 17.000 ;
    END
  END HI[1]
  PIN HI[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 26.770 15.000 27.050 17.000 ;
    END
  END HI[20]
  PIN HI[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 27.690 15.000 27.970 17.000 ;
    END
  END HI[21]
  PIN HI[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 28.610 15.000 28.890 17.000 ;
    END
  END HI[22]
  PIN HI[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 29.530 15.000 29.810 17.000 ;
    END
  END HI[23]
  PIN HI[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 30.450 15.000 30.730 17.000 ;
    END
  END HI[24]
  PIN HI[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 31.370 15.000 31.650 17.000 ;
    END
  END HI[25]
  PIN HI[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 32.290 15.000 32.570 17.000 ;
    END
  END HI[26]
  PIN HI[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 33.210 15.000 33.490 17.000 ;
    END
  END HI[27]
  PIN HI[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 34.130 15.000 34.410 17.000 ;
    END
  END HI[28]
  PIN HI[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.050 15.000 35.330 17.000 ;
    END
  END HI[29]
  PIN HI[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 10.210 15.000 10.490 17.000 ;
    END
  END HI[2]
  PIN HI[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 35.970 15.000 36.250 17.000 ;
    END
  END HI[30]
  PIN HI[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 36.890 15.000 37.170 17.000 ;
    END
  END HI[31]
  PIN HI[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 37.810 15.000 38.090 17.000 ;
    END
  END HI[32]
  PIN HI[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 38.730 15.000 39.010 17.000 ;
    END
  END HI[33]
  PIN HI[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 39.650 15.000 39.930 17.000 ;
    END
  END HI[34]
  PIN HI[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 40.570 15.000 40.850 17.000 ;
    END
  END HI[35]
  PIN HI[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 41.490 15.000 41.770 17.000 ;
    END
  END HI[36]
  PIN HI[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 42.410 15.000 42.690 17.000 ;
    END
  END HI[37]
  PIN HI[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 43.330 15.000 43.610 17.000 ;
    END
  END HI[38]
  PIN HI[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 44.250 15.000 44.530 17.000 ;
    END
  END HI[39]
  PIN HI[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 11.130 15.000 11.410 17.000 ;
    END
  END HI[3]
  PIN HI[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 45.170 15.000 45.450 17.000 ;
    END
  END HI[40]
  PIN HI[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 46.090 15.000 46.370 17.000 ;
    END
  END HI[41]
  PIN HI[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 47.010 15.000 47.290 17.000 ;
    END
  END HI[42]
  PIN HI[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 47.930 15.000 48.210 17.000 ;
    END
  END HI[43]
  PIN HI[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 48.850 15.000 49.130 17.000 ;
    END
  END HI[44]
  PIN HI[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 49.770 15.000 50.050 17.000 ;
    END
  END HI[45]
  PIN HI[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 50.690 15.000 50.970 17.000 ;
    END
  END HI[46]
  PIN HI[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 51.610 15.000 51.890 17.000 ;
    END
  END HI[47]
  PIN HI[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 52.530 15.000 52.810 17.000 ;
    END
  END HI[48]
  PIN HI[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 53.450 15.000 53.730 17.000 ;
    END
  END HI[49]
  PIN HI[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 12.050 15.000 12.330 17.000 ;
    END
  END HI[4]
  PIN HI[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 54.370 15.000 54.650 17.000 ;
    END
  END HI[50]
  PIN HI[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 55.290 15.000 55.570 17.000 ;
    END
  END HI[51]
  PIN HI[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 56.210 15.000 56.490 17.000 ;
    END
  END HI[52]
  PIN HI[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 57.130 15.000 57.410 17.000 ;
    END
  END HI[53]
  PIN HI[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 58.050 15.000 58.330 17.000 ;
    END
  END HI[54]
  PIN HI[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 58.970 15.000 59.250 17.000 ;
    END
  END HI[55]
  PIN HI[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 59.890 15.000 60.170 17.000 ;
    END
  END HI[56]
  PIN HI[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 60.810 15.000 61.090 17.000 ;
    END
  END HI[57]
  PIN HI[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 61.730 15.000 62.010 17.000 ;
    END
  END HI[58]
  PIN HI[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 62.650 15.000 62.930 17.000 ;
    END
  END HI[59]
  PIN HI[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 12.970 15.000 13.250 17.000 ;
    END
  END HI[5]
  PIN HI[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 63.570 15.000 63.850 17.000 ;
    END
  END HI[60]
  PIN HI[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 64.490 15.000 64.770 17.000 ;
    END
  END HI[61]
  PIN HI[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 65.410 15.000 65.690 17.000 ;
    END
  END HI[62]
  PIN HI[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 66.330 15.000 66.610 17.000 ;
    END
  END HI[63]
  PIN HI[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 67.250 15.000 67.530 17.000 ;
    END
  END HI[64]
  PIN HI[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 68.170 15.000 68.450 17.000 ;
    END
  END HI[65]
  PIN HI[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 69.090 15.000 69.370 17.000 ;
    END
  END HI[66]
  PIN HI[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.010 15.000 70.290 17.000 ;
    END
  END HI[67]
  PIN HI[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.930 15.000 71.210 17.000 ;
    END
  END HI[68]
  PIN HI[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 71.850 15.000 72.130 17.000 ;
    END
  END HI[69]
  PIN HI[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 13.890 15.000 14.170 17.000 ;
    END
  END HI[6]
  PIN HI[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 72.770 15.000 73.050 17.000 ;
    END
  END HI[70]
  PIN HI[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 73.690 15.000 73.970 17.000 ;
    END
  END HI[71]
  PIN HI[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 74.610 15.000 74.890 17.000 ;
    END
  END HI[72]
  PIN HI[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 75.530 15.000 75.810 17.000 ;
    END
  END HI[73]
  PIN HI[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 76.450 15.000 76.730 17.000 ;
    END
  END HI[74]
  PIN HI[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 15.000 77.650 17.000 ;
    END
  END HI[75]
  PIN HI[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 78.290 15.000 78.570 17.000 ;
    END
  END HI[76]
  PIN HI[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 79.210 15.000 79.490 17.000 ;
    END
  END HI[77]
  PIN HI[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 80.130 15.000 80.410 17.000 ;
    END
  END HI[78]
  PIN HI[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.050 15.000 81.330 17.000 ;
    END
  END HI[79]
  PIN HI[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 14.810 15.000 15.090 17.000 ;
    END
  END HI[7]
  PIN HI[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.970 15.000 82.250 17.000 ;
    END
  END HI[80]
  PIN HI[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 82.890 15.000 83.170 17.000 ;
    END
  END HI[81]
  PIN HI[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 83.810 15.000 84.090 17.000 ;
    END
  END HI[82]
  PIN HI[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.730 15.000 85.010 17.000 ;
    END
  END HI[83]
  PIN HI[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 85.650 15.000 85.930 17.000 ;
    END
  END HI[84]
  PIN HI[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 86.570 15.000 86.850 17.000 ;
    END
  END HI[85]
  PIN HI[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 87.490 15.000 87.770 17.000 ;
    END
  END HI[86]
  PIN HI[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 88.410 15.000 88.690 17.000 ;
    END
  END HI[87]
  PIN HI[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 89.330 15.000 89.610 17.000 ;
    END
  END HI[88]
  PIN HI[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 90.250 15.000 90.530 17.000 ;
    END
  END HI[89]
  PIN HI[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 15.730 15.000 16.010 17.000 ;
    END
  END HI[8]
  PIN HI[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 91.170 15.000 91.450 17.000 ;
    END
  END HI[90]
  PIN HI[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 16.650 15.000 16.930 17.000 ;
    END
  END HI[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT 5.580 2.480 7.180 11.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 45.580 2.480 47.180 11.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 85.580 2.480 87.180 11.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.140 4.400 99.140 6.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 8.780 2.480 10.380 11.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 48.780 2.480 50.380 11.120 ;
    END
    PORT
      LAYER met2 ;
        RECT 88.780 2.480 90.380 11.120 ;
    END
    PORT
      LAYER met3 ;
        RECT 1.140 7.600 99.140 9.200 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 1.190 2.635 99.090 11.070 ;
      LAYER li1 ;
        RECT 1.380 2.635 98.900 10.965 ;
      LAYER met1 ;
        RECT 1.380 2.480 98.900 12.540 ;
      LAYER met2 ;
        RECT 7.920 14.720 8.090 15.000 ;
        RECT 8.930 14.720 9.010 15.000 ;
        RECT 9.850 14.720 9.930 15.000 ;
        RECT 10.770 14.720 10.850 15.000 ;
        RECT 11.690 14.720 11.770 15.000 ;
        RECT 12.610 14.720 12.690 15.000 ;
        RECT 13.530 14.720 13.610 15.000 ;
        RECT 14.450 14.720 14.530 15.000 ;
        RECT 15.370 14.720 15.450 15.000 ;
        RECT 16.290 14.720 16.370 15.000 ;
        RECT 17.210 14.720 17.290 15.000 ;
        RECT 18.130 14.720 18.210 15.000 ;
        RECT 19.050 14.720 19.130 15.000 ;
        RECT 19.970 14.720 20.050 15.000 ;
        RECT 20.890 14.720 20.970 15.000 ;
        RECT 21.810 14.720 21.890 15.000 ;
        RECT 22.730 14.720 22.810 15.000 ;
        RECT 23.650 14.720 23.730 15.000 ;
        RECT 24.570 14.720 24.650 15.000 ;
        RECT 25.490 14.720 25.570 15.000 ;
        RECT 26.410 14.720 26.490 15.000 ;
        RECT 27.330 14.720 27.410 15.000 ;
        RECT 28.250 14.720 28.330 15.000 ;
        RECT 29.170 14.720 29.250 15.000 ;
        RECT 30.090 14.720 30.170 15.000 ;
        RECT 31.010 14.720 31.090 15.000 ;
        RECT 31.930 14.720 32.010 15.000 ;
        RECT 32.850 14.720 32.930 15.000 ;
        RECT 33.770 14.720 33.850 15.000 ;
        RECT 34.690 14.720 34.770 15.000 ;
        RECT 35.610 14.720 35.690 15.000 ;
        RECT 36.530 14.720 36.610 15.000 ;
        RECT 37.450 14.720 37.530 15.000 ;
        RECT 38.370 14.720 38.450 15.000 ;
        RECT 39.290 14.720 39.370 15.000 ;
        RECT 40.210 14.720 40.290 15.000 ;
        RECT 41.130 14.720 41.210 15.000 ;
        RECT 42.050 14.720 42.130 15.000 ;
        RECT 42.970 14.720 43.050 15.000 ;
        RECT 43.890 14.720 43.970 15.000 ;
        RECT 44.810 14.720 44.890 15.000 ;
        RECT 45.730 14.720 45.810 15.000 ;
        RECT 46.650 14.720 46.730 15.000 ;
        RECT 47.570 14.720 47.650 15.000 ;
        RECT 48.490 14.720 48.570 15.000 ;
        RECT 49.410 14.720 49.490 15.000 ;
        RECT 50.330 14.720 50.410 15.000 ;
        RECT 51.250 14.720 51.330 15.000 ;
        RECT 52.170 14.720 52.250 15.000 ;
        RECT 53.090 14.720 53.170 15.000 ;
        RECT 54.010 14.720 54.090 15.000 ;
        RECT 54.930 14.720 55.010 15.000 ;
        RECT 55.850 14.720 55.930 15.000 ;
        RECT 56.770 14.720 56.850 15.000 ;
        RECT 57.690 14.720 57.770 15.000 ;
        RECT 58.610 14.720 58.690 15.000 ;
        RECT 59.530 14.720 59.610 15.000 ;
        RECT 60.450 14.720 60.530 15.000 ;
        RECT 61.370 14.720 61.450 15.000 ;
        RECT 62.290 14.720 62.370 15.000 ;
        RECT 63.210 14.720 63.290 15.000 ;
        RECT 64.130 14.720 64.210 15.000 ;
        RECT 65.050 14.720 65.130 15.000 ;
        RECT 65.970 14.720 66.050 15.000 ;
        RECT 66.890 14.720 66.970 15.000 ;
        RECT 67.810 14.720 67.890 15.000 ;
        RECT 68.730 14.720 68.810 15.000 ;
        RECT 69.650 14.720 69.730 15.000 ;
        RECT 70.570 14.720 70.650 15.000 ;
        RECT 71.490 14.720 71.570 15.000 ;
        RECT 72.410 14.720 72.490 15.000 ;
        RECT 73.330 14.720 73.410 15.000 ;
        RECT 74.250 14.720 74.330 15.000 ;
        RECT 75.170 14.720 75.250 15.000 ;
        RECT 76.090 14.720 76.170 15.000 ;
        RECT 77.010 14.720 77.090 15.000 ;
        RECT 77.930 14.720 78.010 15.000 ;
        RECT 78.850 14.720 78.930 15.000 ;
        RECT 79.770 14.720 79.850 15.000 ;
        RECT 80.690 14.720 80.770 15.000 ;
        RECT 81.610 14.720 81.690 15.000 ;
        RECT 82.530 14.720 82.610 15.000 ;
        RECT 83.450 14.720 83.530 15.000 ;
        RECT 84.370 14.720 84.450 15.000 ;
        RECT 85.290 14.720 85.370 15.000 ;
        RECT 86.210 14.720 86.290 15.000 ;
        RECT 87.130 14.720 87.210 15.000 ;
        RECT 88.050 14.720 88.130 15.000 ;
        RECT 88.970 14.720 89.050 15.000 ;
        RECT 89.890 14.720 89.970 15.000 ;
        RECT 90.810 14.720 90.890 15.000 ;
        RECT 91.730 14.720 96.960 15.000 ;
        RECT 7.920 11.400 96.960 14.720 ;
        RECT 7.920 3.750 8.500 11.400 ;
        RECT 10.660 3.750 45.300 11.400 ;
        RECT 47.460 3.750 48.500 11.400 ;
        RECT 50.660 3.750 85.300 11.400 ;
        RECT 87.460 3.750 88.500 11.400 ;
        RECT 90.660 3.750 96.960 11.400 ;
  END
END vccd1_tie_high
END LIBRARY

