VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO analog_ctrl_regs_APB
  CLASS BLOCK ;
  FOREIGN analog_ctrl_regs_APB ;
  ORIGIN 0.000 0.000 ;
  SIZE 1605.000 BY 105.000 ;
  PIN IRQ
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END IRQ
  PIN PADDR[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 191.450 0.000 191.730 4.000 ;
    END
  END PADDR[0]
  PIN PADDR[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 228.250 0.000 228.530 4.000 ;
    END
  END PADDR[10]
  PIN PADDR[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END PADDR[11]
  PIN PADDR[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 235.610 0.000 235.890 4.000 ;
    END
  END PADDR[12]
  PIN PADDR[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 239.290 0.000 239.570 4.000 ;
    END
  END PADDR[13]
  PIN PADDR[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END PADDR[14]
  PIN PADDR[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END PADDR[15]
  PIN PADDR[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.330 0.000 250.610 4.000 ;
    END
  END PADDR[16]
  PIN PADDR[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 254.010 0.000 254.290 4.000 ;
    END
  END PADDR[17]
  PIN PADDR[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END PADDR[18]
  PIN PADDR[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END PADDR[19]
  PIN PADDR[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 195.130 0.000 195.410 4.000 ;
    END
  END PADDR[1]
  PIN PADDR[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 0.000 265.330 4.000 ;
    END
  END PADDR[20]
  PIN PADDR[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.730 0.000 269.010 4.000 ;
    END
  END PADDR[21]
  PIN PADDR[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END PADDR[22]
  PIN PADDR[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.090 0.000 276.370 4.000 ;
    END
  END PADDR[23]
  PIN PADDR[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END PADDR[24]
  PIN PADDR[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 0.000 283.730 4.000 ;
    END
  END PADDR[25]
  PIN PADDR[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END PADDR[26]
  PIN PADDR[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 0.000 291.090 4.000 ;
    END
  END PADDR[27]
  PIN PADDR[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.490 0.000 294.770 4.000 ;
    END
  END PADDR[28]
  PIN PADDR[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END PADDR[29]
  PIN PADDR[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 198.810 0.000 199.090 4.000 ;
    END
  END PADDR[2]
  PIN PADDR[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 0.000 302.130 4.000 ;
    END
  END PADDR[30]
  PIN PADDR[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.530 0.000 305.810 4.000 ;
    END
  END PADDR[31]
  PIN PADDR[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 202.490 0.000 202.770 4.000 ;
    END
  END PADDR[3]
  PIN PADDR[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END PADDR[4]
  PIN PADDR[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 209.850 0.000 210.130 4.000 ;
    END
  END PADDR[5]
  PIN PADDR[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 213.530 0.000 213.810 4.000 ;
    END
  END PADDR[6]
  PIN PADDR[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 217.210 0.000 217.490 4.000 ;
    END
  END PADDR[7]
  PIN PADDR[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 220.890 0.000 221.170 4.000 ;
    END
  END PADDR[8]
  PIN PADDR[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END PADDR[9]
  PIN PCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.286700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END PCLK
  PIN PENABLE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END PENABLE
  PIN PRDATA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 320.250 0.000 320.530 4.000 ;
    END
  END PRDATA[0]
  PIN PRDATA[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 357.050 0.000 357.330 4.000 ;
    END
  END PRDATA[10]
  PIN PRDATA[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END PRDATA[11]
  PIN PRDATA[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 364.410 0.000 364.690 4.000 ;
    END
  END PRDATA[12]
  PIN PRDATA[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 368.090 0.000 368.370 4.000 ;
    END
  END PRDATA[13]
  PIN PRDATA[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END PRDATA[14]
  PIN PRDATA[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END PRDATA[15]
  PIN PRDATA[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 379.130 0.000 379.410 4.000 ;
    END
  END PRDATA[16]
  PIN PRDATA[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 382.810 0.000 383.090 4.000 ;
    END
  END PRDATA[17]
  PIN PRDATA[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 386.490 0.000 386.770 4.000 ;
    END
  END PRDATA[18]
  PIN PRDATA[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END PRDATA[19]
  PIN PRDATA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 323.930 0.000 324.210 4.000 ;
    END
  END PRDATA[1]
  PIN PRDATA[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 393.850 0.000 394.130 4.000 ;
    END
  END PRDATA[20]
  PIN PRDATA[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 397.530 0.000 397.810 4.000 ;
    END
  END PRDATA[21]
  PIN PRDATA[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 401.210 0.000 401.490 4.000 ;
    END
  END PRDATA[22]
  PIN PRDATA[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 404.890 0.000 405.170 4.000 ;
    END
  END PRDATA[23]
  PIN PRDATA[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END PRDATA[24]
  PIN PRDATA[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END PRDATA[25]
  PIN PRDATA[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END PRDATA[26]
  PIN PRDATA[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 419.610 0.000 419.890 4.000 ;
    END
  END PRDATA[27]
  PIN PRDATA[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END PRDATA[28]
  PIN PRDATA[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END PRDATA[29]
  PIN PRDATA[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END PRDATA[2]
  PIN PRDATA[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 430.650 0.000 430.930 4.000 ;
    END
  END PRDATA[30]
  PIN PRDATA[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 434.330 0.000 434.610 4.000 ;
    END
  END PRDATA[31]
  PIN PRDATA[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 3.107700 ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END PRDATA[3]
  PIN PRDATA[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END PRDATA[4]
  PIN PRDATA[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 338.650 0.000 338.930 4.000 ;
    END
  END PRDATA[5]
  PIN PRDATA[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END PRDATA[6]
  PIN PRDATA[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 346.010 0.000 346.290 4.000 ;
    END
  END PRDATA[7]
  PIN PRDATA[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 349.690 0.000 349.970 4.000 ;
    END
  END PRDATA[8]
  PIN PRDATA[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END PRDATA[9]
  PIN PREADY
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END PREADY
  PIN PRESETn
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END PRESETn
  PIN PSEL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 312.890 0.000 313.170 4.000 ;
    END
  END PSEL
  PIN PWDATA[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END PWDATA[0]
  PIN PWDATA[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 110.490 0.000 110.770 4.000 ;
    END
  END PWDATA[10]
  PIN PWDATA[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.177200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 114.170 0.000 114.450 4.000 ;
    END
  END PWDATA[11]
  PIN PWDATA[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.177200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 117.850 0.000 118.130 4.000 ;
    END
  END PWDATA[12]
  PIN PWDATA[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 121.530 0.000 121.810 4.000 ;
    END
  END PWDATA[13]
  PIN PWDATA[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 125.210 0.000 125.490 4.000 ;
    END
  END PWDATA[14]
  PIN PWDATA[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END PWDATA[15]
  PIN PWDATA[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 132.570 0.000 132.850 4.000 ;
    END
  END PWDATA[16]
  PIN PWDATA[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.860700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END PWDATA[17]
  PIN PWDATA[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 139.930 0.000 140.210 4.000 ;
    END
  END PWDATA[18]
  PIN PWDATA[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 143.610 0.000 143.890 4.000 ;
    END
  END PWDATA[19]
  PIN PWDATA[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END PWDATA[1]
  PIN PWDATA[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END PWDATA[20]
  PIN PWDATA[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END PWDATA[21]
  PIN PWDATA[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 154.650 0.000 154.930 4.000 ;
    END
  END PWDATA[22]
  PIN PWDATA[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 158.330 0.000 158.610 4.000 ;
    END
  END PWDATA[23]
  PIN PWDATA[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END PWDATA[24]
  PIN PWDATA[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 165.690 0.000 165.970 4.000 ;
    END
  END PWDATA[25]
  PIN PWDATA[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 169.370 0.000 169.650 4.000 ;
    END
  END PWDATA[26]
  PIN PWDATA[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END PWDATA[27]
  PIN PWDATA[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 176.730 0.000 177.010 4.000 ;
    END
  END PWDATA[28]
  PIN PWDATA[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END PWDATA[29]
  PIN PWDATA[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END PWDATA[2]
  PIN PWDATA[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END PWDATA[30]
  PIN PWDATA[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END PWDATA[31]
  PIN PWDATA[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 84.730 0.000 85.010 4.000 ;
    END
  END PWDATA[3]
  PIN PWDATA[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END PWDATA[4]
  PIN PWDATA[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END PWDATA[5]
  PIN PWDATA[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.682200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 95.770 0.000 96.050 4.000 ;
    END
  END PWDATA[6]
  PIN PWDATA[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.177200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 99.450 0.000 99.730 4.000 ;
    END
  END PWDATA[7]
  PIN PWDATA[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END PWDATA[8]
  PIN PWDATA[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.647700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 106.810 0.000 107.090 4.000 ;
    END
  END PWDATA[9]
  PIN PWRITE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.593700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 70.010 0.000 70.290 4.000 ;
    END
  END PWRITE
  PIN adc0_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 438.010 101.000 438.290 105.000 ;
    END
  END adc0_to_analog1
  PIN adc0_to_dac0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 435.250 101.000 435.530 105.000 ;
    END
  END adc0_to_dac0
  PIN adc0_to_gpio1_3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1467.490 101.000 1467.770 105.000 ;
    END
  END adc0_to_gpio1_3[0]
  PIN adc0_to_gpio1_3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1464.730 101.000 1465.010 105.000 ;
    END
  END adc0_to_gpio1_3[1]
  PIN adc0_to_gpio6_4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 117.850 101.000 118.130 105.000 ;
    END
  END adc0_to_gpio6_4[0]
  PIN adc0_to_gpio6_4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 115.090 101.000 115.370 105.000 ;
    END
  END adc0_to_gpio6_4[1]
  PIN adc0_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1185.970 101.000 1186.250 105.000 ;
    END
  END adc0_to_left_vref
  PIN adc0_to_tempsense
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1183.210 101.000 1183.490 105.000 ;
    END
  END adc0_to_tempsense
  PIN adc0_to_vbgtc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1180.450 101.000 1180.730 105.000 ;
    END
  END adc0_to_vbgtc
  PIN adc0_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1188.730 101.000 1189.010 105.000 ;
    END
  END adc0_to_voutref
  PIN adc1_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 443.530 101.000 443.810 105.000 ;
    END
  END adc1_to_analog0
  PIN adc1_to_dac1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 440.770 101.000 441.050 105.000 ;
    END
  END adc1_to_dac1
  PIN adc1_to_gpio1_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1489.570 101.000 1489.850 105.000 ;
    END
  END adc1_to_gpio1_2[0]
  PIN adc1_to_gpio1_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1486.810 101.000 1487.090 105.000 ;
    END
  END adc1_to_gpio1_2[1]
  PIN adc1_to_gpio6_5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 112.330 101.000 112.610 105.000 ;
    END
  END adc1_to_gpio6_5[0]
  PIN adc1_to_gpio6_5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 109.570 101.000 109.850 105.000 ;
    END
  END adc1_to_gpio6_5[1]
  PIN adc1_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1194.250 101.000 1194.530 105.000 ;
    END
  END adc1_to_right_vref
  PIN adc1_to_vbgsc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1191.490 101.000 1191.770 105.000 ;
    END
  END adc1_to_vbgsc
  PIN adc1_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1197.010 101.000 1197.290 105.000 ;
    END
  END adc1_to_vinref
  PIN adc_refh_to_gpio6_6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 106.810 101.000 107.090 105.000 ;
    END
  END adc_refh_to_gpio6_6[0]
  PIN adc_refh_to_gpio6_6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 104.050 101.000 104.330 105.000 ;
    END
  END adc_refh_to_gpio6_6[1]
  PIN adc_refl_to_gpio6_7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 101.290 101.000 101.570 105.000 ;
    END
  END adc_refl_to_gpio6_7[0]
  PIN adc_refl_to_gpio6_7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 98.530 101.000 98.810 105.000 ;
    END
  END adc_refl_to_gpio6_7[1]
  PIN analog0_connect[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 620.170 101.000 620.450 105.000 ;
    END
  END analog0_connect[0]
  PIN analog0_connect[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 617.410 101.000 617.690 105.000 ;
    END
  END analog0_connect[1]
  PIN analog1_connect[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 625.690 101.000 625.970 105.000 ;
    END
  END analog1_connect[0]
  PIN analog1_connect[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 622.930 101.000 623.210 105.000 ;
    END
  END analog1_connect[1]
  PIN audiodac_out_to_analog1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 432.490 101.000 432.770 105.000 ;
    END
  END audiodac_out_to_analog1[0]
  PIN audiodac_out_to_analog1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 429.730 101.000 430.010 105.000 ;
    END
  END audiodac_out_to_analog1[1]
  PIN audiodac_outb_to_analog0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 426.970 101.000 427.250 105.000 ;
    END
  END audiodac_outb_to_analog0[0]
  PIN audiodac_outb_to_analog0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 424.210 101.000 424.490 105.000 ;
    END
  END audiodac_outb_to_analog0[1]
  PIN bandgap_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 716.770 101.000 717.050 105.000 ;
    END
  END bandgap_ena
  PIN bandgap_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 675.370 101.000 675.650 105.000 ;
    END
  END bandgap_sel
  PIN bandgap_trim[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 760.930 101.000 761.210 105.000 ;
    END
  END bandgap_trim[0]
  PIN bandgap_trim[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 733.330 101.000 733.610 105.000 ;
    END
  END bandgap_trim[10]
  PIN bandgap_trim[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 730.570 101.000 730.850 105.000 ;
    END
  END bandgap_trim[11]
  PIN bandgap_trim[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 727.810 101.000 728.090 105.000 ;
    END
  END bandgap_trim[12]
  PIN bandgap_trim[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 725.050 101.000 725.330 105.000 ;
    END
  END bandgap_trim[13]
  PIN bandgap_trim[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 722.290 101.000 722.570 105.000 ;
    END
  END bandgap_trim[14]
  PIN bandgap_trim[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 719.530 101.000 719.810 105.000 ;
    END
  END bandgap_trim[15]
  PIN bandgap_trim[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 758.170 101.000 758.450 105.000 ;
    END
  END bandgap_trim[1]
  PIN bandgap_trim[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 755.410 101.000 755.690 105.000 ;
    END
  END bandgap_trim[2]
  PIN bandgap_trim[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 752.650 101.000 752.930 105.000 ;
    END
  END bandgap_trim[3]
  PIN bandgap_trim[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 749.890 101.000 750.170 105.000 ;
    END
  END bandgap_trim[4]
  PIN bandgap_trim[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 747.130 101.000 747.410 105.000 ;
    END
  END bandgap_trim[5]
  PIN bandgap_trim[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 744.370 101.000 744.650 105.000 ;
    END
  END bandgap_trim[6]
  PIN bandgap_trim[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 741.610 101.000 741.890 105.000 ;
    END
  END bandgap_trim[7]
  PIN bandgap_trim[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 738.850 101.000 739.130 105.000 ;
    END
  END bandgap_trim[8]
  PIN bandgap_trim[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 736.090 101.000 736.370 105.000 ;
    END
  END bandgap_trim[9]
  PIN brownout_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 628.450 101.000 628.730 105.000 ;
    END
  END brownout_ena
  PIN brownout_filt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 664.330 101.000 664.610 105.000 ;
    END
  END brownout_filt
  PIN brownout_isrc_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 647.770 101.000 648.050 105.000 ;
    END
  END brownout_isrc_sel
  PIN brownout_oneshot
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 650.530 101.000 650.810 105.000 ;
    END
  END brownout_oneshot
  PIN brownout_otrip[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 645.010 101.000 645.290 105.000 ;
    END
  END brownout_otrip[0]
  PIN brownout_otrip[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 642.250 101.000 642.530 105.000 ;
    END
  END brownout_otrip[1]
  PIN brownout_otrip[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 639.490 101.000 639.770 105.000 ;
    END
  END brownout_otrip[2]
  PIN brownout_rc_dis
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 656.050 101.000 656.330 105.000 ;
    END
  END brownout_rc_dis
  PIN brownout_rc_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 653.290 101.000 653.570 105.000 ;
    END
  END brownout_rc_ena
  PIN brownout_timeout
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 661.570 101.000 661.850 105.000 ;
    END
  END brownout_timeout
  PIN brownout_unfilt
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 667.090 101.000 667.370 105.000 ;
    END
  END brownout_unfilt
  PIN brownout_vtrip[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 636.730 101.000 637.010 105.000 ;
    END
  END brownout_vtrip[0]
  PIN brownout_vtrip[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 633.970 101.000 634.250 105.000 ;
    END
  END brownout_vtrip[1]
  PIN brownout_vtrip[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 631.210 101.000 631.490 105.000 ;
    END
  END brownout_vtrip[2]
  PIN brownout_vunder
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 658.810 101.000 659.090 105.000 ;
    END
  END brownout_vunder
  PIN comp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 686.410 101.000 686.690 105.000 ;
    END
  END comp_ena
  PIN comp_hyst[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 708.490 101.000 708.770 105.000 ;
    END
  END comp_hyst[0]
  PIN comp_hyst[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 705.730 101.000 706.010 105.000 ;
    END
  END comp_hyst[1]
  PIN comp_n_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1070.050 101.000 1070.330 105.000 ;
    END
  END comp_n_to_analog0
  PIN comp_n_to_dac1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1067.290 101.000 1067.570 105.000 ;
    END
  END comp_n_to_dac1
  PIN comp_n_to_gpio1_4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1461.970 101.000 1462.250 105.000 ;
    END
  END comp_n_to_gpio1_4[0]
  PIN comp_n_to_gpio1_4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1459.210 101.000 1459.490 105.000 ;
    END
  END comp_n_to_gpio1_4[1]
  PIN comp_n_to_gpio6_3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 128.890 101.000 129.170 105.000 ;
    END
  END comp_n_to_gpio6_3[0]
  PIN comp_n_to_gpio6_3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 126.130 101.000 126.410 105.000 ;
    END
  END comp_n_to_gpio6_3[1]
  PIN comp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1078.330 101.000 1078.610 105.000 ;
    END
  END comp_n_to_right_vref
  PIN comp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1072.810 101.000 1073.090 105.000 ;
    END
  END comp_n_to_sio1
  PIN comp_n_to_vbgsc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1075.570 101.000 1075.850 105.000 ;
    END
  END comp_n_to_vbgsc
  PIN comp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1081.090 101.000 1081.370 105.000 ;
    END
  END comp_n_to_vinref
  PIN comp_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 678.130 101.000 678.410 105.000 ;
    END
  END comp_out
  PIN comp_p_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1050.730 101.000 1051.010 105.000 ;
    END
  END comp_p_to_analog1
  PIN comp_p_to_dac0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1047.970 101.000 1048.250 105.000 ;
    END
  END comp_p_to_dac0
  PIN comp_p_to_gpio1_5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1456.450 101.000 1456.730 105.000 ;
    END
  END comp_p_to_gpio1_5[0]
  PIN comp_p_to_gpio1_5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1453.690 101.000 1453.970 105.000 ;
    END
  END comp_p_to_gpio1_5[1]
  PIN comp_p_to_gpio6_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 123.370 101.000 123.650 105.000 ;
    END
  END comp_p_to_gpio6_2[0]
  PIN comp_p_to_gpio6_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 120.610 101.000 120.890 105.000 ;
    END
  END comp_p_to_gpio6_2[1]
  PIN comp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1061.770 101.000 1062.050 105.000 ;
    END
  END comp_p_to_left_vref
  PIN comp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1053.490 101.000 1053.770 105.000 ;
    END
  END comp_p_to_sio0
  PIN comp_p_to_tempsense
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1059.010 101.000 1059.290 105.000 ;
    END
  END comp_p_to_tempsense
  PIN comp_p_to_vbgtc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1056.250 101.000 1056.530 105.000 ;
    END
  END comp_p_to_vbgtc
  PIN comp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1064.530 101.000 1064.810 105.000 ;
    END
  END comp_p_to_voutref
  PIN comp_trim[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 702.970 101.000 703.250 105.000 ;
    END
  END comp_trim[0]
  PIN comp_trim[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 700.210 101.000 700.490 105.000 ;
    END
  END comp_trim[1]
  PIN comp_trim[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 697.450 101.000 697.730 105.000 ;
    END
  END comp_trim[2]
  PIN comp_trim[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 694.690 101.000 694.970 105.000 ;
    END
  END comp_trim[3]
  PIN comp_trim[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 691.930 101.000 692.210 105.000 ;
    END
  END comp_trim[4]
  PIN comp_trim[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 689.170 101.000 689.450 105.000 ;
    END
  END comp_trim[5]
  PIN dac0_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 446.290 101.000 446.570 105.000 ;
    END
  END dac0_to_analog1
  PIN dac0_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1012.090 101.000 1012.370 105.000 ;
    END
  END dac0_to_user
  PIN dac1_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 449.050 101.000 449.330 105.000 ;
    END
  END dac1_to_analog0
  PIN dac1_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1014.850 101.000 1015.130 105.000 ;
    END
  END dac1_to_user
  PIN dac_refh_to_gpio1_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1495.090 101.000 1495.370 105.000 ;
    END
  END dac_refh_to_gpio1_1[0]
  PIN dac_refh_to_gpio1_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1492.330 101.000 1492.610 105.000 ;
    END
  END dac_refh_to_gpio1_1[1]
  PIN dac_refl_to_gpio1_0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1506.130 101.000 1506.410 105.000 ;
    END
  END dac_refl_to_gpio1_0[0]
  PIN dac_refl_to_gpio1_0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1503.370 101.000 1503.650 105.000 ;
    END
  END dac_refl_to_gpio1_0[1]
  PIN ibias_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 766.450 101.000 766.730 105.000 ;
    END
  END ibias_ena
  PIN ibias_ref_select
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 846.490 101.000 846.770 105.000 ;
    END
  END ibias_ref_select
  PIN ibias_snk_ena[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 843.730 101.000 844.010 105.000 ;
    END
  END ibias_snk_ena[0]
  PIN ibias_snk_ena[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 840.970 101.000 841.250 105.000 ;
    END
  END ibias_snk_ena[1]
  PIN ibias_snk_ena[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 838.210 101.000 838.490 105.000 ;
    END
  END ibias_snk_ena[2]
  PIN ibias_snk_ena[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 835.450 101.000 835.730 105.000 ;
    END
  END ibias_snk_ena[3]
  PIN ibias_src_ena[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 832.690 101.000 832.970 105.000 ;
    END
  END ibias_src_ena[0]
  PIN ibias_src_ena[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 805.090 101.000 805.370 105.000 ;
    END
  END ibias_src_ena[10]
  PIN ibias_src_ena[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 802.330 101.000 802.610 105.000 ;
    END
  END ibias_src_ena[11]
  PIN ibias_src_ena[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 799.570 101.000 799.850 105.000 ;
    END
  END ibias_src_ena[12]
  PIN ibias_src_ena[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 796.810 101.000 797.090 105.000 ;
    END
  END ibias_src_ena[13]
  PIN ibias_src_ena[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 794.050 101.000 794.330 105.000 ;
    END
  END ibias_src_ena[14]
  PIN ibias_src_ena[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 791.290 101.000 791.570 105.000 ;
    END
  END ibias_src_ena[15]
  PIN ibias_src_ena[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 788.530 101.000 788.810 105.000 ;
    END
  END ibias_src_ena[16]
  PIN ibias_src_ena[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 785.770 101.000 786.050 105.000 ;
    END
  END ibias_src_ena[17]
  PIN ibias_src_ena[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 783.010 101.000 783.290 105.000 ;
    END
  END ibias_src_ena[18]
  PIN ibias_src_ena[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 780.250 101.000 780.530 105.000 ;
    END
  END ibias_src_ena[19]
  PIN ibias_src_ena[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 829.930 101.000 830.210 105.000 ;
    END
  END ibias_src_ena[1]
  PIN ibias_src_ena[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 777.490 101.000 777.770 105.000 ;
    END
  END ibias_src_ena[20]
  PIN ibias_src_ena[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 774.730 101.000 775.010 105.000 ;
    END
  END ibias_src_ena[21]
  PIN ibias_src_ena[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 771.970 101.000 772.250 105.000 ;
    END
  END ibias_src_ena[22]
  PIN ibias_src_ena[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 769.210 101.000 769.490 105.000 ;
    END
  END ibias_src_ena[23]
  PIN ibias_src_ena[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 827.170 101.000 827.450 105.000 ;
    END
  END ibias_src_ena[2]
  PIN ibias_src_ena[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 824.410 101.000 824.690 105.000 ;
    END
  END ibias_src_ena[3]
  PIN ibias_src_ena[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 821.650 101.000 821.930 105.000 ;
    END
  END ibias_src_ena[4]
  PIN ibias_src_ena[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 818.890 101.000 819.170 105.000 ;
    END
  END ibias_src_ena[5]
  PIN ibias_src_ena[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 816.130 101.000 816.410 105.000 ;
    END
  END ibias_src_ena[6]
  PIN ibias_src_ena[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 813.370 101.000 813.650 105.000 ;
    END
  END ibias_src_ena[7]
  PIN ibias_src_ena[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 810.610 101.000 810.890 105.000 ;
    END
  END ibias_src_ena[8]
  PIN ibias_src_ena[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 807.850 101.000 808.130 105.000 ;
    END
  END ibias_src_ena[9]
  PIN ibias_test_to_gpio1_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1478.530 101.000 1478.810 105.000 ;
    END
  END ibias_test_to_gpio1_2[0]
  PIN ibias_test_to_gpio1_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1475.770 101.000 1476.050 105.000 ;
    END
  END ibias_test_to_gpio1_2[1]
  PIN idac_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 896.170 101.000 896.450 105.000 ;
    END
  END idac_ena
  PIN idac_to_gpio1_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1484.050 101.000 1484.330 105.000 ;
    END
  END idac_to_gpio1_2[0]
  PIN idac_to_gpio1_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1481.290 101.000 1481.570 105.000 ;
    END
  END idac_to_gpio1_2[1]
  PIN idac_to_gpio1_3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1473.010 101.000 1473.290 105.000 ;
    END
  END idac_to_gpio1_3[0]
  PIN idac_to_gpio1_3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1470.250 101.000 1470.530 105.000 ;
    END
  END idac_to_gpio1_3[1]
  PIN idac_value[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 893.410 101.000 893.690 105.000 ;
    END
  END idac_value[0]
  PIN idac_value[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 865.810 101.000 866.090 105.000 ;
    END
  END idac_value[10]
  PIN idac_value[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 863.050 101.000 863.330 105.000 ;
    END
  END idac_value[11]
  PIN idac_value[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 890.650 101.000 890.930 105.000 ;
    END
  END idac_value[1]
  PIN idac_value[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 887.890 101.000 888.170 105.000 ;
    END
  END idac_value[2]
  PIN idac_value[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 885.130 101.000 885.410 105.000 ;
    END
  END idac_value[3]
  PIN idac_value[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 882.370 101.000 882.650 105.000 ;
    END
  END idac_value[4]
  PIN idac_value[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 879.610 101.000 879.890 105.000 ;
    END
  END idac_value[5]
  PIN idac_value[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 876.850 101.000 877.130 105.000 ;
    END
  END idac_value[6]
  PIN idac_value[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 874.090 101.000 874.370 105.000 ;
    END
  END idac_value[7]
  PIN idac_value[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 871.330 101.000 871.610 105.000 ;
    END
  END idac_value[8]
  PIN idac_value[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 868.570 101.000 868.850 105.000 ;
    END
  END idac_value[9]
  PIN ldo_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 763.690 101.000 763.970 105.000 ;
    END
  END ldo_ena
  PIN ldo_ref_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 672.610 101.000 672.890 105.000 ;
    END
  END ldo_ref_sel
  PIN left_hgbw_opamp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 567.730 101.000 568.010 105.000 ;
    END
  END left_hgbw_opamp_ena
  PIN left_hgbw_opamp_n_to_amuxbusB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 363.490 101.000 363.770 105.000 ;
    END
  END left_hgbw_opamp_n_to_amuxbusB
  PIN left_hgbw_opamp_n_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 360.730 101.000 361.010 105.000 ;
    END
  END left_hgbw_opamp_n_to_analog1
  PIN left_hgbw_opamp_n_to_dac1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 357.970 101.000 358.250 105.000 ;
    END
  END left_hgbw_opamp_n_to_dac1
  PIN left_hgbw_opamp_n_to_gpio2_0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1439.890 101.000 1440.170 105.000 ;
    END
  END left_hgbw_opamp_n_to_gpio2_0[0]
  PIN left_hgbw_opamp_n_to_gpio2_0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1437.130 101.000 1437.410 105.000 ;
    END
  END left_hgbw_opamp_n_to_gpio2_0[1]
  PIN left_hgbw_opamp_n_to_gpio5_3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 167.530 101.000 167.810 105.000 ;
    END
  END left_hgbw_opamp_n_to_gpio5_3[0]
  PIN left_hgbw_opamp_n_to_gpio5_3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 164.770 101.000 165.050 105.000 ;
    END
  END left_hgbw_opamp_n_to_gpio5_3[1]
  PIN left_hgbw_opamp_n_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 366.250 101.000 366.530 105.000 ;
    END
  END left_hgbw_opamp_n_to_rheostat_out
  PIN left_hgbw_opamp_n_to_rheostat_tap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 369.010 101.000 369.290 105.000 ;
    END
  END left_hgbw_opamp_n_to_rheostat_tap
  PIN left_hgbw_opamp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1163.890 101.000 1164.170 105.000 ;
    END
  END left_hgbw_opamp_n_to_right_vref
  PIN left_hgbw_opamp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1158.370 101.000 1158.650 105.000 ;
    END
  END left_hgbw_opamp_n_to_sio1
  PIN left_hgbw_opamp_n_to_vbgtc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1161.130 101.000 1161.410 105.000 ;
    END
  END left_hgbw_opamp_n_to_vbgtc
  PIN left_hgbw_opamp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1166.650 101.000 1166.930 105.000 ;
    END
  END left_hgbw_opamp_n_to_vinref
  PIN left_hgbw_opamp_p_to_amuxbusA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 352.450 101.000 352.730 105.000 ;
    END
  END left_hgbw_opamp_p_to_amuxbusA
  PIN left_hgbw_opamp_p_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 349.690 101.000 349.970 105.000 ;
    END
  END left_hgbw_opamp_p_to_analog0
  PIN left_hgbw_opamp_p_to_dac0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 346.930 101.000 347.210 105.000 ;
    END
  END left_hgbw_opamp_p_to_dac0
  PIN left_hgbw_opamp_p_to_gpio2_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1434.370 101.000 1434.650 105.000 ;
    END
  END left_hgbw_opamp_p_to_gpio2_1[0]
  PIN left_hgbw_opamp_p_to_gpio2_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1431.610 101.000 1431.890 105.000 ;
    END
  END left_hgbw_opamp_p_to_gpio2_1[1]
  PIN left_hgbw_opamp_p_to_gpio5_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 173.050 101.000 173.330 105.000 ;
    END
  END left_hgbw_opamp_p_to_gpio5_2[0]
  PIN left_hgbw_opamp_p_to_gpio5_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 170.290 101.000 170.570 105.000 ;
    END
  END left_hgbw_opamp_p_to_gpio5_2[1]
  PIN left_hgbw_opamp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1144.570 101.000 1144.850 105.000 ;
    END
  END left_hgbw_opamp_p_to_left_vref
  PIN left_hgbw_opamp_p_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 355.210 101.000 355.490 105.000 ;
    END
  END left_hgbw_opamp_p_to_rheostat_out
  PIN left_hgbw_opamp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1139.050 101.000 1139.330 105.000 ;
    END
  END left_hgbw_opamp_p_to_sio0
  PIN left_hgbw_opamp_p_to_tempsense
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1141.810 101.000 1142.090 105.000 ;
    END
  END left_hgbw_opamp_p_to_tempsense
  PIN left_hgbw_opamp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1147.330 101.000 1147.610 105.000 ;
    END
  END left_hgbw_opamp_p_to_voutref
  PIN left_hgbw_opamp_to_adc0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 333.130 101.000 333.410 105.000 ;
    END
  END left_hgbw_opamp_to_adc0[0]
  PIN left_hgbw_opamp_to_adc0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 330.370 101.000 330.650 105.000 ;
    END
  END left_hgbw_opamp_to_adc0[1]
  PIN left_hgbw_opamp_to_amuxbusB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 344.170 101.000 344.450 105.000 ;
    END
  END left_hgbw_opamp_to_amuxbusB[0]
  PIN left_hgbw_opamp_to_amuxbusB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 341.410 101.000 341.690 105.000 ;
    END
  END left_hgbw_opamp_to_amuxbusB[1]
  PIN left_hgbw_opamp_to_analog1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 338.650 101.000 338.930 105.000 ;
    END
  END left_hgbw_opamp_to_analog1[0]
  PIN left_hgbw_opamp_to_analog1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 335.890 101.000 336.170 105.000 ;
    END
  END left_hgbw_opamp_to_analog1[1]
  PIN left_hgbw_opamp_to_comp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 327.610 101.000 327.890 105.000 ;
    END
  END left_hgbw_opamp_to_comp_p[0]
  PIN left_hgbw_opamp_to_comp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 324.850 101.000 325.130 105.000 ;
    END
  END left_hgbw_opamp_to_comp_p[1]
  PIN left_hgbw_opamp_to_gpio3_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1387.450 101.000 1387.730 105.000 ;
    END
  END left_hgbw_opamp_to_gpio3_1[0]
  PIN left_hgbw_opamp_to_gpio3_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1384.690 101.000 1384.970 105.000 ;
    END
  END left_hgbw_opamp_to_gpio3_1[1]
  PIN left_hgbw_opamp_to_gpio3_5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1365.370 101.000 1365.650 105.000 ;
    END
  END left_hgbw_opamp_to_gpio3_5[0]
  PIN left_hgbw_opamp_to_gpio3_5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1362.610 101.000 1362.890 105.000 ;
    END
  END left_hgbw_opamp_to_gpio3_5[1]
  PIN left_hgbw_opamp_to_gpio4_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 222.730 101.000 223.010 105.000 ;
    END
  END left_hgbw_opamp_to_gpio4_1[0]
  PIN left_hgbw_opamp_to_gpio4_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 219.970 101.000 220.250 105.000 ;
    END
  END left_hgbw_opamp_to_gpio4_1[1]
  PIN left_hgbw_opamp_to_gpio4_5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 200.650 101.000 200.930 105.000 ;
    END
  END left_hgbw_opamp_to_gpio4_5[0]
  PIN left_hgbw_opamp_to_gpio4_5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 197.890 101.000 198.170 105.000 ;
    END
  END left_hgbw_opamp_to_gpio4_5[1]
  PIN left_hgbw_opamp_to_ulpcomp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 322.090 101.000 322.370 105.000 ;
    END
  END left_hgbw_opamp_to_ulpcomp_p[0]
  PIN left_hgbw_opamp_to_ulpcomp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 319.330 101.000 319.610 105.000 ;
    END
  END left_hgbw_opamp_to_ulpcomp_p[1]
  PIN left_instramp_G1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 551.170 101.000 551.450 105.000 ;
    END
  END left_instramp_G1[0]
  PIN left_instramp_G1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 548.410 101.000 548.690 105.000 ;
    END
  END left_instramp_G1[1]
  PIN left_instramp_G1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 545.650 101.000 545.930 105.000 ;
    END
  END left_instramp_G1[2]
  PIN left_instramp_G1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 542.890 101.000 543.170 105.000 ;
    END
  END left_instramp_G1[3]
  PIN left_instramp_G1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 540.130 101.000 540.410 105.000 ;
    END
  END left_instramp_G1[4]
  PIN left_instramp_G2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 564.970 101.000 565.250 105.000 ;
    END
  END left_instramp_G2[0]
  PIN left_instramp_G2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 562.210 101.000 562.490 105.000 ;
    END
  END left_instramp_G2[1]
  PIN left_instramp_G2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 559.450 101.000 559.730 105.000 ;
    END
  END left_instramp_G2[2]
  PIN left_instramp_G2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 556.690 101.000 556.970 105.000 ;
    END
  END left_instramp_G2[3]
  PIN left_instramp_G2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 553.930 101.000 554.210 105.000 ;
    END
  END left_instramp_G2[4]
  PIN left_instramp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 537.370 101.000 537.650 105.000 ;
    END
  END left_instramp_ena
  PIN left_instramp_n_to_amuxbusB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 261.370 101.000 261.650 105.000 ;
    END
  END left_instramp_n_to_amuxbusB
  PIN left_instramp_n_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 258.610 101.000 258.890 105.000 ;
    END
  END left_instramp_n_to_analog1
  PIN left_instramp_n_to_gpio5_7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 145.450 101.000 145.730 105.000 ;
    END
  END left_instramp_n_to_gpio5_7[0]
  PIN left_instramp_n_to_gpio5_7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 142.690 101.000 142.970 105.000 ;
    END
  END left_instramp_n_to_gpio5_7[1]
  PIN left_instramp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1122.490 101.000 1122.770 105.000 ;
    END
  END left_instramp_n_to_right_vref
  PIN left_instramp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1119.730 101.000 1120.010 105.000 ;
    END
  END left_instramp_n_to_sio1
  PIN left_instramp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1125.250 101.000 1125.530 105.000 ;
    END
  END left_instramp_n_to_vinref
  PIN left_instramp_p_to_amuxbusA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 316.570 101.000 316.850 105.000 ;
    END
  END left_instramp_p_to_amuxbusA
  PIN left_instramp_p_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 313.810 101.000 314.090 105.000 ;
    END
  END left_instramp_p_to_analog0
  PIN left_instramp_p_to_gpio5_6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 150.970 101.000 151.250 105.000 ;
    END
  END left_instramp_p_to_gpio5_6[0]
  PIN left_instramp_p_to_gpio5_6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 148.210 101.000 148.490 105.000 ;
    END
  END left_instramp_p_to_gpio5_6[1]
  PIN left_instramp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1133.530 101.000 1133.810 105.000 ;
    END
  END left_instramp_p_to_left_vref
  PIN left_instramp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1128.010 101.000 1128.290 105.000 ;
    END
  END left_instramp_p_to_sio0
  PIN left_instramp_p_to_tempsense
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1130.770 101.000 1131.050 105.000 ;
    END
  END left_instramp_p_to_tempsense
  PIN left_instramp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1136.290 101.000 1136.570 105.000 ;
    END
  END left_instramp_p_to_voutref
  PIN left_instramp_to_adc0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 244.810 101.000 245.090 105.000 ;
    END
  END left_instramp_to_adc0[0]
  PIN left_instramp_to_adc0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 242.050 101.000 242.330 105.000 ;
    END
  END left_instramp_to_adc0[1]
  PIN left_instramp_to_amuxbusB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 255.850 101.000 256.130 105.000 ;
    END
  END left_instramp_to_amuxbusB[0]
  PIN left_instramp_to_amuxbusB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 253.090 101.000 253.370 105.000 ;
    END
  END left_instramp_to_amuxbusB[1]
  PIN left_instramp_to_analog1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 250.330 101.000 250.610 105.000 ;
    END
  END left_instramp_to_analog1[0]
  PIN left_instramp_to_analog1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 247.570 101.000 247.850 105.000 ;
    END
  END left_instramp_to_analog1[1]
  PIN left_instramp_to_comp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 239.290 101.000 239.570 105.000 ;
    END
  END left_instramp_to_comp_p[0]
  PIN left_instramp_to_comp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 236.530 101.000 236.810 105.000 ;
    END
  END left_instramp_to_comp_p[1]
  PIN left_instramp_to_gpio4_4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 206.170 101.000 206.450 105.000 ;
    END
  END left_instramp_to_gpio4_4[0]
  PIN left_instramp_to_gpio4_4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 203.410 101.000 203.690 105.000 ;
    END
  END left_instramp_to_gpio4_4[1]
  PIN left_instramp_to_ulpcomp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 233.770 101.000 234.050 105.000 ;
    END
  END left_instramp_to_ulpcomp_p[0]
  PIN left_instramp_to_ulpcomp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 231.010 101.000 231.290 105.000 ;
    END
  END left_instramp_to_ulpcomp_p[1]
  PIN left_lp_opamp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 570.490 101.000 570.770 105.000 ;
    END
  END left_lp_opamp_ena
  PIN left_lp_opamp_n_to_amuxbusB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 415.930 101.000 416.210 105.000 ;
    END
  END left_lp_opamp_n_to_amuxbusB
  PIN left_lp_opamp_n_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 413.170 101.000 413.450 105.000 ;
    END
  END left_lp_opamp_n_to_analog1
  PIN left_lp_opamp_n_to_dac1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 410.410 101.000 410.690 105.000 ;
    END
  END left_lp_opamp_n_to_dac1
  PIN left_lp_opamp_n_to_gpio5_5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 156.490 101.000 156.770 105.000 ;
    END
  END left_lp_opamp_n_to_gpio5_5[0]
  PIN left_lp_opamp_n_to_gpio5_5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 153.730 101.000 154.010 105.000 ;
    END
  END left_lp_opamp_n_to_gpio5_5[1]
  PIN left_lp_opamp_n_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 418.690 101.000 418.970 105.000 ;
    END
  END left_lp_opamp_n_to_rheostat_out
  PIN left_lp_opamp_n_to_rheostat_tap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 421.450 101.000 421.730 105.000 ;
    END
  END left_lp_opamp_n_to_rheostat_tap
  PIN left_lp_opamp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1174.930 101.000 1175.210 105.000 ;
    END
  END left_lp_opamp_n_to_right_vref
  PIN left_lp_opamp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1169.410 101.000 1169.690 105.000 ;
    END
  END left_lp_opamp_n_to_sio1
  PIN left_lp_opamp_n_to_vbgsc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1172.170 101.000 1172.450 105.000 ;
    END
  END left_lp_opamp_n_to_vbgsc
  PIN left_lp_opamp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1177.690 101.000 1177.970 105.000 ;
    END
  END left_lp_opamp_n_to_vinref
  PIN left_lp_opamp_p_to_amuxbusA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 404.890 101.000 405.170 105.000 ;
    END
  END left_lp_opamp_p_to_amuxbusA
  PIN left_lp_opamp_p_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 402.130 101.000 402.410 105.000 ;
    END
  END left_lp_opamp_p_to_analog0
  PIN left_lp_opamp_p_to_dac0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 399.370 101.000 399.650 105.000 ;
    END
  END left_lp_opamp_p_to_dac0
  PIN left_lp_opamp_p_to_gpio5_4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 162.010 101.000 162.290 105.000 ;
    END
  END left_lp_opamp_p_to_gpio5_4[0]
  PIN left_lp_opamp_p_to_gpio5_4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 159.250 101.000 159.530 105.000 ;
    END
  END left_lp_opamp_p_to_gpio5_4[1]
  PIN left_lp_opamp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1152.850 101.000 1153.130 105.000 ;
    END
  END left_lp_opamp_p_to_left_vref
  PIN left_lp_opamp_p_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 407.650 101.000 407.930 105.000 ;
    END
  END left_lp_opamp_p_to_rheostat_out
  PIN left_lp_opamp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1150.090 101.000 1150.370 105.000 ;
    END
  END left_lp_opamp_p_to_sio0
  PIN left_lp_opamp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1155.610 101.000 1155.890 105.000 ;
    END
  END left_lp_opamp_p_to_voutref
  PIN left_lp_opamp_to_adc1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 385.570 101.000 385.850 105.000 ;
    END
  END left_lp_opamp_to_adc1[0]
  PIN left_lp_opamp_to_adc1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 382.810 101.000 383.090 105.000 ;
    END
  END left_lp_opamp_to_adc1[1]
  PIN left_lp_opamp_to_amuxbusA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 396.610 101.000 396.890 105.000 ;
    END
  END left_lp_opamp_to_amuxbusA[0]
  PIN left_lp_opamp_to_amuxbusA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 393.850 101.000 394.130 105.000 ;
    END
  END left_lp_opamp_to_amuxbusA[1]
  PIN left_lp_opamp_to_analog0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 391.090 101.000 391.370 105.000 ;
    END
  END left_lp_opamp_to_analog0[0]
  PIN left_lp_opamp_to_analog0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 388.330 101.000 388.610 105.000 ;
    END
  END left_lp_opamp_to_analog0[1]
  PIN left_lp_opamp_to_comp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 380.050 101.000 380.330 105.000 ;
    END
  END left_lp_opamp_to_comp_n[0]
  PIN left_lp_opamp_to_comp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 377.290 101.000 377.570 105.000 ;
    END
  END left_lp_opamp_to_comp_n[1]
  PIN left_lp_opamp_to_gpio3_4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1370.890 101.000 1371.170 105.000 ;
    END
  END left_lp_opamp_to_gpio3_4[0]
  PIN left_lp_opamp_to_gpio3_4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1368.130 101.000 1368.410 105.000 ;
    END
  END left_lp_opamp_to_gpio3_4[1]
  PIN left_lp_opamp_to_gpio4_0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 228.250 101.000 228.530 105.000 ;
    END
  END left_lp_opamp_to_gpio4_0[0]
  PIN left_lp_opamp_to_gpio4_0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 225.490 101.000 225.770 105.000 ;
    END
  END left_lp_opamp_to_gpio4_0[1]
  PIN left_lp_opamp_to_ulpcomp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 374.530 101.000 374.810 105.000 ;
    END
  END left_lp_opamp_to_ulpcomp_n[0]
  PIN left_lp_opamp_to_ulpcomp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 371.770 101.000 372.050 105.000 ;
    END
  END left_lp_opamp_to_ulpcomp_n[1]
  PIN left_rheostat1_b[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 592.570 101.000 592.850 105.000 ;
    END
  END left_rheostat1_b[0]
  PIN left_rheostat1_b[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 589.810 101.000 590.090 105.000 ;
    END
  END left_rheostat1_b[1]
  PIN left_rheostat1_b[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 587.050 101.000 587.330 105.000 ;
    END
  END left_rheostat1_b[2]
  PIN left_rheostat1_b[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 584.290 101.000 584.570 105.000 ;
    END
  END left_rheostat1_b[3]
  PIN left_rheostat1_b[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 581.530 101.000 581.810 105.000 ;
    END
  END left_rheostat1_b[4]
  PIN left_rheostat1_b[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 578.770 101.000 579.050 105.000 ;
    END
  END left_rheostat1_b[5]
  PIN left_rheostat1_b[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 576.010 101.000 576.290 105.000 ;
    END
  END left_rheostat1_b[6]
  PIN left_rheostat1_b[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 573.250 101.000 573.530 105.000 ;
    END
  END left_rheostat1_b[7]
  PIN left_rheostat2_b[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 614.650 101.000 614.930 105.000 ;
    END
  END left_rheostat2_b[0]
  PIN left_rheostat2_b[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 611.890 101.000 612.170 105.000 ;
    END
  END left_rheostat2_b[1]
  PIN left_rheostat2_b[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 609.130 101.000 609.410 105.000 ;
    END
  END left_rheostat2_b[2]
  PIN left_rheostat2_b[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 606.370 101.000 606.650 105.000 ;
    END
  END left_rheostat2_b[3]
  PIN left_rheostat2_b[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 603.610 101.000 603.890 105.000 ;
    END
  END left_rheostat2_b[4]
  PIN left_rheostat2_b[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 600.850 101.000 601.130 105.000 ;
    END
  END left_rheostat2_b[5]
  PIN left_rheostat2_b[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 598.090 101.000 598.370 105.000 ;
    END
  END left_rheostat2_b[6]
  PIN left_rheostat2_b[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 595.330 101.000 595.610 105.000 ;
    END
  END left_rheostat2_b[7]
  PIN left_vref_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1023.130 101.000 1023.410 105.000 ;
    END
  END left_vref_to_user
  PIN overvoltage_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 849.250 101.000 849.530 105.000 ;
    END
  END overvoltage_ena
  PIN overvoltage_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 683.650 101.000 683.930 105.000 ;
    END
  END overvoltage_out
  PIN overvoltage_trim[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 860.290 101.000 860.570 105.000 ;
    END
  END overvoltage_trim[0]
  PIN overvoltage_trim[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 857.530 101.000 857.810 105.000 ;
    END
  END overvoltage_trim[1]
  PIN overvoltage_trim[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 854.770 101.000 855.050 105.000 ;
    END
  END overvoltage_trim[2]
  PIN overvoltage_trim[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 852.010 101.000 852.290 105.000 ;
    END
  END overvoltage_trim[3]
  PIN rdac0_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 465.610 101.000 465.890 105.000 ;
    END
  END rdac0_ena
  PIN rdac0_value[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 498.730 101.000 499.010 105.000 ;
    END
  END rdac0_value[0]
  PIN rdac0_value[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 471.130 101.000 471.410 105.000 ;
    END
  END rdac0_value[10]
  PIN rdac0_value[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 468.370 101.000 468.650 105.000 ;
    END
  END rdac0_value[11]
  PIN rdac0_value[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 495.970 101.000 496.250 105.000 ;
    END
  END rdac0_value[1]
  PIN rdac0_value[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 493.210 101.000 493.490 105.000 ;
    END
  END rdac0_value[2]
  PIN rdac0_value[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 490.450 101.000 490.730 105.000 ;
    END
  END rdac0_value[3]
  PIN rdac0_value[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 487.690 101.000 487.970 105.000 ;
    END
  END rdac0_value[4]
  PIN rdac0_value[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 484.930 101.000 485.210 105.000 ;
    END
  END rdac0_value[5]
  PIN rdac0_value[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 482.170 101.000 482.450 105.000 ;
    END
  END rdac0_value[6]
  PIN rdac0_value[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 479.410 101.000 479.690 105.000 ;
    END
  END rdac0_value[7]
  PIN rdac0_value[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 476.650 101.000 476.930 105.000 ;
    END
  END rdac0_value[8]
  PIN rdac0_value[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 473.890 101.000 474.170 105.000 ;
    END
  END rdac0_value[9]
  PIN rdac1_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 501.490 101.000 501.770 105.000 ;
    END
  END rdac1_ena
  PIN rdac1_value[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 534.610 101.000 534.890 105.000 ;
    END
  END rdac1_value[0]
  PIN rdac1_value[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 507.010 101.000 507.290 105.000 ;
    END
  END rdac1_value[10]
  PIN rdac1_value[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 504.250 101.000 504.530 105.000 ;
    END
  END rdac1_value[11]
  PIN rdac1_value[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 531.850 101.000 532.130 105.000 ;
    END
  END rdac1_value[1]
  PIN rdac1_value[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 529.090 101.000 529.370 105.000 ;
    END
  END rdac1_value[2]
  PIN rdac1_value[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 526.330 101.000 526.610 105.000 ;
    END
  END rdac1_value[3]
  PIN rdac1_value[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 523.570 101.000 523.850 105.000 ;
    END
  END rdac1_value[4]
  PIN rdac1_value[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 520.810 101.000 521.090 105.000 ;
    END
  END rdac1_value[5]
  PIN rdac1_value[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 518.050 101.000 518.330 105.000 ;
    END
  END rdac1_value[6]
  PIN rdac1_value[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 515.290 101.000 515.570 105.000 ;
    END
  END rdac1_value[7]
  PIN rdac1_value[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 512.530 101.000 512.810 105.000 ;
    END
  END rdac1_value[8]
  PIN rdac1_value[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 509.770 101.000 510.050 105.000 ;
    END
  END rdac1_value[9]
  PIN right_hgbw_opamp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 929.290 101.000 929.570 105.000 ;
    END
  END right_hgbw_opamp_ena
  PIN right_hgbw_opamp_n_to_amuxbusB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1293.610 101.000 1293.890 105.000 ;
    END
  END right_hgbw_opamp_n_to_amuxbusB
  PIN right_hgbw_opamp_n_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1290.850 101.000 1291.130 105.000 ;
    END
  END right_hgbw_opamp_n_to_analog1
  PIN right_hgbw_opamp_n_to_dac1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1288.090 101.000 1288.370 105.000 ;
    END
  END right_hgbw_opamp_n_to_dac1
  PIN right_hgbw_opamp_n_to_gpio2_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1428.850 101.000 1429.130 105.000 ;
    END
  END right_hgbw_opamp_n_to_gpio2_2[0]
  PIN right_hgbw_opamp_n_to_gpio2_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1426.090 101.000 1426.370 105.000 ;
    END
  END right_hgbw_opamp_n_to_gpio2_2[1]
  PIN right_hgbw_opamp_n_to_gpio5_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 178.570 101.000 178.850 105.000 ;
    END
  END right_hgbw_opamp_n_to_gpio5_1[0]
  PIN right_hgbw_opamp_n_to_gpio5_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 175.810 101.000 176.090 105.000 ;
    END
  END right_hgbw_opamp_n_to_gpio5_1[1]
  PIN right_hgbw_opamp_n_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1296.370 101.000 1296.650 105.000 ;
    END
  END right_hgbw_opamp_n_to_rheostat_out
  PIN right_hgbw_opamp_n_to_rheostat_tap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1299.130 101.000 1299.410 105.000 ;
    END
  END right_hgbw_opamp_n_to_rheostat_tap
  PIN right_hgbw_opamp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1307.410 101.000 1307.690 105.000 ;
    END
  END right_hgbw_opamp_n_to_right_vref
  PIN right_hgbw_opamp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1301.890 101.000 1302.170 105.000 ;
    END
  END right_hgbw_opamp_n_to_sio1
  PIN right_hgbw_opamp_n_to_vbgsc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1304.650 101.000 1304.930 105.000 ;
    END
  END right_hgbw_opamp_n_to_vbgsc
  PIN right_hgbw_opamp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1310.170 101.000 1310.450 105.000 ;
    END
  END right_hgbw_opamp_n_to_vinref
  PIN right_hgbw_opamp_p_to_amuxbusA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1274.290 101.000 1274.570 105.000 ;
    END
  END right_hgbw_opamp_p_to_amuxbusA
  PIN right_hgbw_opamp_p_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1271.530 101.000 1271.810 105.000 ;
    END
  END right_hgbw_opamp_p_to_analog0
  PIN right_hgbw_opamp_p_to_dac0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1268.770 101.000 1269.050 105.000 ;
    END
  END right_hgbw_opamp_p_to_dac0
  PIN right_hgbw_opamp_p_to_gpio2_3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1423.330 101.000 1423.610 105.000 ;
    END
  END right_hgbw_opamp_p_to_gpio2_3[0]
  PIN right_hgbw_opamp_p_to_gpio2_3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1420.570 101.000 1420.850 105.000 ;
    END
  END right_hgbw_opamp_p_to_gpio2_3[1]
  PIN right_hgbw_opamp_p_to_gpio5_0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 184.090 101.000 184.370 105.000 ;
    END
  END right_hgbw_opamp_p_to_gpio5_0[0]
  PIN right_hgbw_opamp_p_to_gpio5_0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 181.330 101.000 181.610 105.000 ;
    END
  END right_hgbw_opamp_p_to_gpio5_0[1]
  PIN right_hgbw_opamp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1282.570 101.000 1282.850 105.000 ;
    END
  END right_hgbw_opamp_p_to_left_vref
  PIN right_hgbw_opamp_p_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1277.050 101.000 1277.330 105.000 ;
    END
  END right_hgbw_opamp_p_to_rheostat_out
  PIN right_hgbw_opamp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1279.810 101.000 1280.090 105.000 ;
    END
  END right_hgbw_opamp_p_to_sio0
  PIN right_hgbw_opamp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1285.330 101.000 1285.610 105.000 ;
    END
  END right_hgbw_opamp_p_to_voutref
  PIN right_hgbw_opamp_to_adc1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 294.490 101.000 294.770 105.000 ;
    END
  END right_hgbw_opamp_to_adc1[0]
  PIN right_hgbw_opamp_to_adc1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 291.730 101.000 292.010 105.000 ;
    END
  END right_hgbw_opamp_to_adc1[1]
  PIN right_hgbw_opamp_to_amuxbusA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1266.010 101.000 1266.290 105.000 ;
    END
  END right_hgbw_opamp_to_amuxbusA[0]
  PIN right_hgbw_opamp_to_amuxbusA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1263.250 101.000 1263.530 105.000 ;
    END
  END right_hgbw_opamp_to_amuxbusA[1]
  PIN right_hgbw_opamp_to_analog0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1260.490 101.000 1260.770 105.000 ;
    END
  END right_hgbw_opamp_to_analog0[0]
  PIN right_hgbw_opamp_to_analog0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1257.730 101.000 1258.010 105.000 ;
    END
  END right_hgbw_opamp_to_analog0[1]
  PIN right_hgbw_opamp_to_comp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 288.970 101.000 289.250 105.000 ;
    END
  END right_hgbw_opamp_to_comp_n[0]
  PIN right_hgbw_opamp_to_comp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 286.210 101.000 286.490 105.000 ;
    END
  END right_hgbw_opamp_to_comp_n[1]
  PIN right_hgbw_opamp_to_gpio3_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1381.930 101.000 1382.210 105.000 ;
    END
  END right_hgbw_opamp_to_gpio3_2[0]
  PIN right_hgbw_opamp_to_gpio3_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1379.170 101.000 1379.450 105.000 ;
    END
  END right_hgbw_opamp_to_gpio3_2[1]
  PIN right_hgbw_opamp_to_gpio3_6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1359.850 101.000 1360.130 105.000 ;
    END
  END right_hgbw_opamp_to_gpio3_6[0]
  PIN right_hgbw_opamp_to_gpio3_6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1357.090 101.000 1357.370 105.000 ;
    END
  END right_hgbw_opamp_to_gpio3_6[1]
  PIN right_hgbw_opamp_to_gpio4_2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 217.210 101.000 217.490 105.000 ;
    END
  END right_hgbw_opamp_to_gpio4_2[0]
  PIN right_hgbw_opamp_to_gpio4_2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 214.450 101.000 214.730 105.000 ;
    END
  END right_hgbw_opamp_to_gpio4_2[1]
  PIN right_hgbw_opamp_to_gpio4_6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 195.130 101.000 195.410 105.000 ;
    END
  END right_hgbw_opamp_to_gpio4_6[0]
  PIN right_hgbw_opamp_to_gpio4_6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 192.370 101.000 192.650 105.000 ;
    END
  END right_hgbw_opamp_to_gpio4_6[1]
  PIN right_hgbw_opamp_to_ulpcomp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 283.450 101.000 283.730 105.000 ;
    END
  END right_hgbw_opamp_to_ulpcomp_n[0]
  PIN right_hgbw_opamp_to_ulpcomp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 280.690 101.000 280.970 105.000 ;
    END
  END right_hgbw_opamp_to_ulpcomp_n[1]
  PIN right_instramp_G1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 912.730 101.000 913.010 105.000 ;
    END
  END right_instramp_G1[0]
  PIN right_instramp_G1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 909.970 101.000 910.250 105.000 ;
    END
  END right_instramp_G1[1]
  PIN right_instramp_G1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 907.210 101.000 907.490 105.000 ;
    END
  END right_instramp_G1[2]
  PIN right_instramp_G1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 904.450 101.000 904.730 105.000 ;
    END
  END right_instramp_G1[3]
  PIN right_instramp_G1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 901.690 101.000 901.970 105.000 ;
    END
  END right_instramp_G1[4]
  PIN right_instramp_G2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 926.530 101.000 926.810 105.000 ;
    END
  END right_instramp_G2[0]
  PIN right_instramp_G2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 923.770 101.000 924.050 105.000 ;
    END
  END right_instramp_G2[1]
  PIN right_instramp_G2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 921.010 101.000 921.290 105.000 ;
    END
  END right_instramp_G2[2]
  PIN right_instramp_G2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 918.250 101.000 918.530 105.000 ;
    END
  END right_instramp_G2[3]
  PIN right_instramp_G2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 915.490 101.000 915.770 105.000 ;
    END
  END right_instramp_G2[4]
  PIN right_instramp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 898.930 101.000 899.210 105.000 ;
    END
  END right_instramp_ena
  PIN right_instramp_n_to_amuxbusB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1326.730 101.000 1327.010 105.000 ;
    END
  END right_instramp_n_to_amuxbusB
  PIN right_instramp_n_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1323.970 101.000 1324.250 105.000 ;
    END
  END right_instramp_n_to_analog1
  PIN right_instramp_n_to_gpio2_6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1406.770 101.000 1407.050 105.000 ;
    END
  END right_instramp_n_to_gpio2_6[0]
  PIN right_instramp_n_to_gpio2_6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1404.010 101.000 1404.290 105.000 ;
    END
  END right_instramp_n_to_gpio2_6[1]
  PIN right_instramp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1332.250 101.000 1332.530 105.000 ;
    END
  END right_instramp_n_to_right_vref
  PIN right_instramp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1329.490 101.000 1329.770 105.000 ;
    END
  END right_instramp_n_to_sio1
  PIN right_instramp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1335.010 101.000 1335.290 105.000 ;
    END
  END right_instramp_n_to_vinref
  PIN right_instramp_p_to_amuxbusA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1340.530 101.000 1340.810 105.000 ;
    END
  END right_instramp_p_to_amuxbusA
  PIN right_instramp_p_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1337.770 101.000 1338.050 105.000 ;
    END
  END right_instramp_p_to_analog0
  PIN right_instramp_p_to_gpio2_7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1401.250 101.000 1401.530 105.000 ;
    END
  END right_instramp_p_to_gpio2_7[0]
  PIN right_instramp_p_to_gpio2_7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1398.490 101.000 1398.770 105.000 ;
    END
  END right_instramp_p_to_gpio2_7[1]
  PIN right_instramp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1346.050 101.000 1346.330 105.000 ;
    END
  END right_instramp_p_to_left_vref
  PIN right_instramp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1395.730 101.000 1396.010 105.000 ;
    END
  END right_instramp_p_to_sio0
  PIN right_instramp_p_to_tempsense
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1343.290 101.000 1343.570 105.000 ;
    END
  END right_instramp_p_to_tempsense
  PIN right_instramp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1348.810 101.000 1349.090 105.000 ;
    END
  END right_instramp_p_to_voutref
  PIN right_instramp_to_adc1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 311.050 101.000 311.330 105.000 ;
    END
  END right_instramp_to_adc1[0]
  PIN right_instramp_to_adc1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 308.290 101.000 308.570 105.000 ;
    END
  END right_instramp_to_adc1[1]
  PIN right_instramp_to_amuxbusA[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1321.210 101.000 1321.490 105.000 ;
    END
  END right_instramp_to_amuxbusA[0]
  PIN right_instramp_to_amuxbusA[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1318.450 101.000 1318.730 105.000 ;
    END
  END right_instramp_to_amuxbusA[1]
  PIN right_instramp_to_analog0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1315.690 101.000 1315.970 105.000 ;
    END
  END right_instramp_to_analog0[0]
  PIN right_instramp_to_analog0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1312.930 101.000 1313.210 105.000 ;
    END
  END right_instramp_to_analog0[1]
  PIN right_instramp_to_comp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 305.530 101.000 305.810 105.000 ;
    END
  END right_instramp_to_comp_n[0]
  PIN right_instramp_to_comp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 302.770 101.000 303.050 105.000 ;
    END
  END right_instramp_to_comp_n[1]
  PIN right_instramp_to_gpio3_0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1392.970 101.000 1393.250 105.000 ;
    END
  END right_instramp_to_gpio3_0[0]
  PIN right_instramp_to_gpio3_0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1390.210 101.000 1390.490 105.000 ;
    END
  END right_instramp_to_gpio3_0[1]
  PIN right_instramp_to_ulpcomp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 300.010 101.000 300.290 105.000 ;
    END
  END right_instramp_to_ulpcomp_n[0]
  PIN right_instramp_to_ulpcomp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 297.250 101.000 297.530 105.000 ;
    END
  END right_instramp_to_ulpcomp_n[1]
  PIN right_lp_opamp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 932.050 101.000 932.330 105.000 ;
    END
  END right_lp_opamp_ena
  PIN right_lp_opamp_n_to_amuxbusB
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1238.410 101.000 1238.690 105.000 ;
    END
  END right_lp_opamp_n_to_amuxbusB
  PIN right_lp_opamp_n_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1235.650 101.000 1235.930 105.000 ;
    END
  END right_lp_opamp_n_to_analog1
  PIN right_lp_opamp_n_to_dac1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1232.890 101.000 1233.170 105.000 ;
    END
  END right_lp_opamp_n_to_dac1
  PIN right_lp_opamp_n_to_gpio2_4[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1417.810 101.000 1418.090 105.000 ;
    END
  END right_lp_opamp_n_to_gpio2_4[0]
  PIN right_lp_opamp_n_to_gpio2_4[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1415.050 101.000 1415.330 105.000 ;
    END
  END right_lp_opamp_n_to_gpio2_4[1]
  PIN right_lp_opamp_n_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 101.000 1241.450 105.000 ;
    END
  END right_lp_opamp_n_to_rheostat_out
  PIN right_lp_opamp_n_to_rheostat_tap
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1243.930 101.000 1244.210 105.000 ;
    END
  END right_lp_opamp_n_to_rheostat_tap
  PIN right_lp_opamp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1252.210 101.000 1252.490 105.000 ;
    END
  END right_lp_opamp_n_to_right_vref
  PIN right_lp_opamp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1246.690 101.000 1246.970 105.000 ;
    END
  END right_lp_opamp_n_to_sio1
  PIN right_lp_opamp_n_to_vbgtc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1249.450 101.000 1249.730 105.000 ;
    END
  END right_lp_opamp_n_to_vbgtc
  PIN right_lp_opamp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1254.970 101.000 1255.250 105.000 ;
    END
  END right_lp_opamp_n_to_vinref
  PIN right_lp_opamp_p_to_amuxbusA
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1216.330 101.000 1216.610 105.000 ;
    END
  END right_lp_opamp_p_to_amuxbusA
  PIN right_lp_opamp_p_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1213.570 101.000 1213.850 105.000 ;
    END
  END right_lp_opamp_p_to_analog0
  PIN right_lp_opamp_p_to_dac0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1210.810 101.000 1211.090 105.000 ;
    END
  END right_lp_opamp_p_to_dac0
  PIN right_lp_opamp_p_to_gpio2_5[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1412.290 101.000 1412.570 105.000 ;
    END
  END right_lp_opamp_p_to_gpio2_5[0]
  PIN right_lp_opamp_p_to_gpio2_5[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1409.530 101.000 1409.810 105.000 ;
    END
  END right_lp_opamp_p_to_gpio2_5[1]
  PIN right_lp_opamp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1227.370 101.000 1227.650 105.000 ;
    END
  END right_lp_opamp_p_to_left_vref
  PIN right_lp_opamp_p_to_rheostat_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1219.090 101.000 1219.370 105.000 ;
    END
  END right_lp_opamp_p_to_rheostat_out
  PIN right_lp_opamp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1221.850 101.000 1222.130 105.000 ;
    END
  END right_lp_opamp_p_to_sio0
  PIN right_lp_opamp_p_to_tempsense
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1224.610 101.000 1224.890 105.000 ;
    END
  END right_lp_opamp_p_to_tempsense
  PIN right_lp_opamp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1230.130 101.000 1230.410 105.000 ;
    END
  END right_lp_opamp_p_to_voutref
  PIN right_lp_opamp_to_adc0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 277.930 101.000 278.210 105.000 ;
    END
  END right_lp_opamp_to_adc0[0]
  PIN right_lp_opamp_to_adc0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 275.170 101.000 275.450 105.000 ;
    END
  END right_lp_opamp_to_adc0[1]
  PIN right_lp_opamp_to_amuxbusB[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1208.050 101.000 1208.330 105.000 ;
    END
  END right_lp_opamp_to_amuxbusB[0]
  PIN right_lp_opamp_to_amuxbusB[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1205.290 101.000 1205.570 105.000 ;
    END
  END right_lp_opamp_to_amuxbusB[1]
  PIN right_lp_opamp_to_analog1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1202.530 101.000 1202.810 105.000 ;
    END
  END right_lp_opamp_to_analog1[0]
  PIN right_lp_opamp_to_analog1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1199.770 101.000 1200.050 105.000 ;
    END
  END right_lp_opamp_to_analog1[1]
  PIN right_lp_opamp_to_comp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 272.410 101.000 272.690 105.000 ;
    END
  END right_lp_opamp_to_comp_p[0]
  PIN right_lp_opamp_to_comp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 269.650 101.000 269.930 105.000 ;
    END
  END right_lp_opamp_to_comp_p[1]
  PIN right_lp_opamp_to_gpio3_3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1376.410 101.000 1376.690 105.000 ;
    END
  END right_lp_opamp_to_gpio3_3[0]
  PIN right_lp_opamp_to_gpio3_3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1373.650 101.000 1373.930 105.000 ;
    END
  END right_lp_opamp_to_gpio3_3[1]
  PIN right_lp_opamp_to_gpio3_7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1354.330 101.000 1354.610 105.000 ;
    END
  END right_lp_opamp_to_gpio3_7[0]
  PIN right_lp_opamp_to_gpio3_7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1351.570 101.000 1351.850 105.000 ;
    END
  END right_lp_opamp_to_gpio3_7[1]
  PIN right_lp_opamp_to_gpio4_3[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 211.690 101.000 211.970 105.000 ;
    END
  END right_lp_opamp_to_gpio4_3[0]
  PIN right_lp_opamp_to_gpio4_3[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 208.930 101.000 209.210 105.000 ;
    END
  END right_lp_opamp_to_gpio4_3[1]
  PIN right_lp_opamp_to_gpio4_7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 189.610 101.000 189.890 105.000 ;
    END
  END right_lp_opamp_to_gpio4_7[0]
  PIN right_lp_opamp_to_gpio4_7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 186.850 101.000 187.130 105.000 ;
    END
  END right_lp_opamp_to_gpio4_7[1]
  PIN right_lp_opamp_to_ulpcomp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 266.890 101.000 267.170 105.000 ;
    END
  END right_lp_opamp_to_ulpcomp_p[0]
  PIN right_lp_opamp_to_ulpcomp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 264.130 101.000 264.410 105.000 ;
    END
  END right_lp_opamp_to_ulpcomp_p[1]
  PIN right_rheostat1_b[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 954.130 101.000 954.410 105.000 ;
    END
  END right_rheostat1_b[0]
  PIN right_rheostat1_b[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 951.370 101.000 951.650 105.000 ;
    END
  END right_rheostat1_b[1]
  PIN right_rheostat1_b[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 948.610 101.000 948.890 105.000 ;
    END
  END right_rheostat1_b[2]
  PIN right_rheostat1_b[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 945.850 101.000 946.130 105.000 ;
    END
  END right_rheostat1_b[3]
  PIN right_rheostat1_b[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 943.090 101.000 943.370 105.000 ;
    END
  END right_rheostat1_b[4]
  PIN right_rheostat1_b[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 940.330 101.000 940.610 105.000 ;
    END
  END right_rheostat1_b[5]
  PIN right_rheostat1_b[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 937.570 101.000 937.850 105.000 ;
    END
  END right_rheostat1_b[6]
  PIN right_rheostat1_b[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 934.810 101.000 935.090 105.000 ;
    END
  END right_rheostat1_b[7]
  PIN right_rheostat2_b[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 976.210 101.000 976.490 105.000 ;
    END
  END right_rheostat2_b[0]
  PIN right_rheostat2_b[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 973.450 101.000 973.730 105.000 ;
    END
  END right_rheostat2_b[1]
  PIN right_rheostat2_b[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 970.690 101.000 970.970 105.000 ;
    END
  END right_rheostat2_b[2]
  PIN right_rheostat2_b[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 967.930 101.000 968.210 105.000 ;
    END
  END right_rheostat2_b[3]
  PIN right_rheostat2_b[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 965.170 101.000 965.450 105.000 ;
    END
  END right_rheostat2_b[4]
  PIN right_rheostat2_b[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 962.410 101.000 962.690 105.000 ;
    END
  END right_rheostat2_b[5]
  PIN right_rheostat2_b[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 959.650 101.000 959.930 105.000 ;
    END
  END right_rheostat2_b[6]
  PIN right_rheostat2_b[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 956.890 101.000 957.170 105.000 ;
    END
  END right_rheostat2_b[7]
  PIN right_vref_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1020.370 101.000 1020.650 105.000 ;
    END
  END right_vref_to_user
  PIN sio0_connect[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1039.690 101.000 1039.970 105.000 ;
    END
  END sio0_connect[0]
  PIN sio0_connect[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1036.930 101.000 1037.210 105.000 ;
    END
  END sio0_connect[1]
  PIN sio1_connect[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1045.210 101.000 1045.490 105.000 ;
    END
  END sio1_connect[0]
  PIN sio1_connect[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1042.450 101.000 1042.730 105.000 ;
    END
  END sio1_connect[1]
  PIN tempsense_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 462.850 101.000 463.130 105.000 ;
    END
  END tempsense_ena
  PIN tempsense_sel
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 669.850 101.000 670.130 105.000 ;
    END
  END tempsense_sel
  PIN tempsense_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1017.610 101.000 1017.890 105.000 ;
    END
  END tempsense_to_user
  PIN ulpcomp_clk
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 714.010 101.000 714.290 105.000 ;
    END
  END ulpcomp_clk
  PIN ulpcomp_ena
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 711.250 101.000 711.530 105.000 ;
    END
  END ulpcomp_ena
  PIN ulpcomp_n_to_analog0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1105.930 101.000 1106.210 105.000 ;
    END
  END ulpcomp_n_to_analog0
  PIN ulpcomp_n_to_dac1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1103.170 101.000 1103.450 105.000 ;
    END
  END ulpcomp_n_to_dac1
  PIN ulpcomp_n_to_gpio1_6[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1450.930 101.000 1451.210 105.000 ;
    END
  END ulpcomp_n_to_gpio1_6[0]
  PIN ulpcomp_n_to_gpio1_6[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1448.170 101.000 1448.450 105.000 ;
    END
  END ulpcomp_n_to_gpio1_6[1]
  PIN ulpcomp_n_to_gpio6_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 134.410 101.000 134.690 105.000 ;
    END
  END ulpcomp_n_to_gpio6_1[0]
  PIN ulpcomp_n_to_gpio6_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 131.650 101.000 131.930 105.000 ;
    END
  END ulpcomp_n_to_gpio6_1[1]
  PIN ulpcomp_n_to_right_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1114.210 101.000 1114.490 105.000 ;
    END
  END ulpcomp_n_to_right_vref
  PIN ulpcomp_n_to_sio1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1108.690 101.000 1108.970 105.000 ;
    END
  END ulpcomp_n_to_sio1
  PIN ulpcomp_n_to_vbgsc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1111.450 101.000 1111.730 105.000 ;
    END
  END ulpcomp_n_to_vbgsc
  PIN ulpcomp_n_to_vinref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1116.970 101.000 1117.250 105.000 ;
    END
  END ulpcomp_n_to_vinref
  PIN ulpcomp_out
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 680.890 101.000 681.170 105.000 ;
    END
  END ulpcomp_out
  PIN ulpcomp_p_to_analog1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1086.610 101.000 1086.890 105.000 ;
    END
  END ulpcomp_p_to_analog1
  PIN ulpcomp_p_to_dac0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1083.850 101.000 1084.130 105.000 ;
    END
  END ulpcomp_p_to_dac0
  PIN ulpcomp_p_to_gpio1_7[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1445.410 101.000 1445.690 105.000 ;
    END
  END ulpcomp_p_to_gpio1_7[0]
  PIN ulpcomp_p_to_gpio1_7[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1442.650 101.000 1442.930 105.000 ;
    END
  END ulpcomp_p_to_gpio1_7[1]
  PIN ulpcomp_p_to_gpio6_0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 139.930 101.000 140.210 105.000 ;
    END
  END ulpcomp_p_to_gpio6_0[0]
  PIN ulpcomp_p_to_gpio6_0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 137.170 101.000 137.450 105.000 ;
    END
  END ulpcomp_p_to_gpio6_0[1]
  PIN ulpcomp_p_to_left_vref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1097.650 101.000 1097.930 105.000 ;
    END
  END ulpcomp_p_to_left_vref
  PIN ulpcomp_p_to_sio0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1089.370 101.000 1089.650 105.000 ;
    END
  END ulpcomp_p_to_sio0
  PIN ulpcomp_p_to_tempsense
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1094.890 101.000 1095.170 105.000 ;
    END
  END ulpcomp_p_to_tempsense
  PIN ulpcomp_p_to_vbgtc
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1092.130 101.000 1092.410 105.000 ;
    END
  END ulpcomp_p_to_vbgtc
  PIN ulpcomp_p_to_voutref
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1100.410 101.000 1100.690 105.000 ;
    END
  END ulpcomp_p_to_voutref
  PIN user_to_adc0[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1003.810 101.000 1004.090 105.000 ;
    END
  END user_to_adc0[0]
  PIN user_to_adc0[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1001.050 101.000 1001.330 105.000 ;
    END
  END user_to_adc0[1]
  PIN user_to_adc1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1009.330 101.000 1009.610 105.000 ;
    END
  END user_to_adc1[0]
  PIN user_to_adc1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1006.570 101.000 1006.850 105.000 ;
    END
  END user_to_adc1[1]
  PIN user_to_comp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 981.730 101.000 982.010 105.000 ;
    END
  END user_to_comp_n[0]
  PIN user_to_comp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 978.970 101.000 979.250 105.000 ;
    END
  END user_to_comp_n[1]
  PIN user_to_comp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 987.250 101.000 987.530 105.000 ;
    END
  END user_to_comp_p[0]
  PIN user_to_comp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 984.490 101.000 984.770 105.000 ;
    END
  END user_to_comp_p[1]
  PIN user_to_ulpcomp_n[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 992.770 101.000 993.050 105.000 ;
    END
  END user_to_ulpcomp_n[0]
  PIN user_to_ulpcomp_n[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 990.010 101.000 990.290 105.000 ;
    END
  END user_to_ulpcomp_n[1]
  PIN user_to_ulpcomp_p[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 998.290 101.000 998.570 105.000 ;
    END
  END user_to_ulpcomp_p[0]
  PIN user_to_ulpcomp_p[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 995.530 101.000 995.810 105.000 ;
    END
  END user_to_ulpcomp_p[1]
  PIN vbg_test_to_gpio1_1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1500.610 101.000 1500.890 105.000 ;
    END
  END vbg_test_to_gpio1_1[0]
  PIN vbg_test_to_gpio1_1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1497.850 101.000 1498.130 105.000 ;
    END
  END vbg_test_to_gpio1_1[1]
  PIN vbgsc_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1034.170 101.000 1034.450 105.000 ;
    END
  END vbgsc_to_user
  PIN vbgtc_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1031.410 101.000 1031.690 105.000 ;
    END
  END vbgtc_to_user
  PIN vccd0
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 20.580 5.200 22.180 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.180 5.200 175.780 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 327.780 5.200 329.380 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.380 5.200 482.980 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 634.980 5.200 636.580 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 788.580 5.200 790.180 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.180 5.200 943.780 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.380 5.200 1250.980 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1402.980 5.200 1404.580 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1556.580 5.200 1558.180 98.160 ;
    END
  END vccd0
  PIN vccd1_pwr_good
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 454.570 101.000 454.850 105.000 ;
    END
  END vccd1_pwr_good
  PIN vccd2_pwr_good
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 460.090 101.000 460.370 105.000 ;
    END
  END vccd2_pwr_good
  PIN vdda1_pwr_good
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.631200 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 451.810 101.000 452.090 105.000 ;
    END
  END vdda1_pwr_good
  PIN vdda2_pwr_good
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.929700 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 457.330 101.000 457.610 105.000 ;
    END
  END vdda2_pwr_good
  PIN vinref_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1025.890 101.000 1026.170 105.000 ;
    END
  END vinref_to_user
  PIN voutref_to_user
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.434700 ;
    ANTENNADIFFAREA 2.025100 ;
    PORT
      LAYER met2 ;
        RECT 1028.650 101.000 1028.930 105.000 ;
    END
  END voutref_to_user
  PIN vssd0
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 23.880 5.200 25.480 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.480 5.200 179.080 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 331.080 5.200 332.680 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 484.680 5.200 486.280 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.280 5.200 639.880 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 791.880 5.200 793.480 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 945.480 5.200 947.080 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1252.680 5.200 1254.280 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1406.280 5.200 1407.880 98.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 1559.880 5.200 1561.480 98.160 ;
    END
  END vssd0
  OBS
      LAYER nwell ;
        RECT 4.870 5.355 1600.070 98.005 ;
      LAYER li1 ;
        RECT 5.060 5.355 1599.880 98.005 ;
      LAYER met1 ;
        RECT 5.060 0.040 1599.880 104.960 ;
      LAYER met2 ;
        RECT 20.610 100.720 98.250 104.710 ;
        RECT 99.090 100.720 101.010 104.710 ;
        RECT 101.850 100.720 103.770 104.710 ;
        RECT 104.610 100.720 106.530 104.710 ;
        RECT 107.370 100.720 109.290 104.710 ;
        RECT 110.130 100.720 112.050 104.710 ;
        RECT 112.890 100.720 114.810 104.710 ;
        RECT 115.650 100.720 117.570 104.710 ;
        RECT 118.410 100.720 120.330 104.710 ;
        RECT 121.170 100.720 123.090 104.710 ;
        RECT 123.930 100.720 125.850 104.710 ;
        RECT 126.690 100.720 128.610 104.710 ;
        RECT 129.450 100.720 131.370 104.710 ;
        RECT 132.210 100.720 134.130 104.710 ;
        RECT 134.970 100.720 136.890 104.710 ;
        RECT 137.730 100.720 139.650 104.710 ;
        RECT 140.490 100.720 142.410 104.710 ;
        RECT 143.250 100.720 145.170 104.710 ;
        RECT 146.010 100.720 147.930 104.710 ;
        RECT 148.770 100.720 150.690 104.710 ;
        RECT 151.530 100.720 153.450 104.710 ;
        RECT 154.290 100.720 156.210 104.710 ;
        RECT 157.050 100.720 158.970 104.710 ;
        RECT 159.810 100.720 161.730 104.710 ;
        RECT 162.570 100.720 164.490 104.710 ;
        RECT 165.330 100.720 167.250 104.710 ;
        RECT 168.090 100.720 170.010 104.710 ;
        RECT 170.850 100.720 172.770 104.710 ;
        RECT 173.610 100.720 175.530 104.710 ;
        RECT 176.370 100.720 178.290 104.710 ;
        RECT 179.130 100.720 181.050 104.710 ;
        RECT 181.890 100.720 183.810 104.710 ;
        RECT 184.650 100.720 186.570 104.710 ;
        RECT 187.410 100.720 189.330 104.710 ;
        RECT 190.170 100.720 192.090 104.710 ;
        RECT 192.930 100.720 194.850 104.710 ;
        RECT 195.690 100.720 197.610 104.710 ;
        RECT 198.450 100.720 200.370 104.710 ;
        RECT 201.210 100.720 203.130 104.710 ;
        RECT 203.970 100.720 205.890 104.710 ;
        RECT 206.730 100.720 208.650 104.710 ;
        RECT 209.490 100.720 211.410 104.710 ;
        RECT 212.250 100.720 214.170 104.710 ;
        RECT 215.010 100.720 216.930 104.710 ;
        RECT 217.770 100.720 219.690 104.710 ;
        RECT 220.530 100.720 222.450 104.710 ;
        RECT 223.290 100.720 225.210 104.710 ;
        RECT 226.050 100.720 227.970 104.710 ;
        RECT 228.810 100.720 230.730 104.710 ;
        RECT 231.570 100.720 233.490 104.710 ;
        RECT 234.330 100.720 236.250 104.710 ;
        RECT 237.090 100.720 239.010 104.710 ;
        RECT 239.850 100.720 241.770 104.710 ;
        RECT 242.610 100.720 244.530 104.710 ;
        RECT 245.370 100.720 247.290 104.710 ;
        RECT 248.130 100.720 250.050 104.710 ;
        RECT 250.890 100.720 252.810 104.710 ;
        RECT 253.650 100.720 255.570 104.710 ;
        RECT 256.410 100.720 258.330 104.710 ;
        RECT 259.170 100.720 261.090 104.710 ;
        RECT 261.930 100.720 263.850 104.710 ;
        RECT 264.690 100.720 266.610 104.710 ;
        RECT 267.450 100.720 269.370 104.710 ;
        RECT 270.210 100.720 272.130 104.710 ;
        RECT 272.970 100.720 274.890 104.710 ;
        RECT 275.730 100.720 277.650 104.710 ;
        RECT 278.490 100.720 280.410 104.710 ;
        RECT 281.250 100.720 283.170 104.710 ;
        RECT 284.010 100.720 285.930 104.710 ;
        RECT 286.770 100.720 288.690 104.710 ;
        RECT 289.530 100.720 291.450 104.710 ;
        RECT 292.290 100.720 294.210 104.710 ;
        RECT 295.050 100.720 296.970 104.710 ;
        RECT 297.810 100.720 299.730 104.710 ;
        RECT 300.570 100.720 302.490 104.710 ;
        RECT 303.330 100.720 305.250 104.710 ;
        RECT 306.090 100.720 308.010 104.710 ;
        RECT 308.850 100.720 310.770 104.710 ;
        RECT 311.610 100.720 313.530 104.710 ;
        RECT 314.370 100.720 316.290 104.710 ;
        RECT 317.130 100.720 319.050 104.710 ;
        RECT 319.890 100.720 321.810 104.710 ;
        RECT 322.650 100.720 324.570 104.710 ;
        RECT 325.410 100.720 327.330 104.710 ;
        RECT 328.170 100.720 330.090 104.710 ;
        RECT 330.930 100.720 332.850 104.710 ;
        RECT 333.690 100.720 335.610 104.710 ;
        RECT 336.450 100.720 338.370 104.710 ;
        RECT 339.210 100.720 341.130 104.710 ;
        RECT 341.970 100.720 343.890 104.710 ;
        RECT 344.730 100.720 346.650 104.710 ;
        RECT 347.490 100.720 349.410 104.710 ;
        RECT 350.250 100.720 352.170 104.710 ;
        RECT 353.010 100.720 354.930 104.710 ;
        RECT 355.770 100.720 357.690 104.710 ;
        RECT 358.530 100.720 360.450 104.710 ;
        RECT 361.290 100.720 363.210 104.710 ;
        RECT 364.050 100.720 365.970 104.710 ;
        RECT 366.810 100.720 368.730 104.710 ;
        RECT 369.570 100.720 371.490 104.710 ;
        RECT 372.330 100.720 374.250 104.710 ;
        RECT 375.090 100.720 377.010 104.710 ;
        RECT 377.850 100.720 379.770 104.710 ;
        RECT 380.610 100.720 382.530 104.710 ;
        RECT 383.370 100.720 385.290 104.710 ;
        RECT 386.130 100.720 388.050 104.710 ;
        RECT 388.890 100.720 390.810 104.710 ;
        RECT 391.650 100.720 393.570 104.710 ;
        RECT 394.410 100.720 396.330 104.710 ;
        RECT 397.170 100.720 399.090 104.710 ;
        RECT 399.930 100.720 401.850 104.710 ;
        RECT 402.690 100.720 404.610 104.710 ;
        RECT 405.450 100.720 407.370 104.710 ;
        RECT 408.210 100.720 410.130 104.710 ;
        RECT 410.970 100.720 412.890 104.710 ;
        RECT 413.730 100.720 415.650 104.710 ;
        RECT 416.490 100.720 418.410 104.710 ;
        RECT 419.250 100.720 421.170 104.710 ;
        RECT 422.010 100.720 423.930 104.710 ;
        RECT 424.770 100.720 426.690 104.710 ;
        RECT 427.530 100.720 429.450 104.710 ;
        RECT 430.290 100.720 432.210 104.710 ;
        RECT 433.050 100.720 434.970 104.710 ;
        RECT 435.810 100.720 437.730 104.710 ;
        RECT 438.570 100.720 440.490 104.710 ;
        RECT 441.330 100.720 443.250 104.710 ;
        RECT 444.090 100.720 446.010 104.710 ;
        RECT 446.850 100.720 448.770 104.710 ;
        RECT 449.610 100.720 451.530 104.710 ;
        RECT 452.370 100.720 454.290 104.710 ;
        RECT 455.130 100.720 457.050 104.710 ;
        RECT 457.890 100.720 459.810 104.710 ;
        RECT 460.650 100.720 462.570 104.710 ;
        RECT 463.410 100.720 465.330 104.710 ;
        RECT 466.170 100.720 468.090 104.710 ;
        RECT 468.930 100.720 470.850 104.710 ;
        RECT 471.690 100.720 473.610 104.710 ;
        RECT 474.450 100.720 476.370 104.710 ;
        RECT 477.210 100.720 479.130 104.710 ;
        RECT 479.970 100.720 481.890 104.710 ;
        RECT 482.730 100.720 484.650 104.710 ;
        RECT 485.490 100.720 487.410 104.710 ;
        RECT 488.250 100.720 490.170 104.710 ;
        RECT 491.010 100.720 492.930 104.710 ;
        RECT 493.770 100.720 495.690 104.710 ;
        RECT 496.530 100.720 498.450 104.710 ;
        RECT 499.290 100.720 501.210 104.710 ;
        RECT 502.050 100.720 503.970 104.710 ;
        RECT 504.810 100.720 506.730 104.710 ;
        RECT 507.570 100.720 509.490 104.710 ;
        RECT 510.330 100.720 512.250 104.710 ;
        RECT 513.090 100.720 515.010 104.710 ;
        RECT 515.850 100.720 517.770 104.710 ;
        RECT 518.610 100.720 520.530 104.710 ;
        RECT 521.370 100.720 523.290 104.710 ;
        RECT 524.130 100.720 526.050 104.710 ;
        RECT 526.890 100.720 528.810 104.710 ;
        RECT 529.650 100.720 531.570 104.710 ;
        RECT 532.410 100.720 534.330 104.710 ;
        RECT 535.170 100.720 537.090 104.710 ;
        RECT 537.930 100.720 539.850 104.710 ;
        RECT 540.690 100.720 542.610 104.710 ;
        RECT 543.450 100.720 545.370 104.710 ;
        RECT 546.210 100.720 548.130 104.710 ;
        RECT 548.970 100.720 550.890 104.710 ;
        RECT 551.730 100.720 553.650 104.710 ;
        RECT 554.490 100.720 556.410 104.710 ;
        RECT 557.250 100.720 559.170 104.710 ;
        RECT 560.010 100.720 561.930 104.710 ;
        RECT 562.770 100.720 564.690 104.710 ;
        RECT 565.530 100.720 567.450 104.710 ;
        RECT 568.290 100.720 570.210 104.710 ;
        RECT 571.050 100.720 572.970 104.710 ;
        RECT 573.810 100.720 575.730 104.710 ;
        RECT 576.570 100.720 578.490 104.710 ;
        RECT 579.330 100.720 581.250 104.710 ;
        RECT 582.090 100.720 584.010 104.710 ;
        RECT 584.850 100.720 586.770 104.710 ;
        RECT 587.610 100.720 589.530 104.710 ;
        RECT 590.370 100.720 592.290 104.710 ;
        RECT 593.130 100.720 595.050 104.710 ;
        RECT 595.890 100.720 597.810 104.710 ;
        RECT 598.650 100.720 600.570 104.710 ;
        RECT 601.410 100.720 603.330 104.710 ;
        RECT 604.170 100.720 606.090 104.710 ;
        RECT 606.930 100.720 608.850 104.710 ;
        RECT 609.690 100.720 611.610 104.710 ;
        RECT 612.450 100.720 614.370 104.710 ;
        RECT 615.210 100.720 617.130 104.710 ;
        RECT 617.970 100.720 619.890 104.710 ;
        RECT 620.730 100.720 622.650 104.710 ;
        RECT 623.490 100.720 625.410 104.710 ;
        RECT 626.250 100.720 628.170 104.710 ;
        RECT 629.010 100.720 630.930 104.710 ;
        RECT 631.770 100.720 633.690 104.710 ;
        RECT 634.530 100.720 636.450 104.710 ;
        RECT 637.290 100.720 639.210 104.710 ;
        RECT 640.050 100.720 641.970 104.710 ;
        RECT 642.810 100.720 644.730 104.710 ;
        RECT 645.570 100.720 647.490 104.710 ;
        RECT 648.330 100.720 650.250 104.710 ;
        RECT 651.090 100.720 653.010 104.710 ;
        RECT 653.850 100.720 655.770 104.710 ;
        RECT 656.610 100.720 658.530 104.710 ;
        RECT 659.370 100.720 661.290 104.710 ;
        RECT 662.130 100.720 664.050 104.710 ;
        RECT 664.890 100.720 666.810 104.710 ;
        RECT 667.650 100.720 669.570 104.710 ;
        RECT 670.410 100.720 672.330 104.710 ;
        RECT 673.170 100.720 675.090 104.710 ;
        RECT 675.930 100.720 677.850 104.710 ;
        RECT 678.690 100.720 680.610 104.710 ;
        RECT 681.450 100.720 683.370 104.710 ;
        RECT 684.210 100.720 686.130 104.710 ;
        RECT 686.970 100.720 688.890 104.710 ;
        RECT 689.730 100.720 691.650 104.710 ;
        RECT 692.490 100.720 694.410 104.710 ;
        RECT 695.250 100.720 697.170 104.710 ;
        RECT 698.010 100.720 699.930 104.710 ;
        RECT 700.770 100.720 702.690 104.710 ;
        RECT 703.530 100.720 705.450 104.710 ;
        RECT 706.290 100.720 708.210 104.710 ;
        RECT 709.050 100.720 710.970 104.710 ;
        RECT 711.810 100.720 713.730 104.710 ;
        RECT 714.570 100.720 716.490 104.710 ;
        RECT 717.330 100.720 719.250 104.710 ;
        RECT 720.090 100.720 722.010 104.710 ;
        RECT 722.850 100.720 724.770 104.710 ;
        RECT 725.610 100.720 727.530 104.710 ;
        RECT 728.370 100.720 730.290 104.710 ;
        RECT 731.130 100.720 733.050 104.710 ;
        RECT 733.890 100.720 735.810 104.710 ;
        RECT 736.650 100.720 738.570 104.710 ;
        RECT 739.410 100.720 741.330 104.710 ;
        RECT 742.170 100.720 744.090 104.710 ;
        RECT 744.930 100.720 746.850 104.710 ;
        RECT 747.690 100.720 749.610 104.710 ;
        RECT 750.450 100.720 752.370 104.710 ;
        RECT 753.210 100.720 755.130 104.710 ;
        RECT 755.970 100.720 757.890 104.710 ;
        RECT 758.730 100.720 760.650 104.710 ;
        RECT 761.490 100.720 763.410 104.710 ;
        RECT 764.250 100.720 766.170 104.710 ;
        RECT 767.010 100.720 768.930 104.710 ;
        RECT 769.770 100.720 771.690 104.710 ;
        RECT 772.530 100.720 774.450 104.710 ;
        RECT 775.290 100.720 777.210 104.710 ;
        RECT 778.050 100.720 779.970 104.710 ;
        RECT 780.810 100.720 782.730 104.710 ;
        RECT 783.570 100.720 785.490 104.710 ;
        RECT 786.330 100.720 788.250 104.710 ;
        RECT 789.090 100.720 791.010 104.710 ;
        RECT 791.850 100.720 793.770 104.710 ;
        RECT 794.610 100.720 796.530 104.710 ;
        RECT 797.370 100.720 799.290 104.710 ;
        RECT 800.130 100.720 802.050 104.710 ;
        RECT 802.890 100.720 804.810 104.710 ;
        RECT 805.650 100.720 807.570 104.710 ;
        RECT 808.410 100.720 810.330 104.710 ;
        RECT 811.170 100.720 813.090 104.710 ;
        RECT 813.930 100.720 815.850 104.710 ;
        RECT 816.690 100.720 818.610 104.710 ;
        RECT 819.450 100.720 821.370 104.710 ;
        RECT 822.210 100.720 824.130 104.710 ;
        RECT 824.970 100.720 826.890 104.710 ;
        RECT 827.730 100.720 829.650 104.710 ;
        RECT 830.490 100.720 832.410 104.710 ;
        RECT 833.250 100.720 835.170 104.710 ;
        RECT 836.010 100.720 837.930 104.710 ;
        RECT 838.770 100.720 840.690 104.710 ;
        RECT 841.530 100.720 843.450 104.710 ;
        RECT 844.290 100.720 846.210 104.710 ;
        RECT 847.050 100.720 848.970 104.710 ;
        RECT 849.810 100.720 851.730 104.710 ;
        RECT 852.570 100.720 854.490 104.710 ;
        RECT 855.330 100.720 857.250 104.710 ;
        RECT 858.090 100.720 860.010 104.710 ;
        RECT 860.850 100.720 862.770 104.710 ;
        RECT 863.610 100.720 865.530 104.710 ;
        RECT 866.370 100.720 868.290 104.710 ;
        RECT 869.130 100.720 871.050 104.710 ;
        RECT 871.890 100.720 873.810 104.710 ;
        RECT 874.650 100.720 876.570 104.710 ;
        RECT 877.410 100.720 879.330 104.710 ;
        RECT 880.170 100.720 882.090 104.710 ;
        RECT 882.930 100.720 884.850 104.710 ;
        RECT 885.690 100.720 887.610 104.710 ;
        RECT 888.450 100.720 890.370 104.710 ;
        RECT 891.210 100.720 893.130 104.710 ;
        RECT 893.970 100.720 895.890 104.710 ;
        RECT 896.730 100.720 898.650 104.710 ;
        RECT 899.490 100.720 901.410 104.710 ;
        RECT 902.250 100.720 904.170 104.710 ;
        RECT 905.010 100.720 906.930 104.710 ;
        RECT 907.770 100.720 909.690 104.710 ;
        RECT 910.530 100.720 912.450 104.710 ;
        RECT 913.290 100.720 915.210 104.710 ;
        RECT 916.050 100.720 917.970 104.710 ;
        RECT 918.810 100.720 920.730 104.710 ;
        RECT 921.570 100.720 923.490 104.710 ;
        RECT 924.330 100.720 926.250 104.710 ;
        RECT 927.090 100.720 929.010 104.710 ;
        RECT 929.850 100.720 931.770 104.710 ;
        RECT 932.610 100.720 934.530 104.710 ;
        RECT 935.370 100.720 937.290 104.710 ;
        RECT 938.130 100.720 940.050 104.710 ;
        RECT 940.890 100.720 942.810 104.710 ;
        RECT 943.650 100.720 945.570 104.710 ;
        RECT 946.410 100.720 948.330 104.710 ;
        RECT 949.170 100.720 951.090 104.710 ;
        RECT 951.930 100.720 953.850 104.710 ;
        RECT 954.690 100.720 956.610 104.710 ;
        RECT 957.450 100.720 959.370 104.710 ;
        RECT 960.210 100.720 962.130 104.710 ;
        RECT 962.970 100.720 964.890 104.710 ;
        RECT 965.730 100.720 967.650 104.710 ;
        RECT 968.490 100.720 970.410 104.710 ;
        RECT 971.250 100.720 973.170 104.710 ;
        RECT 974.010 100.720 975.930 104.710 ;
        RECT 976.770 100.720 978.690 104.710 ;
        RECT 979.530 100.720 981.450 104.710 ;
        RECT 982.290 100.720 984.210 104.710 ;
        RECT 985.050 100.720 986.970 104.710 ;
        RECT 987.810 100.720 989.730 104.710 ;
        RECT 990.570 100.720 992.490 104.710 ;
        RECT 993.330 100.720 995.250 104.710 ;
        RECT 996.090 100.720 998.010 104.710 ;
        RECT 998.850 100.720 1000.770 104.710 ;
        RECT 1001.610 100.720 1003.530 104.710 ;
        RECT 1004.370 100.720 1006.290 104.710 ;
        RECT 1007.130 100.720 1009.050 104.710 ;
        RECT 1009.890 100.720 1011.810 104.710 ;
        RECT 1012.650 100.720 1014.570 104.710 ;
        RECT 1015.410 100.720 1017.330 104.710 ;
        RECT 1018.170 100.720 1020.090 104.710 ;
        RECT 1020.930 100.720 1022.850 104.710 ;
        RECT 1023.690 100.720 1025.610 104.710 ;
        RECT 1026.450 100.720 1028.370 104.710 ;
        RECT 1029.210 100.720 1031.130 104.710 ;
        RECT 1031.970 100.720 1033.890 104.710 ;
        RECT 1034.730 100.720 1036.650 104.710 ;
        RECT 1037.490 100.720 1039.410 104.710 ;
        RECT 1040.250 100.720 1042.170 104.710 ;
        RECT 1043.010 100.720 1044.930 104.710 ;
        RECT 1045.770 100.720 1047.690 104.710 ;
        RECT 1048.530 100.720 1050.450 104.710 ;
        RECT 1051.290 100.720 1053.210 104.710 ;
        RECT 1054.050 100.720 1055.970 104.710 ;
        RECT 1056.810 100.720 1058.730 104.710 ;
        RECT 1059.570 100.720 1061.490 104.710 ;
        RECT 1062.330 100.720 1064.250 104.710 ;
        RECT 1065.090 100.720 1067.010 104.710 ;
        RECT 1067.850 100.720 1069.770 104.710 ;
        RECT 1070.610 100.720 1072.530 104.710 ;
        RECT 1073.370 100.720 1075.290 104.710 ;
        RECT 1076.130 100.720 1078.050 104.710 ;
        RECT 1078.890 100.720 1080.810 104.710 ;
        RECT 1081.650 100.720 1083.570 104.710 ;
        RECT 1084.410 100.720 1086.330 104.710 ;
        RECT 1087.170 100.720 1089.090 104.710 ;
        RECT 1089.930 100.720 1091.850 104.710 ;
        RECT 1092.690 100.720 1094.610 104.710 ;
        RECT 1095.450 100.720 1097.370 104.710 ;
        RECT 1098.210 100.720 1100.130 104.710 ;
        RECT 1100.970 100.720 1102.890 104.710 ;
        RECT 1103.730 100.720 1105.650 104.710 ;
        RECT 1106.490 100.720 1108.410 104.710 ;
        RECT 1109.250 100.720 1111.170 104.710 ;
        RECT 1112.010 100.720 1113.930 104.710 ;
        RECT 1114.770 100.720 1116.690 104.710 ;
        RECT 1117.530 100.720 1119.450 104.710 ;
        RECT 1120.290 100.720 1122.210 104.710 ;
        RECT 1123.050 100.720 1124.970 104.710 ;
        RECT 1125.810 100.720 1127.730 104.710 ;
        RECT 1128.570 100.720 1130.490 104.710 ;
        RECT 1131.330 100.720 1133.250 104.710 ;
        RECT 1134.090 100.720 1136.010 104.710 ;
        RECT 1136.850 100.720 1138.770 104.710 ;
        RECT 1139.610 100.720 1141.530 104.710 ;
        RECT 1142.370 100.720 1144.290 104.710 ;
        RECT 1145.130 100.720 1147.050 104.710 ;
        RECT 1147.890 100.720 1149.810 104.710 ;
        RECT 1150.650 100.720 1152.570 104.710 ;
        RECT 1153.410 100.720 1155.330 104.710 ;
        RECT 1156.170 100.720 1158.090 104.710 ;
        RECT 1158.930 100.720 1160.850 104.710 ;
        RECT 1161.690 100.720 1163.610 104.710 ;
        RECT 1164.450 100.720 1166.370 104.710 ;
        RECT 1167.210 100.720 1169.130 104.710 ;
        RECT 1169.970 100.720 1171.890 104.710 ;
        RECT 1172.730 100.720 1174.650 104.710 ;
        RECT 1175.490 100.720 1177.410 104.710 ;
        RECT 1178.250 100.720 1180.170 104.710 ;
        RECT 1181.010 100.720 1182.930 104.710 ;
        RECT 1183.770 100.720 1185.690 104.710 ;
        RECT 1186.530 100.720 1188.450 104.710 ;
        RECT 1189.290 100.720 1191.210 104.710 ;
        RECT 1192.050 100.720 1193.970 104.710 ;
        RECT 1194.810 100.720 1196.730 104.710 ;
        RECT 1197.570 100.720 1199.490 104.710 ;
        RECT 1200.330 100.720 1202.250 104.710 ;
        RECT 1203.090 100.720 1205.010 104.710 ;
        RECT 1205.850 100.720 1207.770 104.710 ;
        RECT 1208.610 100.720 1210.530 104.710 ;
        RECT 1211.370 100.720 1213.290 104.710 ;
        RECT 1214.130 100.720 1216.050 104.710 ;
        RECT 1216.890 100.720 1218.810 104.710 ;
        RECT 1219.650 100.720 1221.570 104.710 ;
        RECT 1222.410 100.720 1224.330 104.710 ;
        RECT 1225.170 100.720 1227.090 104.710 ;
        RECT 1227.930 100.720 1229.850 104.710 ;
        RECT 1230.690 100.720 1232.610 104.710 ;
        RECT 1233.450 100.720 1235.370 104.710 ;
        RECT 1236.210 100.720 1238.130 104.710 ;
        RECT 1238.970 100.720 1240.890 104.710 ;
        RECT 1241.730 100.720 1243.650 104.710 ;
        RECT 1244.490 100.720 1246.410 104.710 ;
        RECT 1247.250 100.720 1249.170 104.710 ;
        RECT 1250.010 100.720 1251.930 104.710 ;
        RECT 1252.770 100.720 1254.690 104.710 ;
        RECT 1255.530 100.720 1257.450 104.710 ;
        RECT 1258.290 100.720 1260.210 104.710 ;
        RECT 1261.050 100.720 1262.970 104.710 ;
        RECT 1263.810 100.720 1265.730 104.710 ;
        RECT 1266.570 100.720 1268.490 104.710 ;
        RECT 1269.330 100.720 1271.250 104.710 ;
        RECT 1272.090 100.720 1274.010 104.710 ;
        RECT 1274.850 100.720 1276.770 104.710 ;
        RECT 1277.610 100.720 1279.530 104.710 ;
        RECT 1280.370 100.720 1282.290 104.710 ;
        RECT 1283.130 100.720 1285.050 104.710 ;
        RECT 1285.890 100.720 1287.810 104.710 ;
        RECT 1288.650 100.720 1290.570 104.710 ;
        RECT 1291.410 100.720 1293.330 104.710 ;
        RECT 1294.170 100.720 1296.090 104.710 ;
        RECT 1296.930 100.720 1298.850 104.710 ;
        RECT 1299.690 100.720 1301.610 104.710 ;
        RECT 1302.450 100.720 1304.370 104.710 ;
        RECT 1305.210 100.720 1307.130 104.710 ;
        RECT 1307.970 100.720 1309.890 104.710 ;
        RECT 1310.730 100.720 1312.650 104.710 ;
        RECT 1313.490 100.720 1315.410 104.710 ;
        RECT 1316.250 100.720 1318.170 104.710 ;
        RECT 1319.010 100.720 1320.930 104.710 ;
        RECT 1321.770 100.720 1323.690 104.710 ;
        RECT 1324.530 100.720 1326.450 104.710 ;
        RECT 1327.290 100.720 1329.210 104.710 ;
        RECT 1330.050 100.720 1331.970 104.710 ;
        RECT 1332.810 100.720 1334.730 104.710 ;
        RECT 1335.570 100.720 1337.490 104.710 ;
        RECT 1338.330 100.720 1340.250 104.710 ;
        RECT 1341.090 100.720 1343.010 104.710 ;
        RECT 1343.850 100.720 1345.770 104.710 ;
        RECT 1346.610 100.720 1348.530 104.710 ;
        RECT 1349.370 100.720 1351.290 104.710 ;
        RECT 1352.130 100.720 1354.050 104.710 ;
        RECT 1354.890 100.720 1356.810 104.710 ;
        RECT 1357.650 100.720 1359.570 104.710 ;
        RECT 1360.410 100.720 1362.330 104.710 ;
        RECT 1363.170 100.720 1365.090 104.710 ;
        RECT 1365.930 100.720 1367.850 104.710 ;
        RECT 1368.690 100.720 1370.610 104.710 ;
        RECT 1371.450 100.720 1373.370 104.710 ;
        RECT 1374.210 100.720 1376.130 104.710 ;
        RECT 1376.970 100.720 1378.890 104.710 ;
        RECT 1379.730 100.720 1381.650 104.710 ;
        RECT 1382.490 100.720 1384.410 104.710 ;
        RECT 1385.250 100.720 1387.170 104.710 ;
        RECT 1388.010 100.720 1389.930 104.710 ;
        RECT 1390.770 100.720 1392.690 104.710 ;
        RECT 1393.530 100.720 1395.450 104.710 ;
        RECT 1396.290 100.720 1398.210 104.710 ;
        RECT 1399.050 100.720 1400.970 104.710 ;
        RECT 1401.810 100.720 1403.730 104.710 ;
        RECT 1404.570 100.720 1406.490 104.710 ;
        RECT 1407.330 100.720 1409.250 104.710 ;
        RECT 1410.090 100.720 1412.010 104.710 ;
        RECT 1412.850 100.720 1414.770 104.710 ;
        RECT 1415.610 100.720 1417.530 104.710 ;
        RECT 1418.370 100.720 1420.290 104.710 ;
        RECT 1421.130 100.720 1423.050 104.710 ;
        RECT 1423.890 100.720 1425.810 104.710 ;
        RECT 1426.650 100.720 1428.570 104.710 ;
        RECT 1429.410 100.720 1431.330 104.710 ;
        RECT 1432.170 100.720 1434.090 104.710 ;
        RECT 1434.930 100.720 1436.850 104.710 ;
        RECT 1437.690 100.720 1439.610 104.710 ;
        RECT 1440.450 100.720 1442.370 104.710 ;
        RECT 1443.210 100.720 1445.130 104.710 ;
        RECT 1445.970 100.720 1447.890 104.710 ;
        RECT 1448.730 100.720 1450.650 104.710 ;
        RECT 1451.490 100.720 1453.410 104.710 ;
        RECT 1454.250 100.720 1456.170 104.710 ;
        RECT 1457.010 100.720 1458.930 104.710 ;
        RECT 1459.770 100.720 1461.690 104.710 ;
        RECT 1462.530 100.720 1464.450 104.710 ;
        RECT 1465.290 100.720 1467.210 104.710 ;
        RECT 1468.050 100.720 1469.970 104.710 ;
        RECT 1470.810 100.720 1472.730 104.710 ;
        RECT 1473.570 100.720 1475.490 104.710 ;
        RECT 1476.330 100.720 1478.250 104.710 ;
        RECT 1479.090 100.720 1481.010 104.710 ;
        RECT 1481.850 100.720 1483.770 104.710 ;
        RECT 1484.610 100.720 1486.530 104.710 ;
        RECT 1487.370 100.720 1489.290 104.710 ;
        RECT 1490.130 100.720 1492.050 104.710 ;
        RECT 1492.890 100.720 1494.810 104.710 ;
        RECT 1495.650 100.720 1497.570 104.710 ;
        RECT 1498.410 100.720 1500.330 104.710 ;
        RECT 1501.170 100.720 1503.090 104.710 ;
        RECT 1503.930 100.720 1505.850 104.710 ;
        RECT 1506.690 100.720 1561.450 104.710 ;
        RECT 20.610 4.280 1561.450 100.720 ;
        RECT 20.610 0.010 62.370 4.280 ;
        RECT 63.210 0.010 66.050 4.280 ;
        RECT 66.890 0.010 69.730 4.280 ;
        RECT 70.570 0.010 73.410 4.280 ;
        RECT 74.250 0.010 77.090 4.280 ;
        RECT 77.930 0.010 80.770 4.280 ;
        RECT 81.610 0.010 84.450 4.280 ;
        RECT 85.290 0.010 88.130 4.280 ;
        RECT 88.970 0.010 91.810 4.280 ;
        RECT 92.650 0.010 95.490 4.280 ;
        RECT 96.330 0.010 99.170 4.280 ;
        RECT 100.010 0.010 102.850 4.280 ;
        RECT 103.690 0.010 106.530 4.280 ;
        RECT 107.370 0.010 110.210 4.280 ;
        RECT 111.050 0.010 113.890 4.280 ;
        RECT 114.730 0.010 117.570 4.280 ;
        RECT 118.410 0.010 121.250 4.280 ;
        RECT 122.090 0.010 124.930 4.280 ;
        RECT 125.770 0.010 128.610 4.280 ;
        RECT 129.450 0.010 132.290 4.280 ;
        RECT 133.130 0.010 135.970 4.280 ;
        RECT 136.810 0.010 139.650 4.280 ;
        RECT 140.490 0.010 143.330 4.280 ;
        RECT 144.170 0.010 147.010 4.280 ;
        RECT 147.850 0.010 150.690 4.280 ;
        RECT 151.530 0.010 154.370 4.280 ;
        RECT 155.210 0.010 158.050 4.280 ;
        RECT 158.890 0.010 161.730 4.280 ;
        RECT 162.570 0.010 165.410 4.280 ;
        RECT 166.250 0.010 169.090 4.280 ;
        RECT 169.930 0.010 172.770 4.280 ;
        RECT 173.610 0.010 176.450 4.280 ;
        RECT 177.290 0.010 180.130 4.280 ;
        RECT 180.970 0.010 183.810 4.280 ;
        RECT 184.650 0.010 187.490 4.280 ;
        RECT 188.330 0.010 191.170 4.280 ;
        RECT 192.010 0.010 194.850 4.280 ;
        RECT 195.690 0.010 198.530 4.280 ;
        RECT 199.370 0.010 202.210 4.280 ;
        RECT 203.050 0.010 205.890 4.280 ;
        RECT 206.730 0.010 209.570 4.280 ;
        RECT 210.410 0.010 213.250 4.280 ;
        RECT 214.090 0.010 216.930 4.280 ;
        RECT 217.770 0.010 220.610 4.280 ;
        RECT 221.450 0.010 224.290 4.280 ;
        RECT 225.130 0.010 227.970 4.280 ;
        RECT 228.810 0.010 231.650 4.280 ;
        RECT 232.490 0.010 235.330 4.280 ;
        RECT 236.170 0.010 239.010 4.280 ;
        RECT 239.850 0.010 242.690 4.280 ;
        RECT 243.530 0.010 246.370 4.280 ;
        RECT 247.210 0.010 250.050 4.280 ;
        RECT 250.890 0.010 253.730 4.280 ;
        RECT 254.570 0.010 257.410 4.280 ;
        RECT 258.250 0.010 261.090 4.280 ;
        RECT 261.930 0.010 264.770 4.280 ;
        RECT 265.610 0.010 268.450 4.280 ;
        RECT 269.290 0.010 272.130 4.280 ;
        RECT 272.970 0.010 275.810 4.280 ;
        RECT 276.650 0.010 279.490 4.280 ;
        RECT 280.330 0.010 283.170 4.280 ;
        RECT 284.010 0.010 286.850 4.280 ;
        RECT 287.690 0.010 290.530 4.280 ;
        RECT 291.370 0.010 294.210 4.280 ;
        RECT 295.050 0.010 297.890 4.280 ;
        RECT 298.730 0.010 301.570 4.280 ;
        RECT 302.410 0.010 305.250 4.280 ;
        RECT 306.090 0.010 308.930 4.280 ;
        RECT 309.770 0.010 312.610 4.280 ;
        RECT 313.450 0.010 316.290 4.280 ;
        RECT 317.130 0.010 319.970 4.280 ;
        RECT 320.810 0.010 323.650 4.280 ;
        RECT 324.490 0.010 327.330 4.280 ;
        RECT 328.170 0.010 331.010 4.280 ;
        RECT 331.850 0.010 334.690 4.280 ;
        RECT 335.530 0.010 338.370 4.280 ;
        RECT 339.210 0.010 342.050 4.280 ;
        RECT 342.890 0.010 345.730 4.280 ;
        RECT 346.570 0.010 349.410 4.280 ;
        RECT 350.250 0.010 353.090 4.280 ;
        RECT 353.930 0.010 356.770 4.280 ;
        RECT 357.610 0.010 360.450 4.280 ;
        RECT 361.290 0.010 364.130 4.280 ;
        RECT 364.970 0.010 367.810 4.280 ;
        RECT 368.650 0.010 371.490 4.280 ;
        RECT 372.330 0.010 375.170 4.280 ;
        RECT 376.010 0.010 378.850 4.280 ;
        RECT 379.690 0.010 382.530 4.280 ;
        RECT 383.370 0.010 386.210 4.280 ;
        RECT 387.050 0.010 389.890 4.280 ;
        RECT 390.730 0.010 393.570 4.280 ;
        RECT 394.410 0.010 397.250 4.280 ;
        RECT 398.090 0.010 400.930 4.280 ;
        RECT 401.770 0.010 404.610 4.280 ;
        RECT 405.450 0.010 408.290 4.280 ;
        RECT 409.130 0.010 411.970 4.280 ;
        RECT 412.810 0.010 415.650 4.280 ;
        RECT 416.490 0.010 419.330 4.280 ;
        RECT 420.170 0.010 423.010 4.280 ;
        RECT 423.850 0.010 426.690 4.280 ;
        RECT 427.530 0.010 430.370 4.280 ;
        RECT 431.210 0.010 434.050 4.280 ;
        RECT 434.890 0.010 437.730 4.280 ;
        RECT 438.570 0.010 1561.450 4.280 ;
      LAYER met3 ;
        RECT 20.590 0.175 1561.470 104.545 ;
  END
END analog_ctrl_regs_APB
END LIBRARY

